netcdf press {
dimensions:
	time = UNLIMITED ; // (0 currently)
	bnds = 2 ;
	rlat = 424 ;
	rlon = 436 ;
variables:
	float lon(rlat, rlon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:_CoordinateAxisType = "Lon" ;
	float lat(rlat, rlon) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:_CoordinateAxisType = "Lat" ;
	float rlat(rlat) ;
		rlat:standard_name = "grid_latitude" ;
		rlat:long_name = "rotated latitude" ;
		rlat:units = "degrees" ;
		rlat:axis = "Y" ;
	int rotated_pole ;
		rotated_pole:long_name = "coordinates of the rotated North Pole" ;
		rotated_pole:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_pole:grid_north_pole_latitude = 39.25f ;
		rotated_pole:grid_north_pole_longitude = -162.f ;
	float rlon(rlon) ;
		rlon:standard_name = "grid_longitude" ;
		rlon:long_name = "rotated longitude" ;
		rlon:units = "degrees" ;
		rlon:axis = "X" ;

// global attributes:
		:CDI = "Climate Data Interface version 1.9.8 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.4" ;
		:conventionsURL = "http://www.cfconventions.org/" ;
		:creation_date = "2020-11-23 14:20:57" ;
		:CDO = "Climate Data Operators version 1.9.8 (https://mpimet.mpg.de/cdo)" ;
data:

 lon =
  -10.37361, -10.27498, -10.17626, -10.07746, -9.978562, -9.879581, 
    -9.780514, -9.681359, -9.582117, -9.482788, -9.383372, -9.283871, 
    -9.184281, -9.084607, -8.984845, -8.884998, -8.785065, -8.685045, 
    -8.58494, -8.48475, -8.384474, -8.284113, -8.183666, -8.083135, 
    -7.982519, -7.881818, -7.781033, -7.680163, -7.579209, -7.478171, 
    -7.377049, -7.275844, -7.174555, -7.073182, -6.971726, -6.870188, 
    -6.768566, -6.666862, -6.565075, -6.463205, -6.361254, -6.259221, 
    -6.157105, -6.054909, -5.95263, -5.850271, -5.74783, -5.645308, 
    -5.542706, -5.440024, -5.337261, -5.234418, -5.131495, -5.028493, 
    -4.925411, -4.822249, -4.719009, -4.61569, -4.512292, -4.408816, 
    -4.305262, -4.20163, -4.09792, -3.994133, -3.890268, -3.786326, 
    -3.682307, -3.578212, -3.474041, -3.369793, -3.265469, -3.16107, 
    -3.056595, -2.952045, -2.84742, -2.742721, -2.637947, -2.533099, 
    -2.428177, -2.323181, -2.218112, -2.112969, -2.007754, -1.902466, 
    -1.797106, -1.691674, -1.586169, -1.480593, -1.374946, -1.269228, 
    -1.163439, -1.05758, -0.9516503, -0.8456509, -0.7395817, -0.6334432, 
    -0.5272356, -0.4209593, -0.3146144, -0.2082014, -0.1017204, 0.004828141, 
    0.111444, 0.2181269, 0.3248765, 0.4316925, 0.5385746, 0.6455226, 
    0.752536, 0.8596146, 0.966758, 1.073966, 1.181238, 1.288574, 1.395974, 
    1.503437, 1.610963, 1.718552, 1.826203, 1.933916, 2.041691, 2.149527, 
    2.257423, 2.365381, 2.473399, 2.581477, 2.689614, 2.797811, 2.906067, 
    3.014381, 3.122754, 3.231184, 3.339672, 3.448218, 3.55682, 3.665478, 
    3.774193, 3.882964, 3.99179, 4.100671, 4.209607, 4.318597, 4.427641, 
    4.536738, 4.645889, 4.755093, 4.864349, 4.973658, 5.083017, 5.192429, 
    5.301891, 5.411404, 5.520967, 5.63058, 5.740243, 5.849954, 5.959714, 
    6.069523, 6.179379, 6.289283, 6.399234, 6.509231, 6.619275, 6.729365, 
    6.8395, 6.94968, 7.059906, 7.170175, 7.280488, 7.390845, 7.501245, 
    7.611687, 7.722172, 7.832698, 7.943266, 8.053875, 8.164525, 8.275214, 
    8.385944, 8.496713, 8.607521, 8.718367, 8.829251, 8.940173, 9.051132, 
    9.162128, 9.27316, 9.384229, 9.495333, 9.606471, 9.717645, 9.828852, 
    9.940093, 10.05137, 10.16268, 10.27402, 10.38539, 10.49679, 10.60823, 
    10.71969, 10.83119, 10.94271, 11.05427, 11.16585, 11.27746, 11.3891, 
    11.50077, 11.61247, 11.72419, 11.83594, 11.94771, 12.05951, 12.17133, 
    12.28318, 12.39505, 12.50695, 12.61887, 12.73081, 12.84277, 12.95475, 
    13.06676, 13.17879, 13.29083, 13.4029, 13.51499, 13.62709, 13.73921, 
    13.85136, 13.96351, 14.07569, 14.18788, 14.30009, 14.41231, 14.52455, 
    14.63681, 14.74907, 14.86136, 14.97365, 15.08596, 15.19828, 15.31061, 
    15.42295, 15.53531, 15.64767, 15.76005, 15.87243, 15.98482, 16.09723, 
    16.20963, 16.32205, 16.43448, 16.54691, 16.65935, 16.77179, 16.88424, 
    16.99669, 17.10914, 17.22161, 17.33407, 17.44654, 17.55901, 17.67148, 
    17.78395, 17.89642, 18.0089, 18.12137, 18.23384, 18.34632, 18.45879, 
    18.57125, 18.68372, 18.79618, 18.90864, 19.0211, 19.13355, 19.246, 
    19.35844, 19.47088, 19.58331, 19.69573, 19.80815, 19.92056, 20.03296, 
    20.14535, 20.25773, 20.3701, 20.48247, 20.59482, 20.70716, 20.81949, 
    20.93181, 21.04411, 21.1564, 21.26868, 21.38095, 21.4932, 21.60544, 
    21.71766, 21.82987, 21.94205, 22.05423, 22.16638, 22.27852, 22.39064, 
    22.50274, 22.61483, 22.72689, 22.83894, 22.95096, 23.06296, 23.17494, 
    23.2869, 23.39884, 23.51076, 23.62265, 23.73451, 23.84636, 23.95818, 
    24.06997, 24.18174, 24.29349, 24.4052, 24.5169, 24.62856, 24.74019, 
    24.8518, 24.96338, 25.07493, 25.18645, 25.29794, 25.4094, 25.52083, 
    25.63223, 25.7436, 25.85493, 25.96624, 26.07751, 26.18874, 26.29994, 
    26.41111, 26.52225, 26.63334, 26.74441, 26.85543, 26.96642, 27.07738, 
    27.18829, 27.29917, 27.41001, 27.52081, 27.63157, 27.7423, 27.85298, 
    27.96362, 28.07423, 28.18479, 28.29531, 28.40579, 28.51622, 28.62662, 
    28.73697, 28.84727, 28.95753, 29.06775, 29.17793, 29.28805, 29.39814, 
    29.50817, 29.61816, 29.72811, 29.838, 29.94785, 30.05765, 30.1674, 
    30.27711, 30.38676, 30.49637, 30.60592, 30.71543, 30.82488, 30.93428, 
    31.04364, 31.15294, 31.26218, 31.37138, 31.48052, 31.58961, 31.69865, 
    31.80763, 31.91656, 32.02543, 32.13425, 32.24301, 32.35172, 32.46036, 
    32.56895, 32.67749, 32.78597, 32.89439, 33.00276, 33.11106, 33.21931, 
    33.3275, 33.43562, 33.54369, 33.6517, 33.75965, 33.86753, 33.97536, 
    34.08313, 34.19083, 34.29847, 34.40605, 34.51357, 34.62102, 34.72841, 
    34.83574, 34.943, 35.05019, 35.15733, 35.2644, 35.3714, 35.47834, 
    35.58521, 35.69201, 35.79875, 35.90543, 36.01203, 36.11857, 36.22504, 
    36.33144, 36.43777, 36.54404, 36.65024, 36.75637, 36.86242,
  -10.42116, -10.3224, -10.22354, -10.12459, -10.02556, -9.92644, -9.827231, 
    -9.727936, -9.628552, -9.529082, -9.429524, -9.329881, -9.230149, 
    -9.130331, -9.030426, -8.930435, -8.830358, -8.730193, -8.629944, 
    -8.529608, -8.429186, -8.328679, -8.228086, -8.127408, -8.026645, 
    -7.925797, -7.824863, -7.723845, -7.622743, -7.521556, -7.420285, 
    -7.31893, -7.21749, -7.115967, -7.01436, -6.912671, -6.810897, -6.709041, 
    -6.607102, -6.50508, -6.402975, -6.300788, -6.198519, -6.096168, 
    -5.993735, -5.891221, -5.788625, -5.685948, -5.583189, -5.48035, 
    -5.377431, -5.274431, -5.17135, -5.06819, -4.96495, -4.86163, -4.758231, 
    -4.654753, -4.551195, -4.447559, -4.343844, -4.240052, -4.13618, 
    -4.032231, -3.928205, -3.824101, -3.71992, -3.615661, -3.511327, 
    -3.406915, -3.302427, -3.197864, -3.093224, -2.988509, -2.883719, 
    -2.778854, -2.673914, -2.568899, -2.46381, -2.358647, -2.25341, -2.1481, 
    -2.042717, -1.93726, -1.831731, -1.726129, -1.620456, -1.51471, 
    -1.408892, -1.303004, -1.197044, -1.091013, -0.9849117, -0.8787402, 
    -0.7724987, -0.6661875, -0.5598069, -0.4533572, -0.3468387, -0.2402516, 
    -0.1335963, -0.02687301, 0.07991789, 0.1867761, 0.2937014, 0.4006934, 
    0.5077519, 0.6148764, 0.7220668, 0.8293227, 0.9366438, 1.04403, 1.15148, 
    1.258995, 1.366574, 1.474216, 1.581922, 1.68969, 1.797521, 1.905415, 
    2.01337, 2.121387, 2.229465, 2.337605, 2.445804, 2.554065, 2.662385, 
    2.770764, 2.879203, 2.987701, 3.096257, 3.204872, 3.313544, 3.422274, 
    3.531061, 3.639905, 3.748806, 3.857762, 3.966774, 4.075841, 4.184964, 
    4.29414, 4.403372, 4.512657, 4.621995, 4.731387, 4.840832, 4.950328, 
    5.059877, 5.169477, 5.27913, 5.388832, 5.498585, 5.608388, 5.718241, 
    5.828143, 5.938094, 6.048093, 6.158141, 6.268236, 6.378379, 6.488569, 
    6.598805, 6.709087, 6.819415, 6.929789, 7.040207, 7.15067, 7.261177, 
    7.371727, 7.482321, 7.592958, 7.703638, 7.814359, 7.925122, 8.035926, 
    8.146771, 8.257656, 8.368582, 8.479547, 8.59055, 8.701593, 8.812675, 
    8.923794, 9.034949, 9.146143, 9.257373, 9.368638, 9.47994, 9.591277, 
    9.702648, 9.814054, 9.925494, 10.03697, 10.14847, 10.26001, 10.37158, 
    10.48319, 10.59482, 10.70649, 10.81818, 10.92991, 11.04166, 11.15345, 
    11.26526, 11.3771, 11.48897, 11.60087, 11.71279, 11.82474, 11.93671, 
    12.04871, 12.16074, 12.27279, 12.38486, 12.49696, 12.60908, 12.72122, 
    12.83339, 12.94558, 13.05779, 13.17001, 13.28226, 13.39453, 13.50682, 
    13.61913, 13.73146, 13.8438, 13.95616, 14.06854, 14.18094, 14.29335, 
    14.40578, 14.51822, 14.63068, 14.74315, 14.85564, 14.96814, 15.08065, 
    15.19317, 15.30571, 15.41826, 15.53082, 15.64338, 15.75596, 15.86855, 
    15.98115, 16.09376, 16.20637, 16.31899, 16.43162, 16.54426, 16.6569, 
    16.76955, 16.8822, 16.99486, 17.10752, 17.22019, 17.33286, 17.44553, 
    17.5582, 17.67088, 17.78355, 17.89623, 18.00891, 18.12159, 18.23427, 
    18.34695, 18.45962, 18.5723, 18.68497, 18.79764, 18.9103, 19.02296, 
    19.13562, 19.24827, 19.36092, 19.47356, 19.58619, 19.69882, 19.81144, 
    19.92406, 20.03666, 20.14926, 20.26184, 20.37442, 20.48699, 20.59955, 
    20.71209, 20.82463, 20.93715, 21.04966, 21.16216, 21.27464, 21.38711, 
    21.49957, 21.61201, 21.72443, 21.83684, 21.94923, 22.06161, 22.17397, 
    22.28631, 22.39864, 22.51094, 22.62323, 22.73549, 22.84774, 22.95997, 
    23.07217, 23.18435, 23.29652, 23.40866, 23.52077, 23.63287, 23.74494, 
    23.85699, 23.96901, 24.081, 24.19297, 24.30492, 24.41684, 24.52873, 
    24.64059, 24.75243, 24.86424, 24.97602, 25.08777, 25.19949, 25.31118, 
    25.42284, 25.53447, 25.64607, 25.75763, 25.86917, 25.98067, 26.09214, 
    26.20357, 26.31497, 26.42634, 26.53767, 26.64896, 26.76023, 26.87145, 
    26.98264, 27.09379, 27.2049, 27.31598, 27.42701, 27.53801, 27.64897, 
    27.75989, 27.87077, 27.9816, 28.0924, 28.20316, 28.31387, 28.42455, 
    28.53518, 28.64576, 28.75631, 28.86681, 28.97726, 29.08767, 29.19804, 
    29.30836, 29.41864, 29.52887, 29.63905, 29.74918, 29.85927, 29.96931, 
    30.0793, 30.18925, 30.29914, 30.40899, 30.51878, 30.62852, 30.73822, 
    30.84786, 30.95745, 31.067, 31.17649, 31.28592, 31.3953, 31.50463, 
    31.61391, 31.72313, 31.8323, 31.94142, 32.05047, 32.15948, 32.26842, 
    32.37732, 32.48615, 32.59493, 32.70365, 32.81231, 32.92092, 33.02946, 
    33.13795, 33.24638, 33.35476, 33.46307, 33.57132, 33.6795, 33.78764, 
    33.8957, 34.00371, 34.11166, 34.21954, 34.32736, 34.43512, 34.54282, 
    34.65045, 34.75801, 34.86552, 34.97296, 35.08034, 35.18765, 35.2949, 
    35.40207, 35.50919, 35.61623, 35.72322, 35.83013, 35.93698, 36.04376, 
    36.15047, 36.25712, 36.36369, 36.4702, 36.57664, 36.68301, 36.78931, 
    36.89554,
  -10.46878, -10.36988, -10.27088, -10.1718, -10.07262, -9.973363, -9.874014, 
    -9.774577, -9.675053, -9.575441, -9.475741, -9.375955, -9.276081, 
    -9.17612, -9.076072, -8.975936, -8.875714, -8.775406, -8.675012, 
    -8.57453, -8.473963, -8.373309, -8.272571, -8.171745, -8.070835, 
    -7.969839, -7.868758, -7.767591, -7.66634, -7.565004, -7.463584, 
    -7.362079, -7.260489, -7.158816, -7.057058, -6.955217, -6.853292, 
    -6.751284, -6.649192, -6.547017, -6.444759, -6.342419, -6.239996, 
    -6.137491, -6.034903, -5.932234, -5.829482, -5.726649, -5.623735, 
    -5.52074, -5.417663, -5.314506, -5.211268, -5.107949, -5.004551, 
    -4.901073, -4.797514, -4.693876, -4.590159, -4.486363, -4.382488, 
    -4.278534, -4.174501, -4.070391, -3.966202, -3.861936, -3.757592, 
    -3.653171, -3.548672, -3.444097, -3.339445, -3.234717, -3.129913, 
    -3.025033, -2.920077, -2.815045, -2.709939, -2.604758, -2.499502, 
    -2.394171, -2.288767, -2.183289, -2.077737, -1.972112, -1.866413, 
    -1.760642, -1.654799, -1.548883, -1.442895, -1.336835, -1.230704, 
    -1.124502, -1.018229, -0.9118851, -0.805471, -0.6989869, -0.5924332, 
    -0.4858099, -0.3791174, -0.2723561, -0.1655262, -0.0586281, 0.04833803, 
    0.1553718, 0.262473, 0.3696412, 0.4768762, 0.5841777, 0.6915452, 
    0.7989787, 0.9064776, 1.014042, 1.121671, 1.229364, 1.337122, 1.444944, 
    1.552829, 1.660778, 1.768789, 1.876863, 1.985, 2.093198, 2.201458, 
    2.309779, 2.418161, 2.526604, 2.635107, 2.74367, 2.852292, 2.960973, 
    3.069714, 3.178513, 3.28737, 3.396285, 3.505257, 3.614286, 3.723372, 
    3.832515, 3.941713, 4.050967, 4.160276, 4.26964, 4.379059, 4.488532, 
    4.598058, 4.707638, 4.817271, 4.926957, 5.036695, 5.146485, 5.256326, 
    5.366219, 5.476161, 5.586155, 5.696198, 5.806291, 5.916433, 6.026624, 
    6.136864, 6.247151, 6.357486, 6.467868, 6.578297, 6.688772, 6.799293, 
    6.90986, 7.020472, 7.131128, 7.241829, 7.352574, 7.463363, 7.574194, 
    7.685069, 7.795985, 7.906943, 8.017943, 8.128984, 8.240066, 8.351187, 
    8.462348, 8.573549, 8.684789, 8.796066, 8.907383, 9.018737, 9.130127, 
    9.241555, 9.353019, 9.464519, 9.576054, 9.687624, 9.799229, 9.910868, 
    10.02254, 10.13425, 10.24599, 10.35776, 10.46956, 10.58139, 10.69326, 
    10.80515, 10.91708, 11.02904, 11.14102, 11.25303, 11.36508, 11.47715, 
    11.58924, 11.70137, 11.81352, 11.9257, 12.0379, 12.15012, 12.26238, 
    12.37465, 12.48695, 12.59928, 12.71162, 12.82399, 12.93638, 13.04879, 
    13.16122, 13.27368, 13.38615, 13.49864, 13.61116, 13.72369, 13.83623, 
    13.9488, 14.06138, 14.17398, 14.2866, 14.39923, 14.51188, 14.62454, 
    14.73722, 14.84991, 14.96261, 15.07533, 15.18806, 15.3008, 15.41355, 
    15.52631, 15.63909, 15.75187, 15.86467, 15.97747, 16.09028, 16.2031, 
    16.31593, 16.42876, 16.5416, 16.65445, 16.7673, 16.88016, 16.99302, 
    17.10589, 17.21876, 17.33164, 17.44452, 17.55739, 17.67028, 17.78316, 
    17.89604, 18.00893, 18.12181, 18.2347, 18.34758, 18.46046, 18.57334, 
    18.68622, 18.79909, 18.91196, 19.02483, 19.13769, 19.25055, 19.3634, 
    19.47625, 19.58909, 19.70192, 19.81475, 19.92757, 20.04038, 20.15318, 
    20.26597, 20.37875, 20.49152, 20.60429, 20.71704, 20.82978, 20.9425, 
    21.05522, 21.16792, 21.28061, 21.39328, 21.50594, 21.61859, 21.73122, 
    21.84383, 21.95643, 22.06901, 22.18157, 22.29412, 22.40664, 22.51915, 
    22.63164, 22.74411, 22.85656, 22.96899, 23.0814, 23.19379, 23.30615, 
    23.41849, 23.53081, 23.64311, 23.75538, 23.86763, 23.97985, 24.09205, 
    24.20422, 24.31637, 24.42849, 24.54058, 24.65265, 24.76469, 24.8767, 
    24.98868, 25.10063, 25.21255, 25.32444, 25.4363, 25.54813, 25.65993, 
    25.77169, 25.88343, 25.99513, 26.10679, 26.21843, 26.33003, 26.44159, 
    26.55312, 26.66462, 26.77607, 26.8875, 26.99888, 27.11023, 27.22154, 
    27.33281, 27.44404, 27.55524, 27.66639, 27.77751, 27.88858, 27.99962, 
    28.11061, 28.22156, 28.33247, 28.44334, 28.55416, 28.66495, 28.77568, 
    28.88638, 28.99703, 29.10763, 29.21819, 29.32871, 29.43917, 29.5496, 
    29.65997, 29.7703, 29.88058, 29.99081, 30.10099, 30.21113, 30.32121, 
    30.43125, 30.54123, 30.65117, 30.76105, 30.87089, 30.98067, 31.0904, 
    31.20008, 31.3097, 31.41927, 31.52879, 31.63825, 31.74766, 31.85702, 
    31.96632, 32.07557, 32.18475, 32.29389, 32.40297, 32.51199, 32.62095, 
    32.72985, 32.8387, 32.94749, 33.05622, 33.16489, 33.27351, 33.38206, 
    33.49055, 33.59899, 33.70736, 33.81567, 33.92392, 34.03211, 34.14024, 
    34.2483, 34.3563, 34.46424, 34.57212, 34.67993, 34.78767, 34.89536, 
    35.00298, 35.11053, 35.21802, 35.32544, 35.4328, 35.54009, 35.64732, 
    35.75447, 35.86156, 35.96859, 36.07554, 36.18243, 36.28925, 36.396, 
    36.50268, 36.60929, 36.71584, 36.82231, 36.92871,
  -10.51647, -10.41742, -10.31829, -10.21906, -10.11975, -10.02035, 
    -9.920862, -9.821284, -9.721619, -9.621865, -9.522024, -9.422094, 
    -9.322078, -9.221973, -9.121781, -9.021502, -8.921137, -8.820683, 
    -8.720144, -8.619517, -8.518805, -8.418005, -8.31712, -8.216147, 
    -8.115089, -8.013947, -7.912717, -7.811402, -7.710002, -7.608517, 
    -7.506947, -7.405292, -7.303552, -7.201728, -7.09982, -6.997827, 
    -6.89575, -6.79359, -6.691346, -6.589018, -6.486607, -6.384113, 
    -6.281536, -6.178876, -6.076134, -5.973309, -5.870402, -5.767414, 
    -5.664343, -5.561191, -5.457958, -5.354643, -5.251247, -5.147771, 
    -5.044214, -4.940577, -4.836859, -4.733062, -4.629185, -4.525228, 
    -4.421192, -4.317077, -4.212883, -4.108611, -4.004261, -3.899832, 
    -3.795325, -3.69074, -3.586078, -3.481339, -3.376523, -3.27163, 
    -3.166661, -3.061615, -2.956494, -2.851296, -2.746023, -2.640675, 
    -2.535252, -2.429754, -2.324182, -2.218536, -2.112815, -2.007021, 
    -1.901153, -1.795213, -1.689199, -1.583113, -1.476954, -1.370724, 
    -1.264421, -1.158047, -1.051602, -0.9450859, -0.8384991, -0.7318419, 
    -0.6251147, -0.5183176, -0.4114511, -0.3045154, -0.1975107, -0.09043746, 
    0.0167041, 0.1239137, 0.2311909, 0.3385356, 0.4459474, 0.5534259, 
    0.6609709, 0.768582, 0.8762591, 0.9840016, 1.091809, 1.199682, 1.307619, 
    1.41562, 1.523686, 1.631815, 1.740007, 1.848262, 1.956579, 2.064959, 
    2.173401, 2.281904, 2.390469, 2.499094, 2.60778, 2.716527, 2.825333, 
    2.934198, 3.043123, 3.152106, 3.261148, 3.370248, 3.479406, 3.588621, 
    3.697893, 3.807222, 3.916607, 4.026048, 4.135544, 4.245096, 4.354702, 
    4.464363, 4.574078, 4.683846, 4.793668, 4.903543, 5.01347, 5.12345, 
    5.233481, 5.343564, 5.453697, 5.563881, 5.674116, 5.7844, 5.894733, 
    6.005116, 6.115547, 6.226027, 6.336554, 6.447129, 6.55775, 6.668419, 
    6.779133, 6.889894, 7.0007, 7.11155, 7.222446, 7.333385, 7.444369, 
    7.555395, 7.666465, 7.777577, 7.888731, 7.999927, 8.111163, 8.222442, 
    8.333759, 8.445118, 8.556516, 8.667953, 8.779428, 8.890942, 9.002493, 
    9.114081, 9.225707, 9.33737, 9.449068, 9.560802, 9.672571, 9.784375, 
    9.896214, 10.00809, 10.11999, 10.23193, 10.3439, 10.4559, 10.56794, 
    10.68, 10.7921, 10.90423, 11.01638, 11.12857, 11.24078, 11.35303, 
    11.4653, 11.5776, 11.68993, 11.80228, 11.91466, 12.02706, 12.13949, 
    12.25195, 12.36442, 12.47693, 12.58945, 12.702, 12.81457, 12.92717, 
    13.03978, 13.15242, 13.26507, 13.37775, 13.49045, 13.60316, 13.7159, 
    13.82865, 13.94142, 14.05421, 14.16701, 14.27983, 14.39267, 14.50552, 
    14.61839, 14.73127, 14.84417, 14.95707, 15.07, 15.18293, 15.29588, 
    15.40883, 15.5218, 15.63478, 15.74777, 15.86077, 15.97378, 16.0868, 
    16.19982, 16.31285, 16.4259, 16.53894, 16.65199, 16.76505, 16.87812, 
    16.99119, 17.10426, 17.21734, 17.33042, 17.4435, 17.55659, 17.66968, 
    17.78276, 17.89585, 18.00895, 18.12204, 18.23512, 18.34821, 18.4613, 
    18.57439, 18.68747, 18.80055, 18.91363, 19.0267, 19.13977, 19.25283, 
    19.36589, 19.47894, 19.59199, 19.70502, 19.81806, 19.93108, 20.0441, 
    20.1571, 20.2701, 20.38309, 20.49607, 20.60904, 20.72199, 20.83493, 
    20.94787, 21.06079, 21.17369, 21.28659, 21.39947, 21.51233, 21.62518, 
    21.73801, 21.85083, 21.96363, 22.07642, 22.18919, 22.30194, 22.41467, 
    22.52738, 22.64007, 22.75275, 22.8654, 22.97803, 23.09064, 23.20324, 
    23.3158, 23.42835, 23.54087, 23.65337, 23.76584, 23.8783, 23.99072, 
    24.10312, 24.2155, 24.32784, 24.44017, 24.55246, 24.66473, 24.77697, 
    24.88918, 25.00136, 25.11351, 25.22563, 25.33772, 25.44979, 25.56182, 
    25.67381, 25.78578, 25.89771, 26.00961, 26.12148, 26.23331, 26.34511, 
    26.45687, 26.5686, 26.6803, 26.79195, 26.90357, 27.01516, 27.1267, 
    27.23821, 27.34968, 27.46111, 27.5725, 27.68385, 27.79516, 27.90644, 
    28.01767, 28.12885, 28.24, 28.35111, 28.46217, 28.57319, 28.68417, 
    28.7951, 28.90599, 29.01683, 29.12763, 29.23838, 29.34909, 29.45975, 
    29.57037, 29.68093, 29.79145, 29.90192, 30.01235, 30.12272, 30.23305, 
    30.34332, 30.45355, 30.56373, 30.67385, 30.78393, 30.89395, 31.00392, 
    31.11384, 31.22371, 31.33352, 31.44328, 31.55299, 31.66264, 31.77224, 
    31.88178, 31.99127, 32.1007, 32.21008, 32.3194, 32.42866, 32.53786, 
    32.64701, 32.7561, 32.86514, 32.97411, 33.08303, 33.19188, 33.30068, 
    33.40942, 33.51809, 33.62671, 33.73526, 33.84376, 33.95219, 34.06056, 
    34.16887, 34.27711, 34.3853, 34.49341, 34.60147, 34.70946, 34.81739, 
    34.92525, 35.03305, 35.14078, 35.24844, 35.35604, 35.46358, 35.57105, 
    35.67845, 35.78578, 35.89305, 36.00025, 36.10738, 36.21444, 36.32143, 
    36.42836, 36.53522, 36.642, 36.74872, 36.85537, 36.96194,
  -10.56422, -10.46504, -10.36576, -10.2664, -10.16695, -10.0674, -9.967775, 
    -9.868057, -9.76825, -9.668355, -9.568372, -9.4683, -9.36814, -9.267893, 
    -9.167558, -9.067135, -8.966624, -8.866027, -8.765342, -8.66457, 
    -8.563711, -8.462766, -8.361733, -8.260614, -8.15941, -8.058118, 
    -7.956741, -7.855278, -7.753729, -7.652095, -7.550375, -7.44857, 
    -7.34668, -7.244705, -7.142645, -7.040501, -6.938273, -6.83596, 
    -6.733563, -6.631083, -6.528518, -6.42587, -6.323139, -6.220325, 
    -6.117428, -6.014448, -5.911386, -5.808241, -5.705014, -5.601706, 
    -5.498315, -5.394843, -5.291289, -5.187654, -5.083939, -4.980143, 
    -4.876266, -4.772309, -4.668272, -4.564155, -4.459958, -4.355682, 
    -4.251327, -4.146893, -4.042379, -3.937788, -3.833118, -3.72837, 
    -3.623545, -3.518641, -3.413661, -3.308603, -3.203469, -3.098258, 
    -2.99297, -2.887607, -2.782167, -2.676652, -2.571062, -2.465396, 
    -2.359656, -2.253841, -2.147952, -2.041988, -1.935951, -1.829841, 
    -1.723657, -1.6174, -1.511071, -1.404669, -1.298195, -1.191649, 
    -1.085032, -0.978343, -0.8715832, -0.7647527, -0.6578519, -0.5508809, 
    -0.4438401, -0.3367297, -0.22955, -0.1223015, -0.01498426, 0.0924013, 
    0.1998549, 0.3073762, 0.414965, 0.5226208, 0.6303434, 0.7381326, 
    0.8459879, 0.953909, 1.061896, 1.169948, 1.278064, 1.386246, 1.494491, 
    1.6028, 1.711174, 1.81961, 1.928109, 2.03667, 2.145294, 2.25398, 
    2.362727, 2.471536, 2.580405, 2.689335, 2.798325, 2.907375, 3.016484, 
    3.125653, 3.234879, 3.344165, 3.453508, 3.56291, 3.672368, 3.781883, 
    3.891455, 4.001083, 4.110767, 4.220507, 4.330301, 4.44015, 4.550054, 
    4.660011, 4.770022, 4.880086, 4.990203, 5.100372, 5.210594, 5.320867, 
    5.431191, 5.541566, 5.651992, 5.762467, 5.872993, 5.983568, 6.094191, 
    6.204863, 6.315583, 6.426351, 6.537166, 6.648028, 6.758936, 6.869891, 
    6.980891, 7.091936, 7.203026, 7.31416, 7.425339, 7.536561, 7.647826, 
    7.759134, 7.870484, 7.981876, 8.093309, 8.204784, 8.316299, 8.427855, 
    8.53945, 8.651084, 8.762757, 8.874469, 8.986218, 9.098005, 9.209829, 
    9.321691, 9.433588, 9.545521, 9.65749, 9.769493, 9.881531, 9.993603, 
    10.10571, 10.21785, 10.33002, 10.44222, 10.55446, 10.66672, 10.77902, 
    10.89135, 11.00371, 11.1161, 11.22851, 11.34096, 11.45343, 11.56593, 
    11.67846, 11.79101, 11.9036, 12.0162, 12.12884, 12.24149, 12.35418, 
    12.46688, 12.57961, 12.69236, 12.80514, 12.91794, 13.03076, 13.14359, 
    13.25646, 13.36934, 13.48224, 13.59516, 13.7081, 13.82105, 13.93403, 
    14.04702, 14.16003, 14.27306, 14.3861, 14.49915, 14.61223, 14.72531, 
    14.83841, 14.95153, 15.06465, 15.17779, 15.29095, 15.40411, 15.51728, 
    15.63047, 15.74366, 15.85687, 15.97008, 16.08331, 16.19654, 16.30978, 
    16.42302, 16.53628, 16.64954, 16.7628, 16.87607, 16.98935, 17.10263, 
    17.21591, 17.3292, 17.44249, 17.55578, 17.66907, 17.78237, 17.89566, 
    18.00896, 18.12226, 18.23555, 18.34885, 18.46214, 18.57544, 18.68872, 
    18.80201, 18.91529, 19.02857, 19.14185, 19.25512, 19.36838, 19.48164, 
    19.59489, 19.70814, 19.82137, 19.9346, 20.04782, 20.16104, 20.27424, 
    20.38744, 20.50062, 20.61379, 20.72695, 20.8401, 20.95324, 21.06637, 
    21.17948, 21.29258, 21.40566, 21.51873, 21.63179, 21.74483, 21.85785, 
    21.97085, 22.08384, 22.19682, 22.30977, 22.42271, 22.53562, 22.64852, 
    22.7614, 22.87426, 22.98709, 23.09991, 23.2127, 23.32547, 23.43822, 
    23.55095, 23.66365, 23.77633, 23.88898, 24.00161, 24.11421, 24.22679, 
    24.33934, 24.45187, 24.56436, 24.67683, 24.78927, 24.90168, 25.01407, 
    25.12642, 25.23874, 25.35104, 25.4633, 25.57553, 25.68773, 25.79989, 
    25.91203, 26.02413, 26.13619, 26.24823, 26.36022, 26.47219, 26.58411, 
    26.69601, 26.80786, 26.91968, 27.03146, 27.14321, 27.25491, 27.36658, 
    27.47821, 27.58979, 27.70134, 27.81285, 27.92432, 28.03575, 28.14713, 
    28.25848, 28.36978, 28.48104, 28.59225, 28.70342, 28.81455, 28.92563, 
    29.03667, 29.14766, 29.25861, 29.36951, 29.48037, 29.59117, 29.70193, 
    29.81265, 29.92331, 30.03393, 30.14449, 30.25501, 30.36548, 30.4759, 
    30.58626, 30.69658, 30.80684, 30.91706, 31.02722, 31.13733, 31.24738, 
    31.35739, 31.46733, 31.57723, 31.68707, 31.79686, 31.90659, 32.01626, 
    32.12588, 32.23544, 32.34495, 32.4544, 32.56379, 32.67313, 32.7824, 
    32.89162, 33.00078, 33.10988, 33.21892, 33.3279, 33.43682, 33.54568, 
    33.65448, 33.76322, 33.87189, 33.98051, 34.08906, 34.19755, 34.30597, 
    34.41434, 34.52264, 34.63087, 34.73904, 34.84715, 34.95519, 35.06317, 
    35.17108, 35.27892, 35.3867, 35.49441, 35.60206, 35.70964, 35.81715, 
    35.92459, 36.03196, 36.13927, 36.24651, 36.35368, 36.46078, 36.56781, 
    36.67477, 36.78166, 36.88848, 36.99522,
  -10.61204, -10.51271, -10.4133, -10.3138, -10.21421, -10.11453, -10.01476, 
    -9.914896, -9.814948, -9.714911, -9.614785, -9.514571, -9.414268, 
    -9.313878, -9.213399, -9.112832, -9.012177, -8.911435, -8.810605, 
    -8.709688, -8.608684, -8.507591, -8.406412, -8.305147, -8.203794, 
    -8.102356, -8.00083, -7.899219, -7.797521, -7.695737, -7.593868, 
    -7.491913, -7.389873, -7.287747, -7.185536, -7.08324, -6.98086, 
    -6.878395, -6.775845, -6.673212, -6.570494, -6.467692, -6.364807, 
    -6.261838, -6.158786, -6.055651, -5.952433, -5.849132, -5.745749, 
    -5.642283, -5.538735, -5.435106, -5.331394, -5.227602, -5.123727, 
    -5.019772, -4.915736, -4.811619, -4.707421, -4.603144, -4.498786, 
    -4.394349, -4.289832, -4.185236, -4.08056, -3.975806, -3.870973, 
    -3.766062, -3.661072, -3.556005, -3.45086, -3.345637, -3.240337, 
    -3.13496, -3.029507, -2.923977, -2.818371, -2.712688, -2.60693, 
    -2.501097, -2.395189, -2.289205, -2.183147, -2.077014, -1.970808, 
    -1.864527, -1.758173, -1.651746, -1.545245, -1.438672, -1.332026, 
    -1.225308, -1.118518, -1.011657, -0.9047238, -0.7977198, -0.6906452, 
    -0.5835, -0.4762847, -0.3689994, -0.2616446, -0.1542205, -0.0467274, 
    0.06083436, 0.1684645, 0.2761627, 0.3839287, 0.491762, 0.5996625, 
    0.7076299, 0.8156637, 0.9237637, 1.031929, 1.140161, 1.248457, 1.356819, 
    1.465245, 1.573735, 1.682289, 1.790907, 1.899588, 2.008332, 2.117138, 
    2.226006, 2.334936, 2.443928, 2.552981, 2.662095, 2.771269, 2.880503, 
    2.989798, 3.099151, 3.208563, 3.318035, 3.427564, 3.537152, 3.646796, 
    3.756499, 3.866258, 3.976073, 4.085945, 4.195872, 4.305855, 4.415893, 
    4.525985, 4.636132, 4.746332, 4.856586, 4.966893, 5.077252, 5.187665, 
    5.298128, 5.408644, 5.51921, 5.629827, 5.740495, 5.851212, 5.961979, 
    6.072795, 6.18366, 6.294573, 6.405534, 6.516543, 6.627599, 6.738701, 
    6.84985, 6.961044, 7.072285, 7.183569, 7.294899, 7.406273, 7.517691, 
    7.629152, 7.740656, 7.852203, 7.963791, 8.075421, 8.187093, 8.298805, 
    8.410559, 8.522351, 8.634183, 8.746055, 8.857965, 8.969913, 9.081899, 
    9.193922, 9.305982, 9.418078, 9.53021, 9.642379, 9.754582, 9.86682, 
    9.979093, 10.0914, 10.20374, 10.31611, 10.42851, 10.54095, 10.65342, 
    10.76592, 10.87845, 10.99101, 11.1036, 11.21622, 11.32886, 11.44154, 
    11.55424, 11.66697, 11.77973, 11.89252, 12.00533, 12.11816, 12.23102, 
    12.34391, 12.45682, 12.56975, 12.68271, 12.79569, 12.90869, 13.02171, 
    13.13475, 13.24782, 13.3609, 13.47401, 13.58714, 13.70028, 13.81344, 
    13.92662, 14.03982, 14.15303, 14.26626, 14.37951, 14.49277, 14.60605, 
    14.71934, 14.83265, 14.94597, 15.0593, 15.17265, 15.28601, 15.39937, 
    15.51276, 15.62615, 15.73955, 15.85296, 15.96638, 16.07981, 16.19325, 
    16.30669, 16.42015, 16.53361, 16.64707, 16.76054, 16.87402, 16.9875, 
    17.10099, 17.21448, 17.32797, 17.44147, 17.55497, 17.66847, 17.78197, 
    17.89547, 18.00898, 18.12248, 18.23598, 18.34949, 18.46299, 18.57648, 
    18.68998, 18.80347, 18.91696, 19.03045, 19.14393, 19.25741, 19.37088, 
    19.48434, 19.5978, 19.71125, 19.8247, 19.93813, 20.05156, 20.16498, 
    20.27839, 20.39179, 20.50518, 20.61856, 20.73193, 20.84528, 20.95863, 
    21.07196, 21.18528, 21.29858, 21.41187, 21.52514, 21.6384, 21.75165, 
    21.86488, 21.97809, 22.09128, 22.20446, 22.31762, 22.43076, 22.54388, 
    22.65698, 22.77007, 22.88313, 22.99617, 23.10919, 23.22219, 23.33516, 
    23.44812, 23.56104, 23.67395, 23.78683, 23.89969, 24.01252, 24.12533, 
    24.23811, 24.35086, 24.46359, 24.57629, 24.68896, 24.8016, 24.91422, 
    25.0268, 25.13935, 25.25188, 25.36437, 25.47684, 25.58927, 25.70167, 
    25.81404, 25.92637, 26.03867, 26.15094, 26.26317, 26.37537, 26.48753, 
    26.59966, 26.71175, 26.8238, 26.93582, 27.0478, 27.15974, 27.27164, 
    27.38351, 27.49534, 27.60712, 27.71887, 27.83057, 27.94224, 28.05386, 
    28.16545, 28.27699, 28.38848, 28.49994, 28.61135, 28.72271, 28.83404, 
    28.94531, 29.05655, 29.16774, 29.27888, 29.38997, 29.50102, 29.61202, 
    29.72297, 29.83388, 29.94474, 30.05555, 30.16631, 30.27701, 30.38767, 
    30.49828, 30.60884, 30.71935, 30.82981, 30.94021, 31.05056, 31.16086, 
    31.2711, 31.3813, 31.49143, 31.60152, 31.71155, 31.82152, 31.93144, 
    32.0413, 32.15111, 32.26086, 32.37055, 32.48019, 32.58977, 32.69929, 
    32.80875, 32.91815, 33.0275, 33.13678, 33.24601, 33.35517, 33.46428, 
    33.57332, 33.6823, 33.79122, 33.90008, 34.00887, 34.11761, 34.22628, 
    34.33489, 34.44343, 34.55191, 34.66033, 34.76868, 34.87696, 34.98518, 
    35.09334, 35.20143, 35.30945, 35.41741, 35.5253, 35.63312, 35.74088, 
    35.84856, 35.95618, 36.06374, 36.17122, 36.27863, 36.38597, 36.49325, 
    36.60045, 36.70759, 36.81465, 36.92164, 37.02856,
  -10.65992, -10.56046, -10.46091, -10.36127, -10.26153, -10.16171, -10.0618, 
    -9.961802, -9.861712, -9.761533, -9.661265, -9.560909, -9.460464, 
    -9.35993, -9.259307, -9.158596, -9.057797, -8.95691, -8.855935, 
    -8.754872, -8.653722, -8.552484, -8.451158, -8.349745, -8.248245, 
    -8.146659, -8.044985, -7.943225, -7.841378, -7.739445, -7.637426, 
    -7.535321, -7.43313, -7.330854, -7.228492, -7.126044, -7.023512, 
    -6.920895, -6.818192, -6.715405, -6.612534, -6.509579, -6.406539, 
    -6.303416, -6.200209, -6.096918, -5.993544, -5.890087, -5.786547, 
    -5.682925, -5.57922, -5.475432, -5.371563, -5.267612, -5.163579, 
    -5.059464, -4.955268, -4.850991, -4.746634, -4.642195, -4.537677, 
    -4.433078, -4.328399, -4.223641, -4.118803, -4.013885, -3.90889, 
    -3.803814, -3.698661, -3.593429, -3.488119, -3.382731, -3.277266, 
    -3.171723, -3.066104, -2.960407, -2.854634, -2.748785, -2.642859, 
    -2.536858, -2.430781, -2.324628, -2.218401, -2.112099, -2.005723, 
    -1.899272, -1.792747, -1.686149, -1.579477, -1.472732, -1.365915, 
    -1.259024, -1.152062, -1.045027, -0.9379212, -0.8307436, -0.7234948, 
    -0.6161753, -0.5087852, -0.4013249, -0.2937947, -0.1861949, -0.07852568, 
    0.0292125, 0.1370194, 0.2448947, 0.3528381, 0.4608492, 0.5689278, 
    0.6770736, 0.7852862, 0.8935652, 1.00191, 1.110322, 1.218798, 1.32734, 
    1.435947, 1.544618, 1.653353, 1.762153, 1.871016, 1.979942, 2.088931, 
    2.197982, 2.307096, 2.416271, 2.525508, 2.634806, 2.744164, 2.853583, 
    2.963063, 3.072601, 3.182199, 3.291857, 3.401572, 3.511346, 3.621178, 
    3.731068, 3.841014, 3.951018, 4.061077, 4.171193, 4.281364, 4.391591, 
    4.501873, 4.612208, 4.722599, 4.833042, 4.94354, 5.05409, 5.164692, 
    5.275347, 5.386054, 5.496812, 5.607621, 5.718481, 5.829391, 5.940351, 
    6.051359, 6.162417, 6.273524, 6.384679, 6.495881, 6.607131, 6.718428, 
    6.829772, 6.941161, 7.052596, 7.164076, 7.275602, 7.387172, 7.498785, 
    7.610443, 7.722143, 7.833887, 7.945672, 8.0575, 8.169369, 8.281279, 
    8.393229, 8.505219, 8.61725, 8.72932, 8.841429, 8.953575, 9.065761, 
    9.177983, 9.290242, 9.402538, 9.514871, 9.627239, 9.739643, 9.852081, 
    9.964554, 10.07706, 10.1896, 10.30217, 10.41478, 10.52742, 10.64009, 
    10.75279, 10.86552, 10.97828, 11.09107, 11.20389, 11.31674, 11.42962, 
    11.54253, 11.65546, 11.76842, 11.88141, 11.99443, 12.10746, 12.22053, 
    12.33362, 12.44673, 12.55987, 12.67303, 12.78621, 12.89942, 13.01265, 
    13.1259, 13.23917, 13.35246, 13.46577, 13.5791, 13.69245, 13.80581, 
    13.9192, 14.0326, 14.14602, 14.25946, 14.37291, 14.48638, 14.59986, 
    14.71336, 14.82687, 14.9404, 15.05394, 15.16749, 15.28106, 15.39463, 
    15.50822, 15.62182, 15.73542, 15.84904, 15.96267, 16.07631, 16.18995, 
    16.3036, 16.41726, 16.53093, 16.6446, 16.75828, 16.87197, 16.98565, 
    17.09935, 17.21305, 17.32675, 17.44045, 17.55416, 17.66786, 17.78157, 
    17.89528, 18.00899, 18.1227, 18.23641, 18.35012, 18.46383, 18.57754, 
    18.69124, 18.80494, 18.91864, 19.03233, 19.14602, 19.2597, 19.37338, 
    19.48705, 19.60072, 19.71437, 19.82803, 19.94167, 20.05531, 20.16893, 
    20.28255, 20.39615, 20.50975, 20.62333, 20.73691, 20.85047, 20.96402, 
    21.07756, 21.19108, 21.30459, 21.41809, 21.53157, 21.64504, 21.75849, 
    21.87192, 21.98534, 22.09874, 22.21212, 22.32549, 22.43883, 22.55216, 
    22.66547, 22.77875, 22.89202, 23.00526, 23.11849, 23.23169, 23.34487, 
    23.45803, 23.57116, 23.68427, 23.79736, 23.91042, 24.02345, 24.13646, 
    24.24945, 24.3624, 24.47533, 24.58824, 24.70111, 24.81396, 24.92677, 
    25.03956, 25.15232, 25.26504, 25.37774, 25.4904, 25.60303, 25.71564, 
    25.8282, 25.94074, 26.05324, 26.16571, 26.27814, 26.39054, 26.5029, 
    26.61523, 26.72752, 26.83977, 26.95199, 27.06417, 27.17631, 27.28841, 
    27.40047, 27.5125, 27.62448, 27.73643, 27.84833, 27.96019, 28.07201, 
    28.18379, 28.29553, 28.40722, 28.51887, 28.63048, 28.74204, 28.85356, 
    28.96503, 29.07646, 29.18785, 29.29918, 29.41047, 29.52171, 29.63291, 
    29.74405, 29.85515, 29.9662, 30.07721, 30.18816, 30.29906, 30.40991, 
    30.52071, 30.63146, 30.74216, 30.85281, 30.9634, 31.07394, 31.18443, 
    31.29487, 31.40525, 31.51558, 31.62585, 31.73607, 31.84623, 31.95634, 
    32.06639, 32.17638, 32.28632, 32.3962, 32.50602, 32.61579, 32.72549, 
    32.83514, 32.94473, 33.05426, 33.16373, 33.27314, 33.38249, 33.49178, 
    33.601, 33.71017, 33.81927, 33.92831, 34.03729, 34.14621, 34.25506, 
    34.36385, 34.47258, 34.58124, 34.68983, 34.79837, 34.90683, 35.01523, 
    35.12357, 35.23183, 35.34004, 35.44817, 35.55624, 35.66424, 35.77217, 
    35.88004, 35.98783, 36.09556, 36.20322, 36.31081, 36.41833, 36.52578, 
    36.63316, 36.74046, 36.8477, 36.95487, 37.06196,
  -10.70787, -10.60827, -10.50858, -10.4088, -10.30893, -10.20897, -10.10891, 
    -10.00877, -9.908543, -9.808223, -9.707812, -9.607313, -9.506725, 
    -9.406048, -9.305282, -9.204427, -9.103484, -9.002452, -8.901332, 
    -8.800123, -8.698827, -8.597442, -8.49597, -8.39441, -8.292763, 
    -8.191028, -8.089206, -7.987298, -7.885302, -7.783219, -7.68105, 
    -7.578795, -7.476454, -7.374026, -7.271513, -7.168914, -7.066229, 
    -6.963459, -6.860604, -6.757664, -6.654639, -6.55153, -6.448336, 
    -6.345058, -6.241696, -6.138249, -6.03472, -5.931107, -5.82741, -5.72363, 
    -5.619768, -5.515823, -5.411795, -5.307685, -5.203493, -5.099219, 
    -4.994864, -4.890427, -4.785909, -4.68131, -4.57663, -4.47187, -4.367029, 
    -4.262108, -4.157108, -4.052028, -3.946868, -3.841629, -3.736311, 
    -3.630915, -3.52544, -3.419887, -3.314256, -3.208548, -3.102762, 
    -2.996898, -2.890958, -2.784941, -2.678848, -2.572678, -2.466433, 
    -2.360111, -2.253715, -2.147243, -2.040697, -1.934076, -1.82738, 
    -1.720611, -1.613768, -1.506851, -1.399861, -1.292799, -1.185663, 
    -1.078455, -0.9711757, -0.8638242, -0.7564012, -0.6489071, -0.5413421, 
    -0.4337066, -0.3260008, -0.2182249, -0.1103795, -0.002464646, 0.1055192, 
    0.2135718, 0.3216929, 0.429882, 0.5381389, 0.6464634, 0.7548549, 
    0.8633133, 0.9718382, 1.080429, 1.189086, 1.297809, 1.406596, 1.515449, 
    1.624366, 1.733347, 1.842392, 1.951501, 2.060673, 2.169907, 2.279204, 
    2.388563, 2.497984, 2.607467, 2.71701, 2.826614, 2.936279, 3.046003, 
    3.155787, 3.265631, 3.375533, 3.485494, 3.595513, 3.70559, 3.815724, 
    3.925916, 4.036164, 4.146468, 4.256828, 4.367244, 4.477715, 4.588241, 
    4.698821, 4.809455, 4.920143, 5.030884, 5.141678, 5.252524, 5.363422, 
    5.474372, 5.585373, 5.696425, 5.807528, 5.918681, 6.029883, 6.141135, 
    6.252435, 6.363784, 6.475181, 6.586625, 6.698116, 6.809655, 6.921239, 
    7.03287, 7.144547, 7.256268, 7.368033, 7.479844, 7.591698, 7.703595, 
    7.815536, 7.927518, 8.039543, 8.15161, 8.263718, 8.375867, 8.488055, 
    8.600285, 8.712553, 8.824861, 8.937207, 9.049591, 9.162013, 9.274473, 
    9.386969, 9.499501, 9.61207, 9.724674, 9.837314, 9.949986, 10.06269, 
    10.17544, 10.28821, 10.40102, 10.51386, 10.62673, 10.73963, 10.85257, 
    10.96553, 11.07853, 11.19155, 11.3046, 11.41768, 11.53079, 11.64393, 
    11.7571, 11.87029, 11.9835, 12.09675, 12.21002, 12.32331, 12.43663, 
    12.54997, 12.66333, 12.77672, 12.89013, 13.00357, 13.11702, 13.2305, 
    13.34399, 13.45751, 13.57104, 13.6846, 13.79817, 13.91176, 14.02537, 
    14.139, 14.25264, 14.3663, 14.47997, 14.59366, 14.70737, 14.82109, 
    14.93482, 15.04857, 15.16232, 15.2761, 15.38988, 15.50367, 15.61748, 
    15.73129, 15.84512, 15.95895, 16.0728, 16.18665, 16.30051, 16.41437, 
    16.52825, 16.64213, 16.75601, 16.86991, 16.9838, 17.0977, 17.21161, 
    17.32552, 17.43943, 17.55334, 17.66726, 17.78117, 17.89509, 18.00901, 
    18.12293, 18.23685, 18.35076, 18.46468, 18.57859, 18.6925, 18.80641, 
    18.92031, 19.03421, 19.14811, 19.262, 19.37589, 19.48977, 19.60364, 
    19.7175, 19.83136, 19.94521, 20.05906, 20.17289, 20.28671, 20.40053, 
    20.51433, 20.62812, 20.7419, 20.85567, 20.96943, 21.08317, 21.1969, 
    21.31062, 21.42432, 21.53801, 21.65168, 21.76534, 21.87898, 21.9926, 
    22.10621, 22.2198, 22.33337, 22.44692, 22.56045, 22.67396, 22.78746, 
    22.90093, 23.01438, 23.12781, 23.24121, 23.3546, 23.46796, 23.5813, 
    23.69461, 23.8079, 23.92117, 24.03441, 24.14762, 24.26081, 24.37397, 
    24.4871, 24.60021, 24.71328, 24.82633, 24.93935, 25.05234, 25.1653, 
    25.27823, 25.39113, 25.50399, 25.61683, 25.72963, 25.8424, 25.95514, 
    26.06784, 26.18051, 26.29314, 26.40574, 26.5183, 26.63083, 26.74332, 
    26.85577, 26.96819, 27.08057, 27.19291, 27.30521, 27.41747, 27.52969, 
    27.64188, 27.75402, 27.86612, 27.97818, 28.0902, 28.20218, 28.31411, 
    28.426, 28.53785, 28.64965, 28.76141, 28.87312, 28.98479, 29.09641, 
    29.20799, 29.31952, 29.43101, 29.54244, 29.65383, 29.76517, 29.87647, 
    29.98771, 30.09891, 30.21005, 30.32114, 30.43219, 30.54318, 30.65412, 
    30.76501, 30.87585, 30.98664, 31.09737, 31.20805, 31.31867, 31.42925, 
    31.53976, 31.65023, 31.76063, 31.87099, 31.98128, 32.09152, 32.2017, 
    32.31182, 32.42189, 32.5319, 32.64186, 32.75175, 32.86158, 32.97136, 
    33.08107, 33.19073, 33.30032, 33.40985, 33.51933, 33.62874, 33.73809, 
    33.84738, 33.9566, 34.06576, 34.17486, 34.2839, 34.39287, 34.50177, 
    34.61061, 34.71939, 34.82811, 34.93675, 35.04533, 35.15385, 35.26229, 
    35.37068, 35.47899, 35.58724, 35.69542, 35.80352, 35.91157, 36.01954, 
    36.12745, 36.23528, 36.34304, 36.45074, 36.55836, 36.66592, 36.7734, 
    36.88081, 36.98815, 37.09542,
  -10.75589, -10.65615, -10.55632, -10.4564, -10.35639, -10.25629, -10.1561, 
    -10.05581, -9.955441, -9.854979, -9.754427, -9.653786, -9.553055, 
    -9.452234, -9.351324, -9.250325, -9.149238, -9.04806, -8.946795, 
    -8.845441, -8.743999, -8.642467, -8.540849, -8.439141, -8.337346, 
    -8.235464, -8.133493, -8.031436, -7.929292, -7.82706, -7.724741, 
    -7.622335, -7.519844, -7.417265, -7.3146, -7.211849, -7.109013, -7.00609, 
    -6.903082, -6.799989, -6.69681, -6.593547, -6.490198, -6.386765, 
    -6.283248, -6.179646, -6.07596, -5.972191, -5.868338, -5.7644, -5.660381, 
    -5.556278, -5.452092, -5.347823, -5.243472, -5.139039, -5.034523, 
    -4.929926, -4.825248, -4.720488, -4.615647, -4.510725, -4.405722, 
    -4.300639, -4.195475, -4.090232, -3.984909, -3.879506, -3.774024, 
    -3.668463, -3.562823, -3.457105, -3.351308, -3.245433, -3.13948, 
    -3.03345, -2.927343, -2.821158, -2.714897, -2.608559, -2.502145, 
    -2.395654, -2.289088, -2.182447, -2.07573, -1.968939, -1.862072, 
    -1.755132, -1.648117, -1.541028, -1.433866, -1.326631, -1.219322, 
    -1.111941, -1.004488, -0.8969622, -0.7893648, -0.6816959, -0.5739558, 
    -0.4661447, -0.3582631, -0.2503111, -0.1422891, -0.03419743, 0.07396364, 
    0.1821938, 0.2904927, 0.3988601, 0.5072955, 0.6157989, 0.7243696, 
    0.8330076, 0.9417124, 1.050484, 1.159321, 1.268225, 1.377193, 1.486228, 
    1.595326, 1.70449, 1.813717, 1.923009, 2.032364, 2.141782, 2.251263, 
    2.360806, 2.470411, 2.580078, 2.689807, 2.799596, 2.909446, 3.019357, 
    3.129327, 3.239357, 3.349446, 3.459594, 3.569801, 3.680065, 3.790388, 
    3.900767, 4.011204, 4.121697, 4.232246, 4.342852, 4.453513, 4.564229, 
    4.674999, 4.785824, 4.896702, 5.007635, 5.11862, 5.229658, 5.340748, 
    5.45189, 5.563084, 5.674329, 5.785625, 5.89697, 6.008366, 6.119812, 
    6.231306, 6.342849, 6.454441, 6.56608, 6.677766, 6.7895, 6.90128, 
    7.013107, 7.124979, 7.236897, 7.348859, 7.460865, 7.572917, 7.685011, 
    7.797149, 7.909329, 8.021552, 8.133817, 8.246123, 8.358471, 8.470859, 
    8.583286, 8.695754, 8.808261, 8.920807, 9.033391, 9.146013, 9.258673, 
    9.371369, 9.484102, 9.596871, 9.709677, 9.822516, 9.935391, 10.0483, 
    10.16124, 10.27422, 10.38723, 10.50027, 10.61335, 10.72645, 10.83959, 
    10.95275, 11.06595, 11.17918, 11.29244, 11.40572, 11.51903, 11.63238, 
    11.74574, 11.85914, 11.97256, 12.08601, 12.19948, 12.31298, 12.4265, 
    12.54005, 12.65362, 12.76721, 12.88083, 12.99447, 13.10813, 13.22181, 
    13.33551, 13.44923, 13.56297, 13.67673, 13.79051, 13.90431, 14.01813, 
    14.13196, 14.24581, 14.35967, 14.47355, 14.58745, 14.70136, 14.81529, 
    14.92923, 15.04318, 15.15715, 15.27112, 15.38512, 15.49912, 15.61313, 
    15.72715, 15.84118, 15.95523, 16.06928, 16.18334, 16.29741, 16.41148, 
    16.52556, 16.63965, 16.75374, 16.86784, 16.98195, 17.09606, 17.21017, 
    17.32429, 17.4384, 17.55253, 17.66665, 17.78078, 17.8949, 18.00903, 
    18.12315, 18.23728, 18.3514, 18.46553, 18.57965, 18.69377, 18.80788, 
    18.922, 19.0361, 19.15021, 19.26431, 19.3784, 19.49249, 19.60657, 
    19.72064, 19.83471, 19.94876, 20.06281, 20.17685, 20.29089, 20.40491, 
    20.51892, 20.63292, 20.7469, 20.86088, 20.97485, 21.0888, 21.20273, 
    21.31666, 21.43057, 21.54446, 21.65834, 21.7722, 21.88605, 21.99988, 
    22.11369, 22.22749, 22.34126, 22.45502, 22.56876, 22.68248, 22.79618, 
    22.90985, 23.02351, 23.13714, 23.25076, 23.36435, 23.47791, 23.59146, 
    23.70498, 23.81847, 23.93194, 24.04538, 24.1588, 24.27219, 24.38556, 
    24.49889, 24.6122, 24.72548, 24.83873, 24.95196, 25.06515, 25.17831, 
    25.29144, 25.40454, 25.51761, 25.63065, 25.74365, 25.85662, 25.96956, 
    26.08247, 26.19534, 26.30817, 26.42097, 26.53373, 26.64646, 26.75915, 
    26.87181, 26.98442, 27.097, 27.20954, 27.32204, 27.4345, 27.54692, 
    27.6593, 27.77164, 27.88394, 27.9962, 28.10842, 28.22059, 28.33272, 
    28.44481, 28.55685, 28.66886, 28.78081, 28.89272, 29.00459, 29.11641, 
    29.22818, 29.3399, 29.45158, 29.56322, 29.6748, 29.78633, 29.89782, 
    30.00926, 30.12065, 30.23198, 30.34327, 30.45451, 30.56569, 30.67683, 
    30.78791, 30.89894, 31.00992, 31.12084, 31.23171, 31.34253, 31.45329, 
    31.564, 31.67465, 31.78524, 31.89578, 32.00627, 32.1167, 32.22707, 
    32.33738, 32.44764, 32.55783, 32.66797, 32.77805, 32.88807, 32.99803, 
    33.10793, 33.21777, 33.32756, 33.43727, 33.54693, 33.65652, 33.76606, 
    33.87553, 33.98494, 34.09428, 34.20356, 34.31278, 34.42194, 34.53102, 
    34.64005, 34.74901, 34.8579, 34.96673, 35.07549, 35.18418, 35.29281, 
    35.40137, 35.50986, 35.61829, 35.72664, 35.83493, 35.94315, 36.0513, 
    36.15938, 36.26739, 36.37533, 36.4832, 36.591, 36.69873, 36.80639, 
    36.91397, 37.02149, 37.12893,
  -10.80398, -10.7041, -10.60413, -10.50407, -10.40392, -10.30368, -10.20334, 
    -10.10292, -10.00241, -9.901803, -9.801109, -9.700325, -9.599451, 
    -9.498487, -9.397433, -9.29629, -9.195058, -9.093737, -8.992326, 
    -8.890826, -8.789237, -8.68756, -8.585794, -8.48394, -8.381997, 
    -8.279967, -8.177849, -8.075643, -7.973348, -7.870967, -7.768498, 
    -7.665943, -7.5633, -7.46057, -7.357754, -7.254851, -7.151862, -7.048787, 
    -6.945626, -6.84238, -6.739047, -6.635629, -6.532126, -6.428538, 
    -6.324865, -6.221108, -6.117266, -6.01334, -5.90933, -5.805236, 
    -5.701058, -5.596797, -5.492453, -5.388025, -5.283515, -5.178923, 
    -5.074247, -4.96949, -4.864651, -4.759729, -4.654727, -4.549643, 
    -4.444478, -4.339232, -4.233906, -4.1285, -4.023012, -3.917446, 
    -3.811799, -3.706073, -3.600268, -3.494384, -3.388422, -3.28238, 
    -3.176261, -3.070064, -2.963789, -2.857436, -2.751007, -2.6445, 
    -2.537917, -2.431258, -2.324522, -2.217711, -2.110824, -2.003861, 
    -1.896824, -1.789712, -1.682525, -1.575264, -1.46793, -1.360522, 
    -1.25304, -1.145485, -1.037858, -0.930158, -0.8223859, -0.714542, 
    -0.6066265, -0.4986398, -0.3905821, -0.2824537, -0.174255, -0.06598622, 
    0.04235228, 0.1507602, 0.2592372, 0.367783, 0.4763973, 0.5850797, 
    0.69383, 0.8026478, 0.9115327, 1.020484, 1.129503, 1.238587, 1.347738, 
    1.456953, 1.566234, 1.67558, 1.784991, 1.894465, 2.004003, 2.113605, 
    2.22327, 2.332998, 2.442788, 2.55264, 2.662553, 2.772528, 2.882565, 
    2.992661, 3.102818, 3.213035, 3.323311, 3.433646, 3.544041, 3.654493, 
    3.765004, 3.875572, 3.986198, 4.09688, 4.207619, 4.318414, 4.429265, 
    4.540171, 4.651132, 4.762148, 4.873218, 4.984341, 5.095519, 5.206748, 
    5.318031, 5.429366, 5.540752, 5.65219, 5.76368, 5.875219, 5.986809, 
    6.098448, 6.210137, 6.321875, 6.433661, 6.545495, 6.657377, 6.769307, 
    6.881283, 6.993305, 7.105374, 7.217488, 7.329647, 7.441851, 7.5541, 
    7.666391, 7.778727, 7.891106, 8.003527, 8.11599, 8.228495, 8.341041, 
    8.453628, 8.566256, 8.678923, 8.791629, 8.904375, 9.017159, 9.129981, 
    9.242842, 9.355739, 9.468673, 9.581643, 9.69465, 9.807692, 9.920768, 
    10.03388, 10.14702, 10.2602, 10.37341, 10.48666, 10.59994, 10.71324, 
    10.82658, 10.93995, 11.05336, 11.16679, 11.28025, 11.39373, 11.50725, 
    11.6208, 11.73437, 11.84797, 11.9616, 12.07525, 12.18893, 12.30263, 
    12.41636, 12.53011, 12.64389, 12.75769, 12.87151, 12.98535, 13.09922, 
    13.2131, 13.32701, 13.44094, 13.55489, 13.66885, 13.78284, 13.89684, 
    14.01087, 14.1249, 14.23896, 14.35303, 14.46712, 14.58123, 14.69534, 
    14.80948, 14.92363, 15.03779, 15.15196, 15.26615, 15.38034, 15.49455, 
    15.60877, 15.723, 15.83724, 15.95149, 16.06575, 16.18002, 16.2943, 
    16.40858, 16.52287, 16.63717, 16.75147, 16.86578, 16.98009, 17.0944, 
    17.20873, 17.32305, 17.43738, 17.55171, 17.66604, 17.78037, 17.89471, 
    18.00904, 18.12338, 18.23771, 18.35205, 18.46638, 18.58071, 18.69503, 
    18.80936, 18.92368, 19.03799, 19.15231, 19.26661, 19.38091, 19.49521, 
    19.6095, 19.72378, 19.83805, 19.95232, 20.06658, 20.18083, 20.29507, 
    20.4093, 20.52351, 20.63772, 20.75192, 20.8661, 20.98027, 21.09443, 
    21.20858, 21.32271, 21.43682, 21.55093, 21.66501, 21.77908, 21.89314, 
    22.00717, 22.12119, 22.23519, 22.34917, 22.46314, 22.57708, 22.69101, 
    22.80491, 22.9188, 23.03266, 23.1465, 23.26032, 23.37411, 23.48788, 
    23.60163, 23.71536, 23.82906, 23.94273, 24.05638, 24.17, 24.2836, 
    24.39717, 24.51071, 24.62422, 24.7377, 24.85116, 24.96458, 25.07798, 
    25.19135, 25.30468, 25.41798, 25.53126, 25.6445, 25.7577, 25.87088, 
    25.98402, 26.09712, 26.21019, 26.32323, 26.43623, 26.54919, 26.66212, 
    26.77501, 26.88787, 27.00068, 27.11346, 27.2262, 27.3389, 27.45156, 
    27.56418, 27.67677, 27.7893, 27.9018, 28.01426, 28.12667, 28.23905, 
    28.35137, 28.46366, 28.5759, 28.6881, 28.80025, 28.91236, 29.02442, 
    29.13643, 29.2484, 29.36032, 29.4722, 29.58402, 29.6958, 29.80753, 
    29.91921, 30.03085, 30.14243, 30.25396, 30.36544, 30.47687, 30.58825, 
    30.69958, 30.81085, 30.92207, 31.03324, 31.14436, 31.25542, 31.36642, 
    31.47738, 31.58827, 31.69912, 31.8099, 31.92063, 32.03131, 32.14192, 
    32.25248, 32.36298, 32.47343, 32.58381, 32.69414, 32.80441, 32.91461, 
    33.02476, 33.13485, 33.24487, 33.35484, 33.46474, 33.57458, 33.68436, 
    33.79408, 33.90374, 34.01333, 34.12286, 34.23232, 34.34172, 34.45106, 
    34.56033, 34.66953, 34.77867, 34.88774, 34.99675, 35.1057, 35.21457, 
    35.32338, 35.43212, 35.54079, 35.64939, 35.75793, 35.86639, 35.97479, 
    36.08312, 36.19138, 36.29956, 36.40768, 36.51573, 36.6237, 36.73161, 
    36.83944, 36.9472, 37.05489, 37.1625,
  -10.85213, -10.75212, -10.65201, -10.55181, -10.45152, -10.35113, 
    -10.25066, -10.1501, -10.04944, -9.948696, -9.847859, -9.746933, 
    -9.645916, -9.544808, -9.443611, -9.342324, -9.240947, -9.139481, 
    -9.037925, -8.936279, -8.834544, -8.73272, -8.630808, -8.528807, 
    -8.426716, -8.324537, -8.222271, -8.119915, -8.017472, -7.914941, 
    -7.812323, -7.709617, -7.606823, -7.503942, -7.400974, -7.29792, 
    -7.194778, -7.091551, -6.988236, -6.884836, -6.78135, -6.677778, 
    -6.574121, -6.470377, -6.366549, -6.262636, -6.158638, -6.054555, 
    -5.950388, -5.846137, -5.741801, -5.637382, -5.532879, -5.428293, 
    -5.323623, -5.218871, -5.114036, -5.009118, -4.904118, -4.799036, 
    -4.693871, -4.588625, -4.483298, -4.37789, -4.2724, -4.16683, -4.061179, 
    -3.955448, -3.849637, -3.743746, -3.637776, -3.531726, -3.425597, 
    -3.31939, -3.213104, -3.106739, -3.000296, -2.893776, -2.787178, 
    -2.680503, -2.573751, -2.466922, -2.360016, -2.253035, -2.145977, 
    -2.038844, -1.931635, -1.824352, -1.716993, -1.60956, -1.502053, 
    -1.394471, -1.286816, -1.179088, -1.071286, -0.9634118, -0.8554649, 
    -0.7474458, -0.6393547, -0.5311921, -0.4229581, -0.3146531, -0.2062774, 
    -0.09783138, 0.01068477, 0.1192707, 0.227926, 0.3366505, 0.4454438, 
    0.5543056, 0.6632355, 0.7722334, 0.8812987, 0.9904311, 1.09963, 1.208896, 
    1.318228, 1.427626, 1.53709, 1.646618, 1.756211, 1.865869, 1.975591, 
    2.085377, 2.195226, 2.305138, 2.415113, 2.525151, 2.63525, 2.745411, 
    2.855633, 2.965916, 3.07626, 3.186664, 3.297127, 3.407651, 3.518233, 
    3.628874, 3.739573, 3.85033, 3.961145, 4.072017, 4.182946, 4.293931, 
    4.404972, 4.516068, 4.627221, 4.738428, 4.849689, 4.961004, 5.072373, 
    5.183795, 5.295271, 5.406798, 5.518378, 5.63001, 5.741693, 5.853426, 
    5.965209, 6.077044, 6.188927, 6.30086, 6.412841, 6.524871, 6.636949, 
    6.749074, 6.861247, 6.973465, 7.085731, 7.198042, 7.310399, 7.4228, 
    7.535246, 7.647736, 7.76027, 7.872847, 7.985466, 8.098128, 8.210832, 
    8.323577, 8.436364, 8.549191, 8.662058, 8.774964, 8.887911, 9.000896, 
    9.113918, 9.226979, 9.340078, 9.453214, 9.566385, 9.679593, 9.792837, 
    9.906116, 10.01943, 10.13278, 10.24616, 10.35957, 10.47302, 10.5865, 
    10.70001, 10.81355, 10.92713, 11.04073, 11.15437, 11.26803, 11.38173, 
    11.49545, 11.6092, 11.72297, 11.83678, 11.95061, 12.06447, 12.17835, 
    12.29226, 12.40619, 12.52015, 12.63413, 12.74814, 12.86217, 12.97622, 
    13.09029, 13.20438, 13.3185, 13.43263, 13.54678, 13.66096, 13.77515, 
    13.88936, 14.00359, 14.11784, 14.2321, 14.34638, 14.46068, 14.57499, 
    14.68932, 14.80366, 14.91801, 15.03238, 15.14676, 15.26116, 15.37556, 
    15.48998, 15.60441, 15.71885, 15.83329, 15.94775, 16.06222, 16.1767, 
    16.29118, 16.40567, 16.52017, 16.63468, 16.74919, 16.8637, 16.97823, 
    17.09275, 17.20728, 17.32181, 17.43635, 17.55089, 17.66543, 17.77997, 
    17.89452, 18.00906, 18.1236, 18.23815, 18.35269, 18.46723, 18.58177, 
    18.6963, 18.81084, 18.92537, 19.03989, 19.15441, 19.26893, 19.38344, 
    19.49794, 19.61244, 19.72693, 19.84141, 19.95589, 20.07035, 20.18481, 
    20.29926, 20.41369, 20.52812, 20.64254, 20.75694, 20.87133, 20.98571, 
    21.10008, 21.21443, 21.32877, 21.44309, 21.5574, 21.6717, 21.78597, 
    21.90023, 22.01448, 22.12871, 22.24291, 22.3571, 22.47128, 22.58543, 
    22.69956, 22.81367, 22.92776, 23.04183, 23.15587, 23.2699, 23.3839, 
    23.49788, 23.61183, 23.72576, 23.83966, 23.95354, 24.0674, 24.18122, 
    24.29502, 24.4088, 24.52254, 24.63626, 24.74995, 24.86361, 24.97724, 
    25.09084, 25.20441, 25.31795, 25.43145, 25.54493, 25.65837, 25.77178, 
    25.88516, 25.9985, 26.1118, 26.22508, 26.33832, 26.45152, 26.56469, 
    26.67781, 26.79091, 26.90396, 27.01698, 27.12996, 27.2429, 27.3558, 
    27.46866, 27.58148, 27.69426, 27.807, 27.9197, 28.03235, 28.14496, 
    28.25753, 28.37006, 28.48254, 28.59498, 28.70738, 28.81973, 28.93203, 
    29.04429, 29.1565, 29.26867, 29.38078, 29.49285, 29.60488, 29.71685, 
    29.82877, 29.94065, 30.05248, 30.16425, 30.27598, 30.38765, 30.49928, 
    30.61085, 30.72237, 30.83383, 30.94525, 31.05661, 31.16792, 31.27917, 
    31.39037, 31.50151, 31.6126, 31.72363, 31.83461, 31.94553, 32.05639, 
    32.16719, 32.27794, 32.38863, 32.49926, 32.60984, 32.72035, 32.8308, 
    32.9412, 33.05153, 33.16181, 33.27202, 33.38217, 33.49226, 33.60229, 
    33.71225, 33.82215, 33.932, 34.04177, 34.15148, 34.26113, 34.37071, 
    34.48023, 34.58968, 34.69907, 34.80839, 34.91765, 35.02684, 35.13596, 
    35.24501, 35.354, 35.46292, 35.57177, 35.68055, 35.78926, 35.89791, 
    36.00648, 36.11499, 36.22343, 36.33179, 36.44008, 36.54831, 36.65646, 
    36.76454, 36.87255, 36.98048, 37.08834, 37.19613,
  -10.90036, -10.8002, -10.69995, -10.59961, -10.49918, -10.39866, -10.29805, 
    -10.19734, -10.09655, -9.995657, -9.894679, -9.79361, -9.69245, 
    -9.591199, -9.489858, -9.388426, -9.286904, -9.185293, -9.083591, 
    -8.9818, -8.879919, -8.777949, -8.675889, -8.573741, -8.471502, 
    -8.369176, -8.266761, -8.164256, -8.061664, -7.958983, -7.856215, 
    -7.753358, -7.650414, -7.547381, -7.444262, -7.341055, -7.237762, 
    -7.134381, -7.030914, -6.92736, -6.82372, -6.719994, -6.616181, 
    -6.512283, -6.408299, -6.30423, -6.200076, -6.095836, -5.991512, 
    -5.887103, -5.78261, -5.678032, -5.573371, -5.468626, -5.363797, 
    -5.258884, -5.153889, -5.04881, -4.94365, -4.838406, -4.73308, -4.627672, 
    -4.522182, -4.416611, -4.310958, -4.205225, -4.09941, -3.993514, 
    -3.887538, -3.781482, -3.675347, -3.569131, -3.462836, -3.356462, 
    -3.250008, -3.143476, -3.036866, -2.930178, -2.823411, -2.716567, 
    -2.609646, -2.502647, -2.395572, -2.28842, -2.181191, -2.073887, 
    -1.966507, -1.859052, -1.751521, -1.643915, -1.536235, -1.42848, 
    -1.320652, -1.212749, -1.104773, -0.9967241, -0.8886021, -0.7804075, 
    -0.6721408, -0.563802, -0.4553915, -0.3469097, -0.2383569, -0.1297333, 
    -0.02103924, 0.08772489, 0.1965588, 0.3054622, 0.4144348, 0.5234761, 
    0.6325861, 0.7417641, 0.85101, 0.9603235, 1.069704, 1.179152, 1.288666, 
    1.398246, 1.507892, 1.617603, 1.72738, 1.837221, 1.947127, 2.057097, 
    2.167131, 2.277228, 2.387388, 2.497611, 2.607896, 2.718243, 2.828652, 
    2.939121, 3.049652, 3.160244, 3.270895, 3.381606, 3.492377, 3.603206, 
    3.714094, 3.825041, 3.936045, 4.047107, 4.158226, 4.269401, 4.380633, 
    4.49192, 4.603264, 4.714662, 4.826116, 4.937623, 5.049184, 5.1608, 
    5.272468, 5.384188, 5.495962, 5.607787, 5.719663, 5.831591, 5.94357, 
    6.055598, 6.167677, 6.279805, 6.391982, 6.504208, 6.616481, 6.728803, 
    6.841172, 6.953588, 7.06605, 7.178558, 7.291112, 7.403712, 7.516356, 
    7.629044, 7.741776, 7.854552, 7.96737, 8.080232, 8.193134, 8.30608, 
    8.419065, 8.532093, 8.64516, 8.758267, 8.871414, 8.9846, 9.097824, 
    9.211086, 9.324386, 9.437723, 9.551097, 9.664507, 9.777953, 9.891434, 
    10.00495, 10.1185, 10.23209, 10.3457, 10.45935, 10.57304, 10.68675, 
    10.8005, 10.91428, 11.02809, 11.14192, 11.25579, 11.36969, 11.48362, 
    11.59757, 11.71156, 11.82557, 11.9396, 12.05367, 12.16776, 12.28187, 
    12.39601, 12.51017, 12.62436, 12.73857, 12.85281, 12.96706, 13.08134, 
    13.19564, 13.30996, 13.4243, 13.53867, 13.65305, 13.76745, 13.88187, 
    13.9963, 14.11076, 14.22523, 14.33972, 14.45422, 14.56874, 14.68327, 
    14.79782, 14.91239, 15.02696, 15.14155, 15.25616, 15.37077, 15.4854, 
    15.60003, 15.71468, 15.82934, 15.94401, 16.05868, 16.17337, 16.28806, 
    16.40276, 16.51747, 16.63218, 16.7469, 16.86163, 16.97636, 17.09109, 
    17.20583, 17.32058, 17.43532, 17.55007, 17.66482, 17.77957, 17.89432, 
    18.00908, 18.12383, 18.23858, 18.35333, 18.46808, 18.58283, 18.69758, 
    18.81232, 18.92706, 19.04179, 19.15652, 19.27125, 19.38597, 19.50068, 
    19.61538, 19.73008, 19.84477, 19.95946, 20.07413, 20.1888, 20.30346, 
    20.4181, 20.53274, 20.64736, 20.76197, 20.87657, 20.99116, 21.10574, 
    21.2203, 21.33484, 21.44938, 21.56389, 21.67839, 21.79288, 21.90735, 
    22.0218, 22.13623, 22.25065, 22.36505, 22.47943, 22.59378, 22.70812, 
    22.82244, 22.93674, 23.05101, 23.16527, 23.2795, 23.3937, 23.50789, 
    23.62205, 23.73618, 23.85029, 23.96438, 24.07844, 24.19247, 24.30648, 
    24.42045, 24.5344, 24.64833, 24.76222, 24.87609, 24.98992, 25.10372, 
    25.21749, 25.33124, 25.44495, 25.55863, 25.67227, 25.78588, 25.89946, 
    26.01301, 26.12652, 26.23999, 26.35344, 26.46684, 26.58021, 26.69354, 
    26.80683, 26.92009, 27.03331, 27.14649, 27.25963, 27.37273, 27.48579, 
    27.59881, 27.71179, 27.82473, 27.93762, 28.05048, 28.16329, 28.27606, 
    28.38878, 28.50147, 28.6141, 28.72669, 28.83924, 28.95174, 29.0642, 
    29.17661, 29.28897, 29.40128, 29.51355, 29.62577, 29.73794, 29.85006, 
    29.96213, 30.07415, 30.18612, 30.29804, 30.40991, 30.52172, 30.63349, 
    30.7452, 30.85686, 30.96847, 31.08002, 31.19152, 31.30296, 31.41435, 
    31.52569, 31.63697, 31.74819, 31.85936, 31.97046, 32.08152, 32.19251, 
    32.30345, 32.41433, 32.52515, 32.63591, 32.74661, 32.85725, 32.96783, 
    33.07836, 33.18882, 33.29922, 33.40955, 33.51983, 33.63004, 33.74019, 
    33.85028, 33.9603, 34.07026, 34.18016, 34.28999, 34.39976, 34.50946, 
    34.61909, 34.72866, 34.83817, 34.9476, 35.05697, 35.16628, 35.27551, 
    35.38468, 35.49378, 35.60281, 35.71177, 35.82066, 35.92949, 36.03824, 
    36.14692, 36.25553, 36.36407, 36.47255, 36.58094, 36.68927, 36.79753, 
    36.90571, 37.01382, 37.12186, 37.22982,
  -10.94865, -10.84836, -10.74797, -10.64749, -10.54692, -10.44626, -10.3455, 
    -10.24466, -10.14372, -10.04269, -9.941566, -9.840355, -9.739052, 
    -9.637657, -9.536173, -9.434597, -9.332931, -9.231174, -9.129327, 
    -9.02739, -8.925363, -8.823246, -8.72104, -8.618743, -8.516357, 
    -8.413882, -8.311318, -8.208666, -8.105924, -8.003094, -7.900175, 
    -7.797167, -7.694072, -7.590889, -7.487617, -7.384259, -7.280813, 
    -7.177279, -7.073658, -6.969951, -6.866157, -6.762276, -6.658309, 
    -6.554255, -6.450116, -6.345891, -6.24158, -6.137184, -6.032702, 
    -5.928136, -5.823484, -5.718749, -5.613928, -5.509024, -5.404036, 
    -5.298964, -5.193808, -5.088569, -4.983246, -4.877841, -4.772354, 
    -4.666784, -4.561131, -4.455397, -4.349581, -4.243683, -4.137704, 
    -4.031644, -3.925504, -3.819282, -3.712981, -3.606599, -3.500138, 
    -3.393596, -3.286976, -3.180277, -3.073498, -2.966642, -2.859706, 
    -2.752693, -2.645602, -2.538434, -2.431189, -2.323866, -2.216467, 
    -2.108991, -2.00144, -1.893812, -1.786109, -1.67833, -1.570477, 
    -1.462549, -1.354546, -1.24647, -1.138319, -1.030095, -0.921798, 
    -0.8134278, -0.704985, -0.5964699, -0.4878827, -0.3792239, -0.2704936, 
    -0.1616923, -0.05282013, 0.05612245, 0.1651352, 0.2742177, 0.3833698, 
    0.492591, 0.601881, 0.7112396, 0.8206664, 0.930161, 1.039723, 1.149352, 
    1.259049, 1.368811, 1.47864, 1.588535, 1.698495, 1.80852, 1.91861, 
    2.028765, 2.138983, 2.249266, 2.359611, 2.47002, 2.580491, 2.691025, 
    2.80162, 2.912277, 3.022995, 3.133774, 3.244613, 3.355513, 3.466472, 
    3.57749, 3.688568, 3.799704, 3.910898, 4.02215, 4.133459, 4.244825, 
    4.356247, 4.467727, 4.579261, 4.690852, 4.802497, 4.914197, 5.025951, 
    5.137759, 5.24962, 5.361535, 5.473502, 5.585521, 5.697592, 5.809714, 
    5.921887, 6.034111, 6.146385, 6.258709, 6.371082, 6.483504, 6.595974, 
    6.708492, 6.821058, 6.933671, 7.046331, 7.159037, 7.271789, 7.384586, 
    7.497428, 7.610315, 7.723246, 7.836221, 7.949239, 8.0623, 8.175403, 
    8.288548, 8.401733, 8.514961, 8.628229, 8.741537, 8.854885, 8.968272, 
    9.081697, 9.195162, 9.308663, 9.422202, 9.535778, 9.649391, 9.76304, 
    9.876723, 9.990442, 10.1042, 10.21798, 10.33181, 10.44566, 10.55955, 
    10.67347, 10.78742, 10.9014, 11.01541, 11.12946, 11.24353, 11.35763, 
    11.47177, 11.58593, 11.70011, 11.81433, 11.92857, 12.04284, 12.15714, 
    12.27146, 12.3858, 12.50017, 12.61457, 12.72899, 12.84343, 12.95789, 
    13.07238, 13.18688, 13.30141, 13.41596, 13.53053, 13.64512, 13.75973, 
    13.87435, 13.989, 14.10366, 14.21834, 14.33304, 14.44775, 14.56248, 
    14.67722, 14.79198, 14.90675, 15.02154, 15.13633, 15.25115, 15.36597, 
    15.4808, 15.59565, 15.71051, 15.82537, 15.94025, 16.05514, 16.17003, 
    16.28493, 16.39984, 16.51476, 16.62968, 16.74461, 16.85955, 16.97449, 
    17.08943, 17.20438, 17.31933, 17.43429, 17.54925, 17.66421, 17.77917, 
    17.89413, 18.00909, 18.12406, 18.23902, 18.35398, 18.46894, 18.58389, 
    18.69885, 18.8138, 18.92875, 19.04369, 19.15863, 19.27357, 19.3885, 
    19.50342, 19.61834, 19.73324, 19.84814, 19.96304, 20.07792, 20.1928, 
    20.30766, 20.42252, 20.53736, 20.65219, 20.76702, 20.88183, 20.99662, 
    21.11141, 21.22618, 21.34093, 21.45567, 21.5704, 21.68511, 21.7998, 
    21.91448, 22.02914, 22.14378, 22.2584, 22.37301, 22.48759, 22.60216, 
    22.71671, 22.83123, 22.94573, 23.06022, 23.17468, 23.28911, 23.40353, 
    23.51792, 23.63229, 23.74663, 23.86094, 23.97523, 24.0895, 24.20374, 
    24.31795, 24.43213, 24.54629, 24.66042, 24.77452, 24.88858, 25.00262, 
    25.11663, 25.23061, 25.34456, 25.45847, 25.57235, 25.6862, 25.80002, 
    25.9138, 26.02755, 26.14126, 26.25494, 26.36858, 26.48219, 26.59576, 
    26.70929, 26.82279, 26.93625, 27.04967, 27.16305, 27.27639, 27.38969, 
    27.50295, 27.61617, 27.72935, 27.84249, 27.95559, 28.06864, 28.18165, 
    28.29462, 28.40755, 28.52042, 28.63326, 28.74605, 28.8588, 28.97149, 
    29.08415, 29.19675, 29.30931, 29.42182, 29.53428, 29.6467, 29.75906, 
    29.87138, 29.98364, 30.09586, 30.20802, 30.32014, 30.4322, 30.54421, 
    30.65617, 30.76808, 30.87993, 30.99173, 31.10348, 31.21517, 31.3268, 
    31.43839, 31.54991, 31.66138, 31.77279, 31.88415, 31.99545, 32.1067, 
    32.21788, 32.32901, 32.44007, 32.55108, 32.66203, 32.77292, 32.88375, 
    32.99452, 33.10523, 33.21588, 33.32647, 33.43699, 33.54745, 33.65785, 
    33.76818, 33.87846, 33.98866, 34.09881, 34.20889, 34.3189, 34.42885, 
    34.53874, 34.64856, 34.75831, 34.86799, 34.97761, 35.08716, 35.19665, 
    35.30606, 35.41541, 35.52469, 35.6339, 35.74304, 35.85211, 35.96112, 
    36.07005, 36.17891, 36.2877, 36.39642, 36.50507, 36.61364, 36.72215, 
    36.83057, 36.93893, 37.04722, 37.15543, 37.26357,
  -10.99701, -10.89658, -10.79605, -10.69544, -10.59472, -10.49392, 
    -10.39303, -10.29204, -10.19096, -10.08979, -9.988524, -9.88717, 
    -9.785724, -9.684186, -9.582557, -9.480837, -9.379026, -9.277124, 
    -9.175132, -9.07305, -8.970876, -8.868612, -8.766258, -8.663815, 
    -8.561281, -8.458658, -8.355946, -8.253143, -8.150252, -8.047272, 
    -7.944203, -7.841045, -7.737799, -7.634464, -7.531041, -7.42753, 
    -7.323932, -7.220245, -7.116471, -7.01261, -6.908661, -6.804626, 
    -6.700504, -6.596295, -6.492, -6.387619, -6.283151, -6.178598, -6.073959, 
    -5.969235, -5.864426, -5.759531, -5.654552, -5.549489, -5.444341, 
    -5.339108, -5.233792, -5.128393, -5.022909, -4.917343, -4.811693, 
    -4.70596, -4.600145, -4.494247, -4.388268, -4.282207, -4.176064, 
    -4.069839, -3.963533, -3.857146, -3.750679, -3.644131, -3.537503, 
    -3.430795, -3.324007, -3.21714, -3.110193, -3.003168, -2.896064, 
    -2.788882, -2.681621, -2.574283, -2.466867, -2.359374, -2.251803, 
    -2.144156, -2.036433, -1.928633, -1.820757, -1.712806, -1.604779, 
    -1.496678, -1.388501, -1.28025, -1.171925, -1.063526, -0.9550529, 
    -0.8465068, -0.7378878, -0.6291961, -0.5204321, -0.4115959, -0.302688, 
    -0.1937087, -0.08465826, 0.02446301, 0.1336548, 0.2429167, 0.3522485, 
    0.4616497, 0.5711202, 0.6806595, 0.7902674, 0.8999435, 1.009687, 
    1.119499, 1.229378, 1.339323, 1.449335, 1.559413, 1.669557, 1.779766, 
    1.890041, 2.00038, 2.110784, 2.221251, 2.331783, 2.442378, 2.553035, 
    2.663755, 2.774538, 2.885382, 2.996288, 3.107255, 3.218282, 3.32937, 
    3.440518, 3.551726, 3.662993, 3.774319, 3.885703, 3.997145, 4.108645, 
    4.220202, 4.331816, 4.443487, 4.555213, 4.666996, 4.778833, 4.890726, 
    5.002673, 5.114675, 5.226729, 5.338838, 5.450999, 5.563212, 5.675478, 
    5.787795, 5.900164, 6.012583, 6.125052, 6.237572, 6.350142, 6.462759, 
    6.575427, 6.688142, 6.800905, 6.913716, 7.026573, 7.139477, 7.252427, 
    7.365423, 7.478464, 7.59155, 7.70468, 7.817854, 7.931072, 8.044333, 
    8.157636, 8.270981, 8.384368, 8.497796, 8.611265, 8.724774, 8.838323, 
    8.951912, 9.065539, 9.179205, 9.292909, 9.406651, 9.52043, 9.634245, 
    9.748096, 9.861983, 9.975905, 10.08986, 10.20385, 10.31788, 10.43194, 
    10.54603, 10.66015, 10.77431, 10.8885, 11.00272, 11.11696, 11.23124, 
    11.34555, 11.45989, 11.57426, 11.68865, 11.80307, 11.91752, 12.032, 
    12.1465, 12.26103, 12.37558, 12.49016, 12.60476, 12.71938, 12.83403, 
    12.9487, 13.06339, 13.17811, 13.29284, 13.4076, 13.52238, 13.63718, 
    13.75199, 13.86683, 13.98168, 14.09655, 14.21144, 14.32634, 14.44127, 
    14.5562, 14.67115, 14.78612, 14.9011, 15.0161, 15.1311, 15.24613, 
    15.36116, 15.4762, 15.59126, 15.70632, 15.8214, 15.93649, 16.05158, 
    16.16669, 16.2818, 16.39692, 16.51204, 16.62718, 16.74232, 16.85746, 
    16.97261, 17.08777, 17.20293, 17.31809, 17.43325, 17.54842, 17.66359, 
    17.77876, 17.89394, 18.00911, 18.12428, 18.23945, 18.35463, 18.4698, 
    18.58496, 18.70013, 18.81529, 18.93045, 19.0456, 19.16075, 19.2759, 
    19.39104, 19.50617, 19.62129, 19.73641, 19.85152, 19.96663, 20.08172, 
    20.1968, 20.31188, 20.42694, 20.542, 20.65704, 20.77207, 20.88709, 
    21.00209, 21.11709, 21.23207, 21.34703, 21.46198, 21.57691, 21.69183, 
    21.80674, 21.92162, 22.03649, 22.15134, 22.26617, 22.38098, 22.49578, 
    22.61055, 22.72531, 22.84004, 22.95475, 23.06944, 23.18411, 23.29875, 
    23.41337, 23.52797, 23.64254, 23.75709, 23.87162, 23.98611, 24.10059, 
    24.21503, 24.32945, 24.44384, 24.5582, 24.67253, 24.78684, 24.90111, 
    25.01535, 25.12957, 25.24375, 25.3579, 25.47202, 25.58611, 25.70016, 
    25.81418, 25.92817, 26.04212, 26.15603, 26.26992, 26.38376, 26.49757, 
    26.61134, 26.72508, 26.83878, 26.95244, 27.06606, 27.17964, 27.29318, 
    27.40669, 27.52015, 27.63357, 27.74695, 27.86029, 27.97359, 28.08684, 
    28.20005, 28.31322, 28.42634, 28.53942, 28.65245, 28.76544, 28.87839, 
    28.99128, 29.10413, 29.21694, 29.32969, 29.4424, 29.55506, 29.66767, 
    29.78023, 29.89274, 30.0052, 30.11761, 30.22997, 30.34229, 30.45454, 
    30.56675, 30.6789, 30.791, 30.90305, 31.01504, 31.12698, 31.23886, 
    31.35069, 31.46246, 31.57418, 31.68584, 31.79745, 31.909, 32.02049, 
    32.13192, 32.24329, 32.35461, 32.46587, 32.57707, 32.68821, 32.79929, 
    32.9103, 33.02126, 33.13216, 33.24299, 33.35376, 33.46447, 33.57512, 
    33.68571, 33.79623, 33.90668, 34.01708, 34.12741, 34.23767, 34.34787, 
    34.458, 34.56807, 34.67807, 34.78801, 34.89788, 35.00768, 35.11741, 
    35.22707, 35.33667, 35.4462, 35.55566, 35.66505, 35.77437, 35.88362, 
    35.9928, 36.10191, 36.21095, 36.31992, 36.42882, 36.53764, 36.64639, 
    36.75507, 36.86368, 36.97222, 37.08068, 37.18906, 37.29738,
  -11.04545, -10.94487, -10.84421, -10.74345, -10.6426, -10.54166, -10.44062, 
    -10.33949, -10.23827, -10.13696, -10.03555, -9.934054, -9.832465, 
    -9.730783, -9.629011, -9.527146, -9.425191, -9.323144, -9.221006, 
    -9.118777, -9.016458, -8.914047, -8.811547, -8.708956, -8.606275, 
    -8.503503, -8.400641, -8.29769, -8.19465, -8.091519, -7.9883, -7.884992, 
    -7.781594, -7.678108, -7.574533, -7.47087, -7.367119, -7.263279, 
    -7.159352, -7.055336, -6.951234, -6.847044, -6.742766, -6.638402, 
    -6.533951, -6.429414, -6.32479, -6.22008, -6.115283, -6.010402, 
    -5.905434, -5.800381, -5.695243, -5.59002, -5.484712, -5.37932, 
    -5.273843, -5.168283, -5.062638, -4.956909, -4.851098, -4.745203, 
    -4.639225, -4.533164, -4.427021, -4.320795, -4.214487, -4.108098, 
    -4.001626, -3.895074, -3.788441, -3.681727, -3.574932, -3.468057, 
    -3.361101, -3.254066, -3.146952, -3.039758, -2.932485, -2.825133, 
    -2.717703, -2.610194, -2.502608, -2.394943, -2.287202, -2.179383, 
    -2.071488, -1.963516, -1.855467, -1.747342, -1.639142, -1.530867, 
    -1.422516, -1.31409, -1.20559, -1.097016, -0.9883671, -0.879645, 
    -0.7708496, -0.6619811, -0.5530399, -0.4440263, -0.3349406, -0.225783, 
    -0.116554, -0.007253821, 0.1021172, 0.2115587, 0.3210705, 0.4306521, 
    0.5403032, 0.6500235, 0.7598128, 0.8696705, 0.9795964, 1.08959, 1.199652, 
    1.30978, 1.419976, 1.530237, 1.640565, 1.750959, 1.861418, 1.971943, 
    2.082532, 2.193185, 2.303902, 2.414683, 2.525528, 2.636435, 2.747405, 
    2.858437, 2.96953, 3.080685, 3.191902, 3.303179, 3.414516, 3.525913, 
    3.637369, 3.748885, 3.86046, 3.972093, 4.083784, 4.195532, 4.307338, 
    4.4192, 4.531119, 4.643094, 4.755125, 4.86721, 4.979351, 5.091545, 
    5.203794, 5.316096, 5.428452, 5.54086, 5.653321, 5.765833, 5.878397, 
    5.991013, 6.103678, 6.216394, 6.32916, 6.441975, 6.554839, 6.667752, 
    6.780713, 6.893721, 7.006777, 7.119879, 7.233027, 7.346222, 7.459463, 
    7.572748, 7.686077, 7.799451, 7.912868, 8.02633, 8.139833, 8.253379, 
    8.366967, 8.480597, 8.594267, 8.707977, 8.821729, 8.935519, 9.049349, 
    9.163217, 9.277123, 9.391068, 9.50505, 9.619068, 9.733123, 9.847214, 
    9.96134, 10.0755, 10.1897, 10.30393, 10.41819, 10.53249, 10.64681, 
    10.76118, 10.87557, 10.98999, 11.10445, 11.21893, 11.33345, 11.44799, 
    11.56256, 11.67716, 11.79179, 11.90645, 12.02113, 12.13584, 12.25057, 
    12.36533, 12.48011, 12.59492, 12.70976, 12.82461, 12.93949, 13.05439, 
    13.16932, 13.28426, 13.39923, 13.51421, 13.62922, 13.74424, 13.85929, 
    13.97435, 14.08943, 14.20452, 14.31964, 14.43477, 14.54991, 14.66508, 
    14.78025, 14.89544, 15.01065, 15.12586, 15.24109, 15.35634, 15.47159, 
    15.58686, 15.70213, 15.81742, 15.93272, 16.04802, 16.16334, 16.27866, 
    16.39399, 16.50933, 16.62467, 16.74002, 16.85538, 16.97074, 17.0861, 
    17.20147, 17.31684, 17.43222, 17.5476, 17.66298, 17.77836, 17.89374, 
    18.00913, 18.12451, 18.23989, 18.35527, 18.47065, 18.58603, 18.70141, 
    18.81678, 18.93215, 19.04751, 19.16287, 19.27823, 19.39358, 19.50892, 
    19.62426, 19.73958, 19.85491, 19.97022, 20.08552, 20.20082, 20.3161, 
    20.43138, 20.54664, 20.66189, 20.77713, 20.89236, 21.00758, 21.12278, 
    21.23797, 21.35314, 21.4683, 21.58344, 21.69857, 21.81368, 21.92878, 
    22.04386, 22.15891, 22.27395, 22.38898, 22.50398, 22.61896, 22.73392, 
    22.84887, 22.96379, 23.07868, 23.19356, 23.30841, 23.42324, 23.53804, 
    23.65282, 23.76758, 23.88231, 23.99701, 24.11169, 24.22635, 24.34097, 
    24.45556, 24.57013, 24.68467, 24.79918, 24.91366, 25.02811, 25.14253, 
    25.25692, 25.37127, 25.4856, 25.59989, 25.71415, 25.82837, 25.94256, 
    26.05672, 26.17084, 26.28492, 26.39897, 26.51298, 26.62696, 26.7409, 
    26.8548, 26.96866, 27.08248, 27.19627, 27.31001, 27.42372, 27.53738, 
    27.651, 27.76459, 27.87812, 27.99162, 28.10508, 28.21848, 28.33185, 
    28.44518, 28.55845, 28.67169, 28.78487, 28.89802, 29.01111, 29.12416, 
    29.23716, 29.35011, 29.46302, 29.57587, 29.68868, 29.80144, 29.91415, 
    30.0268, 30.13941, 30.25197, 30.36447, 30.47692, 30.58932, 30.70167, 
    30.81396, 30.92621, 31.03839, 31.15052, 31.2626, 31.37462, 31.48659, 
    31.5985, 31.71035, 31.82215, 31.93389, 32.04557, 32.15719, 32.26876, 
    32.38026, 32.49171, 32.6031, 32.71443, 32.8257, 32.9369, 33.04805, 
    33.15913, 33.27015, 33.38111, 33.49201, 33.60284, 33.71362, 33.82432, 
    33.93497, 34.04554, 34.15606, 34.26651, 34.37689, 34.48721, 34.59746, 
    34.70765, 34.81776, 34.92781, 35.0378, 35.14771, 35.25756, 35.36734, 
    35.47705, 35.58669, 35.69626, 35.80576, 35.91519, 36.02455, 36.13384, 
    36.24305, 36.3522, 36.46128, 36.57028, 36.67921, 36.78806, 36.89685, 
    37.00556, 37.1142, 37.22276, 37.33125,
  -11.09395, -10.99324, -10.89244, -10.79154, -10.69055, -10.58946, 
    -10.48829, -10.38702, -10.28565, -10.1842, -10.08265, -9.981009, 
    -9.879277, -9.777452, -9.675535, -9.573526, -9.471426, -9.369234, 
    -9.266951, -9.164577, -9.06211, -8.959553, -8.856905, -8.754167, 
    -8.651337, -8.548417, -8.445407, -8.342307, -8.239117, -8.135837, 
    -8.032467, -7.929008, -7.825459, -7.721821, -7.618094, -7.514279, 
    -7.410375, -7.306382, -7.202301, -7.098132, -6.993875, -6.88953, 
    -6.785098, -6.680578, -6.575971, -6.471277, -6.366497, -6.261629, 
    -6.156676, -6.051636, -5.94651, -5.841298, -5.736001, -5.630619, 
    -5.525151, -5.419598, -5.313961, -5.208239, -5.102433, -4.996542, 
    -4.890568, -4.784511, -4.67837, -4.572145, -4.465838, -4.359448, 
    -4.252976, -4.146422, -4.039785, -3.933067, -3.826268, -3.719387, 
    -3.612425, -3.505383, -3.39826, -3.291057, -3.183774, -3.076411, 
    -2.968969, -2.861447, -2.753847, -2.646168, -2.538411, -2.430576, 
    -2.322663, -2.214672, -2.106604, -1.99846, -1.890238, -1.78194, 
    -1.673566, -1.565117, -1.456591, -1.347991, -1.239316, -1.130565, 
    -1.021741, -0.9128428, -0.8038707, -0.6948252, -0.5857067, -0.4765153, 
    -0.3672515, -0.2579155, -0.1485077, -0.0390284, 0.07052212, 0.1801435, 
    0.2898355, 0.3995976, 0.5094296, 0.6193312, 0.729302, 0.8393417, 0.94945, 
    1.059626, 1.169871, 1.280183, 1.390562, 1.501007, 1.61152, 1.722098, 
    1.832742, 1.943452, 2.054227, 2.165066, 2.27597, 2.386937, 2.497968, 
    2.609063, 2.72022, 2.83144, 2.942722, 3.054066, 3.165471, 3.276937, 
    3.388463, 3.500051, 3.611697, 3.723403, 3.835169, 3.946992, 4.058875, 
    4.170815, 4.282812, 4.394867, 4.506979, 4.619146, 4.731369, 4.843648, 
    4.955983, 5.068371, 5.180814, 5.293311, 5.405861, 5.518465, 5.631121, 
    5.743829, 5.856589, 5.9694, 6.082262, 6.195175, 6.308137, 6.42115, 
    6.534211, 6.647322, 6.76048, 6.873687, 6.986941, 7.100242, 7.21359, 
    7.326983, 7.440423, 7.553908, 7.667438, 7.781012, 7.894629, 8.008291, 
    8.121995, 8.235743, 8.349531, 8.463363, 8.577234, 8.691147, 8.8051, 
    8.919093, 9.033125, 9.147197, 9.261306, 9.375454, 9.489638, 9.603861, 
    9.71812, 9.832415, 9.946745, 10.06111, 10.17551, 10.28994, 10.40441, 
    10.51891, 10.63345, 10.74801, 10.86261, 10.97724, 11.0919, 11.20659, 
    11.32131, 11.43606, 11.55084, 11.66565, 11.78049, 11.89535, 12.01024, 
    12.12515, 12.2401, 12.35506, 12.47005, 12.58507, 12.70011, 12.81518, 
    12.93026, 13.04537, 13.1605, 13.27566, 13.39083, 13.50603, 13.62124, 
    13.73647, 13.85173, 13.967, 14.08229, 14.19759, 14.31292, 14.42826, 
    14.54361, 14.65898, 14.77437, 14.88977, 15.00519, 15.12061, 15.23605, 
    15.35151, 15.46697, 15.58245, 15.69793, 15.81343, 15.92894, 16.04445, 
    16.15998, 16.27551, 16.39105, 16.5066, 16.62215, 16.73771, 16.85328, 
    16.96885, 17.08443, 17.20001, 17.31559, 17.43118, 17.54677, 17.66236, 
    17.77795, 17.89355, 18.00914, 18.12474, 18.24033, 18.35592, 18.47152, 
    18.5871, 18.70269, 18.81827, 18.93385, 19.04943, 19.165, 19.28057, 
    19.39612, 19.51168, 19.62723, 19.74277, 19.8583, 19.97382, 20.08933, 
    20.20484, 20.32034, 20.43582, 20.55129, 20.66676, 20.78221, 20.89765, 
    21.01307, 21.12848, 21.24388, 21.35927, 21.47464, 21.58999, 21.70533, 
    21.82065, 21.93595, 22.05124, 22.16651, 22.28176, 22.39699, 22.5122, 
    22.62739, 22.74256, 22.85771, 22.97284, 23.08794, 23.20303, 23.31809, 
    23.43312, 23.54814, 23.66313, 23.77809, 23.89303, 24.00794, 24.12282, 
    24.23768, 24.35251, 24.46732, 24.58209, 24.69683, 24.81155, 24.92624, 
    25.04089, 25.15552, 25.27011, 25.38467, 25.4992, 25.6137, 25.72816, 
    25.84259, 25.95698, 26.07134, 26.18567, 26.29996, 26.41421, 26.52843, 
    26.6426, 26.75675, 26.87085, 26.98491, 27.09894, 27.21293, 27.32688, 
    27.44078, 27.55465, 27.66847, 27.78225, 27.89599, 28.00969, 28.12335, 
    28.23696, 28.35052, 28.46405, 28.57752, 28.69096, 28.80434, 28.91768, 
    29.03098, 29.14422, 29.25742, 29.37057, 29.48368, 29.59673, 29.70973, 
    29.82269, 29.93559, 30.04845, 30.16125, 30.274, 30.3867, 30.49935, 
    30.61195, 30.72449, 30.83698, 30.94941, 31.06179, 31.17412, 31.28639, 
    31.3986, 31.51076, 31.62286, 31.73491, 31.8469, 31.95883, 32.0707, 
    32.18251, 32.29427, 32.40597, 32.5176, 32.62918, 32.7407, 32.85216, 
    32.96355, 33.07489, 33.18616, 33.29737, 33.40852, 33.5196, 33.63062, 
    33.74158, 33.85247, 33.9633, 34.07407, 34.18476, 34.2954, 34.40597, 
    34.51647, 34.6269, 34.73727, 34.84757, 34.95781, 35.06797, 35.17807, 
    35.2881, 35.39806, 35.50795, 35.61777, 35.72752, 35.8372, 35.94681, 
    36.05635, 36.16582, 36.27522, 36.38454, 36.49379, 36.60297, 36.71208, 
    36.82111, 36.93007, 37.03896, 37.14777, 37.25651, 37.36517,
  -11.14253, -11.04168, -10.94073, -10.83969, -10.73856, -10.63734, 
    -10.53602, -10.43461, -10.33311, -10.23151, -10.12982, -10.02804, 
    -9.92616, -9.824191, -9.722131, -9.619977, -9.517733, -9.415395, 
    -9.312966, -9.210445, -9.107833, -9.005129, -8.902333, -8.799447, 
    -8.69647, -8.593402, -8.490243, -8.386993, -8.283653, -8.180223, 
    -8.076703, -7.973093, -7.869393, -7.765604, -7.661725, -7.557757, 
    -7.4537, -7.349554, -7.245319, -7.140996, -7.036585, -6.932085, 
    -6.827497, -6.722822, -6.618059, -6.513209, -6.408271, -6.303247, 
    -6.198135, -6.092937, -5.987653, -5.882283, -5.776826, -5.671284, 
    -5.565657, -5.459943, -5.354145, -5.248262, -5.142294, -5.036242, 
    -4.930106, -4.823885, -4.717581, -4.611193, -4.504722, -4.398168, 
    -4.291531, -4.184812, -4.07801, -3.971126, -3.86416, -3.757112, 
    -3.649983, -3.542773, -3.435483, -3.328111, -3.220659, -3.113128, 
    -3.005516, -2.897825, -2.790055, -2.682205, -2.574277, -2.466271, 
    -2.358186, -2.250023, -2.141783, -2.033466, -1.925071, -1.8166, 
    -1.708052, -1.599428, -1.490728, -1.381952, -1.273102, -1.164176, 
    -1.055175, -0.9461005, -0.8369516, -0.7277288, -0.6184327, -0.5090634, 
    -0.3996213, -0.2901067, -0.1805198, -0.0708611, 0.03886915, 0.1486706, 
    0.258543, 0.368486, 0.4784991, 0.5885822, 0.6987349, 0.8089568, 
    0.9192476, 1.029607, 1.140034, 1.25053, 1.361093, 1.471723, 1.58242, 
    1.693183, 1.804012, 1.914908, 2.025868, 2.136894, 2.247984, 2.359138, 
    2.470357, 2.581639, 2.692984, 2.804392, 2.915863, 3.027395, 3.13899, 
    3.250645, 3.362361, 3.474138, 3.585976, 3.697872, 3.809829, 3.921844, 
    4.033918, 4.14605, 4.25824, 4.370487, 4.482791, 4.595151, 4.707569, 
    4.820041, 4.93257, 5.045152, 5.15779, 5.270482, 5.383227, 5.496026, 
    5.608877, 5.721781, 5.834737, 5.947745, 6.060804, 6.173913, 6.287074, 
    6.400283, 6.513543, 6.626851, 6.740208, 6.853613, 6.967066, 7.080566, 
    7.194113, 7.307707, 7.421346, 7.535031, 7.648761, 7.762535, 7.876354, 
    7.990216, 8.104122, 8.21807, 8.332061, 8.446094, 8.560168, 8.674283, 
    8.788439, 8.902635, 9.01687, 9.131144, 9.245457, 9.359808, 9.474196, 
    9.588623, 9.703086, 9.817585, 9.93212, 10.04669, 10.16129, 10.27594, 
    10.39061, 10.50531, 10.62006, 10.73483, 10.84963, 10.96447, 11.07933, 
    11.19423, 11.30916, 11.42412, 11.5391, 11.65412, 11.76916, 11.88423, 
    11.99932, 12.11445, 12.2296, 12.34477, 12.45997, 12.5752, 12.69045, 
    12.80572, 12.92102, 13.03633, 13.15168, 13.26704, 13.38242, 13.49782, 
    13.61325, 13.72869, 13.84415, 13.95963, 14.07513, 14.19065, 14.30618, 
    14.42173, 14.5373, 14.65288, 14.76848, 14.88409, 14.99971, 15.11535, 
    15.231, 15.34667, 15.46234, 15.57803, 15.69373, 15.80943, 15.92515, 
    16.04088, 16.15661, 16.27236, 16.38811, 16.50387, 16.61963, 16.73541, 
    16.85118, 16.96697, 17.08275, 17.19855, 17.31434, 17.43014, 17.54594, 
    17.66174, 17.77755, 17.89335, 18.00916, 18.12497, 18.24077, 18.35658, 
    18.47238, 18.58818, 18.70398, 18.81977, 18.93556, 19.05135, 19.16713, 
    19.28291, 19.39868, 19.51444, 19.6302, 19.74595, 19.86169, 19.97743, 
    20.09315, 20.20887, 20.32458, 20.44027, 20.55596, 20.67163, 20.78729, 
    20.90294, 21.01858, 21.1342, 21.24981, 21.3654, 21.48098, 21.59655, 
    21.71209, 21.82762, 21.94314, 22.05863, 22.17411, 22.28957, 22.40501, 
    22.52043, 22.63583, 22.75121, 22.86657, 22.98191, 23.09722, 23.21251, 
    23.32778, 23.44303, 23.55825, 23.67345, 23.78862, 23.90376, 24.01888, 
    24.13398, 24.24904, 24.36408, 24.47909, 24.59407, 24.70902, 24.82395, 
    24.93884, 25.0537, 25.16853, 25.28333, 25.3981, 25.51283, 25.62753, 
    25.7422, 25.85684, 25.97144, 26.086, 26.20053, 26.31502, 26.42948, 
    26.5439, 26.65828, 26.77263, 26.88693, 27.0012, 27.11543, 27.22962, 
    27.34377, 27.45788, 27.57195, 27.68597, 27.79996, 27.9139, 28.0278, 
    28.14165, 28.25546, 28.36923, 28.48296, 28.59663, 28.71027, 28.82385, 
    28.93739, 29.05088, 29.16433, 29.27773, 29.39108, 29.50438, 29.61763, 
    29.73083, 29.84398, 29.95708, 30.07014, 30.18313, 30.29608, 30.40898, 
    30.52182, 30.63461, 30.74735, 30.86003, 30.97266, 31.08523, 31.19775, 
    31.31022, 31.42263, 31.53498, 31.64727, 31.75951, 31.87169, 31.98381, 
    32.09588, 32.20789, 32.31983, 32.43172, 32.54355, 32.65532, 32.76702, 
    32.87867, 32.99025, 33.10178, 33.21323, 33.32463, 33.43597, 33.54724, 
    33.65845, 33.76959, 33.88067, 33.99169, 34.10264, 34.21352, 34.32434, 
    34.4351, 34.54578, 34.6564, 34.76695, 34.87744, 34.98785, 35.0982, 
    35.20848, 35.3187, 35.42884, 35.53891, 35.64891, 35.75884, 35.8687, 
    35.97849, 36.08821, 36.19786, 36.30743, 36.41694, 36.52637, 36.63573, 
    36.74501, 36.85422, 36.96336, 37.07242, 37.18141, 37.29033, 37.39916,
  -11.19117, -11.09018, -10.9891, -10.88792, -10.78665, -10.68529, -10.58383, 
    -10.48228, -10.38063, -10.27889, -10.17706, -10.07513, -9.973113, 
    -9.871001, -9.768797, -9.666499, -9.564109, -9.461627, -9.359052, 
    -9.256385, -9.153626, -9.050776, -8.947833, -8.844799, -8.741673, 
    -8.638456, -8.535149, -8.43175, -8.32826, -8.22468, -8.12101, -8.017249, 
    -7.913397, -7.809456, -7.705426, -7.601305, -7.497095, -7.392796, 
    -7.288407, -7.18393, -7.079364, -6.97471, -6.869967, -6.765135, 
    -6.660216, -6.55521, -6.450115, -6.344933, -6.239664, -6.134308, 
    -6.028865, -5.923336, -5.81772, -5.712018, -5.60623, -5.500357, 
    -5.394397, -5.288353, -5.182223, -5.076009, -4.96971, -4.863327, 
    -4.756859, -4.650308, -4.543673, -4.436954, -4.330152, -4.223267, 
    -4.1163, -4.009249, -3.902117, -3.794903, -3.687607, -3.580229, -3.47277, 
    -3.365231, -3.25761, -3.149909, -3.042128, -2.934267, -2.826326, 
    -2.718306, -2.610207, -2.502029, -2.393772, -2.285438, -2.177025, 
    -2.068534, -1.959966, -1.851321, -1.742599, -1.633801, -1.524926, 
    -1.415975, -1.306949, -1.197847, -1.08867, -0.9794185, -0.8700925, 
    -0.7606924, -0.6512184, -0.5416709, -0.4320503, -0.3223567, -0.2125906, 
    -0.1027523, 0.007157928, 0.1171397, 0.2271928, 0.3373168, 0.4475114, 
    0.5577762, 0.668111, 0.7785153, 0.8889889, 0.9995313, 1.110142, 1.220822, 
    1.331569, 1.442383, 1.553265, 1.664214, 1.775229, 1.88631, 1.997456, 
    2.108668, 2.219945, 2.331287, 2.442693, 2.554163, 2.665696, 2.777293, 
    2.888952, 3.000674, 3.112458, 3.224303, 3.336209, 3.448177, 3.560205, 
    3.672292, 3.78444, 3.896647, 4.008913, 4.121237, 4.233619, 4.346059, 
    4.458556, 4.571111, 4.683721, 4.796388, 4.90911, 5.021888, 5.13472, 
    5.247607, 5.360548, 5.473542, 5.58659, 5.69969, 5.812843, 5.926047, 
    6.039303, 6.15261, 6.265968, 6.379375, 6.492833, 6.60634, 6.719895, 
    6.833499, 6.947152, 7.060851, 7.174598, 7.288391, 7.402231, 7.516116, 
    7.630046, 7.744022, 7.858042, 7.972106, 8.086213, 8.200363, 8.314556, 
    8.428791, 8.543067, 8.657385, 8.771744, 8.886143, 9.000581, 9.115059, 
    9.229575, 9.344131, 9.458724, 9.573354, 9.688022, 9.802726, 9.917465, 
    10.03224, 10.14705, 10.2619, 10.37678, 10.49169, 10.60663, 10.72161, 
    10.83662, 10.95167, 11.06674, 11.18184, 11.29698, 11.41214, 11.52734, 
    11.64256, 11.75781, 11.87309, 11.98839, 12.10372, 12.21908, 12.33446, 
    12.44987, 12.56531, 12.68076, 12.79625, 12.91175, 13.02728, 13.14283, 
    13.2584, 13.37399, 13.48961, 13.60524, 13.72089, 13.83657, 13.95226, 
    14.06796, 14.18369, 14.29944, 14.4152, 14.53097, 14.64676, 14.76257, 
    14.87839, 14.99423, 15.11008, 15.22594, 15.34181, 15.4577, 15.5736, 
    15.68951, 15.80543, 15.92136, 16.03729, 16.15324, 16.2692, 16.38516, 
    16.50113, 16.61711, 16.73309, 16.84908, 16.96508, 17.08108, 17.19708, 
    17.31309, 17.4291, 17.54511, 17.66113, 17.77714, 17.89316, 18.00918, 
    18.12519, 18.24121, 18.35723, 18.47324, 18.58925, 18.70526, 18.82127, 
    18.93727, 19.05327, 19.16927, 19.28525, 19.40124, 19.51721, 19.63318, 
    19.74915, 19.8651, 19.98104, 20.09698, 20.21291, 20.32883, 20.44473, 
    20.56063, 20.67652, 20.79239, 20.90825, 21.0241, 21.13993, 21.25575, 
    21.37155, 21.48734, 21.60312, 21.71887, 21.83462, 21.95034, 22.06605, 
    22.18173, 22.2974, 22.41305, 22.52868, 22.64429, 22.75988, 22.87545, 
    22.991, 23.10652, 23.22202, 23.3375, 23.45296, 23.56838, 23.68379, 
    23.79917, 23.91452, 24.02985, 24.14515, 24.26043, 24.37567, 24.49089, 
    24.60608, 24.72124, 24.83637, 24.95147, 25.06653, 25.18157, 25.29658, 
    25.41155, 25.52649, 25.6414, 25.75627, 25.87111, 25.98592, 26.10069, 
    26.21542, 26.33012, 26.44478, 26.55941, 26.67399, 26.78854, 26.90305, 
    27.01752, 27.13196, 27.24635, 27.3607, 27.47501, 27.58928, 27.70351, 
    27.8177, 27.93184, 28.04594, 28.16, 28.27401, 28.38798, 28.5019, 
    28.61578, 28.72961, 28.8434, 28.95714, 29.07083, 29.18447, 29.29807, 
    29.41162, 29.52512, 29.63857, 29.75197, 29.86532, 29.97861, 30.09186, 
    30.20506, 30.3182, 30.4313, 30.54433, 30.65732, 30.77025, 30.88313, 
    30.99596, 31.10872, 31.22144, 31.3341, 31.4467, 31.55924, 31.67173, 
    31.78416, 31.89654, 32.00885, 32.12111, 32.2333, 32.34544, 32.45752, 
    32.56954, 32.6815, 32.79339, 32.90523, 33.017, 33.12872, 33.24036, 
    33.35195, 33.46347, 33.57493, 33.68633, 33.79766, 33.90893, 34.02013, 
    34.13127, 34.24234, 34.35334, 34.46428, 34.57515, 34.68596, 34.79669, 
    34.90736, 35.01796, 35.12849, 35.23895, 35.34935, 35.45967, 35.56992, 
    35.68011, 35.79022, 35.90026, 36.01023, 36.12013, 36.22996, 36.33971, 
    36.44939, 36.55901, 36.66854, 36.778, 36.88739, 36.9967, 37.10595, 
    37.21511, 37.3242, 37.43322,
  -11.23989, -11.13876, -11.03754, -10.93622, -10.83481, -10.73331, 
    -10.63171, -10.53001, -10.42823, -10.32635, -10.22437, -10.1223, 
    -10.02014, -9.917883, -9.815535, -9.713092, -9.610558, -9.50793, 
    -9.40521, -9.302396, -9.199491, -9.096493, -8.993403, -8.890222, 
    -8.786948, -8.683582, -8.580126, -8.476578, -8.372938, -8.269208, 
    -8.165387, -8.061475, -7.957472, -7.853379, -7.749196, -7.644923, 
    -7.54056, -7.436108, -7.331565, -7.226933, -7.122213, -7.017404, 
    -6.912505, -6.807518, -6.702443, -6.597279, -6.492028, -6.386688, 
    -6.281261, -6.175747, -6.070146, -5.964457, -5.858682, -5.75282, 
    -5.646872, -5.540838, -5.434717, -5.328511, -5.22222, -5.115843, 
    -5.009382, -4.902835, -4.796204, -4.689489, -4.58269, -4.475806, 
    -4.368839, -4.261789, -4.154655, -4.047439, -3.94014, -3.832759, 
    -3.725296, -3.61775, -3.510123, -3.402415, -3.294626, -3.186755, 
    -3.078804, -2.970773, -2.862662, -2.754471, -2.6462, -2.537851, 
    -2.429422, -2.320915, -2.212329, -2.103665, -1.994924, -1.886105, 
    -1.777208, -1.668235, -1.559186, -1.450059, -1.340857, -1.231579, 
    -1.122226, -1.012797, -0.9032939, -0.7937161, -0.6840641, -0.5743383, 
    -0.4645388, -0.3546661, -0.2447206, -0.1347024, -0.02461194, 0.08555045, 
    0.1957844, 0.3060897, 0.4164659, 0.5269127, 0.6374299, 0.7480169, 
    0.8586735, 0.9693994, 1.080194, 1.191057, 1.301989, 1.412988, 1.524055, 
    1.635189, 1.74639, 1.857657, 1.96899, 2.080389, 2.191854, 2.303383, 
    2.414977, 2.526634, 2.638356, 2.750142, 2.86199, 2.973901, 3.085875, 
    3.19791, 3.310007, 3.422165, 3.534384, 3.646663, 3.759002, 3.871401, 
    3.983859, 4.096375, 4.208951, 4.321584, 4.434275, 4.547022, 4.659827, 
    4.772688, 4.885605, 4.998578, 5.111605, 5.224688, 5.337824, 5.451015, 
    5.564259, 5.677556, 5.790905, 5.904307, 6.01776, 6.131265, 6.24482, 
    6.358426, 6.472082, 6.585788, 6.699543, 6.813346, 6.927197, 7.041097, 
    7.155044, 7.269037, 7.383077, 7.497163, 7.611295, 7.725471, 7.839693, 
    7.953958, 8.068267, 8.18262, 8.297015, 8.411452, 8.525932, 8.640452, 
    8.755014, 8.869617, 8.98426, 9.098941, 9.213662, 9.328422, 9.443219, 
    9.558054, 9.672927, 9.787836, 9.902781, 10.01776, 10.13278, 10.24783, 
    10.36291, 10.47803, 10.59319, 10.70837, 10.82359, 10.93884, 11.05412, 
    11.16943, 11.28477, 11.40014, 11.51554, 11.63097, 11.74643, 11.86192, 
    11.97743, 12.09297, 12.20854, 12.32413, 12.43975, 12.55539, 12.67106, 
    12.78675, 12.90247, 13.0182, 13.13396, 13.24974, 13.36555, 13.48137, 
    13.59721, 13.71308, 13.82896, 13.94486, 14.06078, 14.17672, 14.29267, 
    14.40864, 14.52463, 14.64064, 14.75665, 14.87269, 14.98873, 15.10479, 
    15.22087, 15.33695, 15.45305, 15.56916, 15.68528, 15.80141, 15.91755, 
    16.0337, 16.14986, 16.26603, 16.38221, 16.49839, 16.61458, 16.73078, 
    16.84698, 16.96318, 17.0794, 17.19561, 17.31183, 17.42805, 17.54428, 
    17.66051, 17.77673, 17.89296, 18.00919, 18.12542, 18.24165, 18.35788, 
    18.47411, 18.59033, 18.70655, 18.82277, 18.93899, 19.0552, 19.1714, 
    19.28761, 19.4038, 19.51999, 19.63617, 19.75234, 19.86851, 19.98467, 
    20.10082, 20.21696, 20.33309, 20.44921, 20.56531, 20.68141, 20.79749, 
    20.91357, 21.02962, 21.14567, 21.2617, 21.37772, 21.49372, 21.6097, 
    21.72567, 21.84162, 21.95756, 22.07347, 22.18937, 22.30525, 22.42111, 
    22.53695, 22.65277, 22.76857, 22.88435, 23.00011, 23.11584, 23.23155, 
    23.34724, 23.4629, 23.57854, 23.69415, 23.80974, 23.92531, 24.04084, 
    24.15635, 24.27183, 24.38729, 24.50271, 24.61811, 24.73348, 24.84881, 
    24.96412, 25.0794, 25.19464, 25.30985, 25.42503, 25.54018, 25.65529, 
    25.77037, 25.88542, 26.00043, 26.1154, 26.23034, 26.34525, 26.46011, 
    26.57494, 26.68973, 26.80449, 26.9192, 27.03388, 27.14851, 27.26311, 
    27.37766, 27.49218, 27.60665, 27.72108, 27.83547, 27.94982, 28.06412, 
    28.17838, 28.29259, 28.40676, 28.52089, 28.63497, 28.749, 28.86298, 
    28.97692, 29.09081, 29.20466, 29.31845, 29.4322, 29.5459, 29.65955, 
    29.77315, 29.88669, 30.00019, 30.11364, 30.22703, 30.34037, 30.45366, 
    30.56689, 30.68008, 30.7932, 30.90628, 31.0193, 31.13226, 31.24517, 
    31.35802, 31.47082, 31.58356, 31.69624, 31.80886, 31.92143, 32.03394, 
    32.14638, 32.25877, 32.3711, 32.48337, 32.59558, 32.70773, 32.81982, 
    32.93184, 33.0438, 33.15571, 33.26754, 33.37932, 33.49103, 33.60268, 
    33.71426, 33.82578, 33.93724, 34.04863, 34.15995, 34.27121, 34.3824, 
    34.49352, 34.60458, 34.71556, 34.82648, 34.93734, 35.04812, 35.15884, 
    35.26948, 35.38006, 35.49056, 35.601, 35.71136, 35.82166, 35.93188, 
    36.04203, 36.15211, 36.26212, 36.37205, 36.48191, 36.5917, 36.70142, 
    36.81105, 36.92062, 37.03011, 37.13953, 37.24887, 37.35814, 37.46733,
  -11.28868, -11.18741, -11.08605, -10.9846, -10.88305, -10.7814, -10.67966, 
    -10.57782, -10.47589, -10.37387, -10.27175, -10.16954, -10.06724, 
    -9.964837, -9.862344, -9.759757, -9.657078, -9.554304, -9.451438, 
    -9.348479, -9.245427, -9.142282, -9.039045, -8.935716, -8.832294, 
    -8.72878, -8.625175, -8.521477, -8.417687, -8.313807, -8.209835, 
    -8.105772, -8.001617, -7.897373, -7.793038, -7.688612, -7.584096, 
    -7.47949, -7.374794, -7.270008, -7.165132, -7.060167, -6.955113, 
    -6.849971, -6.744739, -6.639419, -6.53401, -6.428513, -6.322928, 
    -6.217256, -6.111495, -6.005648, -5.899713, -5.793691, -5.687582, 
    -5.581387, -5.475106, -5.368738, -5.262285, -5.155746, -5.049121, 
    -4.942412, -4.835617, -4.728738, -4.621774, -4.514726, -4.407594, 
    -4.300378, -4.193079, -4.085696, -3.97823, -3.870682, -3.76305, 
    -3.655337, -3.547542, -3.439665, -3.331706, -3.223666, -3.115546, 
    -3.007344, -2.899062, -2.7907, -2.682258, -2.573736, -2.465136, 
    -2.356456, -2.247697, -2.13886, -2.029945, -1.920951, -1.811881, 
    -1.702732, -1.593507, -1.484205, -1.374827, -1.265373, -1.155843, 
    -1.046237, -0.9365563, -0.8268005, -0.7169703, -0.6070658, -0.4970873, 
    -0.3870353, -0.27691, -0.1667117, -0.05644082, 0.05390239, 0.1643176, 
    0.2748044, 0.3853625, 0.4959916, 0.6066913, 0.7174613, 0.8283012, 
    0.9392107, 1.050189, 1.161237, 1.272353, 1.383538, 1.49479, 1.60611, 
    1.717497, 1.82895, 1.94047, 2.052056, 2.163708, 2.275425, 2.387207, 
    2.499053, 2.610964, 2.722938, 2.834976, 2.947077, 3.05924, 3.171466, 
    3.283753, 3.396102, 3.508512, 3.620983, 3.733514, 3.846105, 3.958756, 
    4.071465, 4.184234, 4.29706, 4.409945, 4.522887, 4.635886, 4.748942, 
    4.862054, 4.975222, 5.088445, 5.201723, 5.315055, 5.428442, 5.541883, 
    5.655377, 5.768923, 5.882523, 5.996174, 6.109877, 6.22363, 6.337435, 
    6.45129, 6.565195, 6.679149, 6.793151, 6.907203, 7.021302, 7.135449, 
    7.249644, 7.363884, 7.478172, 7.592505, 7.706883, 7.821306, 7.935774, 
    8.050285, 8.164841, 8.279438, 8.394079, 8.508761, 8.623487, 8.738252, 
    8.853058, 8.967904, 9.08279, 9.197716, 9.31268, 9.427683, 9.542723, 
    9.657801, 9.772915, 9.888066, 10.00325, 10.11848, 10.23373, 10.34902, 
    10.46435, 10.57971, 10.6951, 10.81053, 10.92598, 11.04147, 11.15699, 
    11.27254, 11.38812, 11.50373, 11.61937, 11.73503, 11.85073, 11.96645, 
    12.0822, 12.19798, 12.31378, 12.42961, 12.54546, 12.66134, 12.77724, 
    12.89316, 13.00911, 13.12508, 13.24107, 13.35708, 13.47312, 13.58917, 
    13.70525, 13.82134, 13.93745, 14.05358, 14.16973, 14.2859, 14.40208, 
    14.51828, 14.63449, 14.75072, 14.86697, 14.98323, 15.0995, 15.21578, 
    15.33208, 15.44839, 15.56471, 15.68105, 15.79739, 15.91374, 16.03011, 
    16.14648, 16.26286, 16.37925, 16.49564, 16.61204, 16.72845, 16.84487, 
    16.96129, 17.07771, 17.19414, 17.31057, 17.42701, 17.54344, 17.65988, 
    17.77633, 17.89277, 18.00921, 18.12565, 18.24209, 18.35854, 18.47498, 
    18.59141, 18.70785, 18.82428, 18.94071, 19.05713, 19.17355, 19.28996, 
    19.40637, 19.52277, 19.63917, 19.75555, 19.87193, 19.9883, 20.10466, 
    20.22101, 20.33735, 20.45369, 20.57001, 20.68632, 20.80261, 20.91889, 
    21.03517, 21.15142, 21.26766, 21.38389, 21.5001, 21.6163, 21.73248, 
    21.84864, 21.96479, 22.08092, 22.19703, 22.31312, 22.42919, 22.54524, 
    22.66127, 22.77728, 22.89327, 23.00923, 23.12518, 23.2411, 23.357, 
    23.47287, 23.58872, 23.70454, 23.82034, 23.93611, 24.05186, 24.16757, 
    24.28326, 24.39893, 24.51456, 24.63017, 24.74574, 24.86128, 24.9768, 
    25.09228, 25.20773, 25.32315, 25.43854, 25.55389, 25.66921, 25.7845, 
    25.89975, 26.01497, 26.13015, 26.2453, 26.3604, 26.47548, 26.59051, 
    26.70551, 26.82047, 26.93538, 27.05027, 27.16511, 27.27991, 27.39466, 
    27.50938, 27.62406, 27.73869, 27.85328, 27.96783, 28.08234, 28.1968, 
    28.31121, 28.42558, 28.53991, 28.65419, 28.76842, 28.88261, 28.99675, 
    29.11084, 29.22489, 29.33888, 29.45283, 29.56672, 29.68057, 29.79437, 
    29.90811, 30.02181, 30.13545, 30.24904, 30.36258, 30.47606, 30.5895, 
    30.70288, 30.8162, 30.92947, 31.04268, 31.15584, 31.26895, 31.38199, 
    31.49498, 31.60792, 31.72079, 31.83361, 31.94637, 32.05907, 32.17171, 
    32.28429, 32.39681, 32.50927, 32.62167, 32.73401, 32.84629, 32.95851, 
    33.07066, 33.18275, 33.29478, 33.40674, 33.51864, 33.63048, 33.74225, 
    33.85396, 33.9656, 34.07718, 34.18869, 34.30013, 34.4115, 34.52281, 
    34.63406, 34.74523, 34.85633, 34.96737, 35.07834, 35.18924, 35.30006, 
    35.41082, 35.52151, 35.63213, 35.74268, 35.85315, 35.96356, 36.07389, 
    36.18415, 36.29433, 36.40445, 36.51449, 36.62445, 36.73435, 36.84417, 
    36.95391, 37.06358, 37.17317, 37.28269, 37.39214, 37.5015,
  -11.33754, -11.23614, -11.13464, -11.03304, -10.93135, -10.82957, 
    -10.72768, -10.62571, -10.52364, -10.42147, -10.31921, -10.21686, 
    -10.11441, -10.01186, -9.909226, -9.806495, -9.703671, -9.600752, 
    -9.49774, -9.394634, -9.291435, -9.188144, -9.08476, -8.981282, 
    -8.877711, -8.774049, -8.670295, -8.566447, -8.462508, -8.358478, 
    -8.254354, -8.150141, -8.045835, -7.941438, -7.83695, -7.732372, 
    -7.627702, -7.522943, -7.418093, -7.313152, -7.208122, -7.103002, 
    -6.997793, -6.892494, -6.787106, -6.681628, -6.576062, -6.470407, 
    -6.364665, -6.258833, -6.152915, -6.046907, -5.940813, -5.834631, 
    -5.728362, -5.622006, -5.515563, -5.409034, -5.302418, -5.195716, 
    -5.088929, -4.982056, -4.875098, -4.768054, -4.660926, -4.553713, 
    -4.446415, -4.339034, -4.231568, -4.124019, -4.016387, -3.90867, 
    -3.800872, -3.69299, -3.585026, -3.47698, -3.368852, -3.260643, 
    -3.152352, -3.04398, -2.935527, -2.826994, -2.71838, -2.609687, 
    -2.500913, -2.392061, -2.283129, -2.174118, -2.065029, -1.955861, 
    -1.846616, -1.737292, -1.627892, -1.518414, -1.40886, -1.299229, 
    -1.189521, -1.079738, -0.9698799, -0.859946, -0.7499372, -0.6398539, 
    -0.5296962, -0.4194646, -0.3091593, -0.1987807, -0.08832908, 0.02219518, 
    0.1327918, 0.2434604, 0.3542006, 0.4650122, 0.5758948, 0.686848, 
    0.7978715, 0.9089649, 1.020128, 1.13136, 1.242661, 1.354031, 1.465469, 
    1.576975, 1.688548, 1.800188, 1.911895, 2.023669, 2.135508, 2.247413, 
    2.359383, 2.471418, 2.583518, 2.695682, 2.807909, 2.9202, 3.032554, 
    3.14497, 3.257449, 3.369989, 3.482591, 3.595254, 3.707977, 3.82076, 
    3.933604, 4.046507, 4.159469, 4.272489, 4.385568, 4.498704, 4.611897, 
    4.725148, 4.838456, 4.951819, 5.065238, 5.178712, 5.292242, 5.405825, 
    5.519463, 5.633154, 5.746898, 5.860695, 5.974545, 6.088446, 6.202398, 
    6.316401, 6.430456, 6.54456, 6.658713, 6.772916, 6.887168, 7.001468, 
    7.115816, 7.230211, 7.344654, 7.459142, 7.573677, 7.688257, 7.802883, 
    7.917552, 8.032267, 8.147025, 8.261826, 8.37667, 8.491556, 8.606484, 
    8.721455, 8.836465, 8.951515, 9.066607, 9.181737, 9.296906, 9.412114, 
    9.52736, 9.642644, 9.757964, 9.873322, 9.988714, 10.10414, 10.21961, 
    10.33511, 10.45064, 10.56621, 10.68181, 10.79744, 10.9131, 11.0288, 
    11.14453, 11.26028, 11.37607, 11.49189, 11.60774, 11.72361, 11.83952, 
    11.95545, 12.07141, 12.18739, 12.3034, 12.41944, 12.5355, 12.65159, 
    12.7677, 12.88384, 12.99999, 13.11617, 13.23238, 13.3486, 13.46485, 
    13.58111, 13.6974, 13.8137, 13.93003, 14.04637, 14.16273, 14.27911, 
    14.3955, 14.51191, 14.62834, 14.74478, 14.86124, 14.97771, 15.09419, 
    15.21069, 15.3272, 15.44372, 15.56026, 15.6768, 15.79336, 15.90993, 
    16.0265, 16.14309, 16.25968, 16.37628, 16.49289, 16.6095, 16.72612, 
    16.84275, 16.95938, 17.07602, 17.19266, 17.30931, 17.42596, 17.54261, 
    17.65926, 17.77592, 17.89257, 18.00923, 18.12588, 18.24254, 18.35919, 
    18.47585, 18.59249, 18.70914, 18.82579, 18.94243, 19.05906, 19.1757, 
    19.29232, 19.40895, 19.52556, 19.64217, 19.75877, 19.87536, 19.99194, 
    20.10851, 20.22508, 20.34163, 20.45818, 20.57471, 20.69123, 20.80774, 
    20.92423, 21.04072, 21.15719, 21.27364, 21.39008, 21.5065, 21.62291, 
    21.7393, 21.85568, 21.97204, 22.08838, 22.2047, 22.321, 22.43728, 
    22.55354, 22.66978, 22.78601, 22.9022, 23.01838, 23.13453, 23.25067, 
    23.36677, 23.48286, 23.59892, 23.71495, 23.83096, 23.94694, 24.06289, 
    24.17882, 24.29472, 24.41059, 24.52643, 24.64225, 24.75803, 24.87378, 
    24.98951, 25.1052, 25.22086, 25.33648, 25.45208, 25.56764, 25.68317, 
    25.79866, 25.91412, 26.02954, 26.14493, 26.26028, 26.3756, 26.49087, 
    26.60611, 26.72131, 26.83648, 26.9516, 27.06669, 27.18173, 27.29674, 
    27.4117, 27.52662, 27.6415, 27.75634, 27.87113, 27.98588, 28.10059, 
    28.21525, 28.32987, 28.44444, 28.55897, 28.67345, 28.78789, 28.90228, 
    29.01661, 29.13091, 29.24515, 29.35935, 29.47349, 29.58759, 29.70164, 
    29.81563, 29.92957, 30.04347, 30.15731, 30.2711, 30.38483, 30.49852, 
    30.61215, 30.72572, 30.83924, 30.95271, 31.06612, 31.17947, 31.29277, 
    31.40601, 31.5192, 31.63232, 31.74539, 31.8584, 31.97136, 32.08425, 
    32.19708, 32.30986, 32.42257, 32.53522, 32.64782, 32.76035, 32.87282, 
    32.98522, 33.09757, 33.20985, 33.32206, 33.43422, 33.54631, 33.65833, 
    33.77029, 33.88219, 33.99401, 34.10578, 34.21748, 34.32911, 34.44067, 
    34.55216, 34.66359, 34.77495, 34.88624, 34.99746, 35.10861, 35.2197, 
    35.33071, 35.44165, 35.55252, 35.66332, 35.77405, 35.88471, 35.99529, 
    36.1058, 36.21625, 36.32661, 36.4369, 36.54713, 36.65727, 36.76735, 
    36.87734, 36.98726, 37.09711, 37.20688, 37.31657, 37.42619, 37.53574,
  -11.38648, -11.28494, -11.1833, -11.08156, -10.97973, -10.8778, -10.77578, 
    -10.67366, -10.57145, -10.46914, -10.36674, -10.26424, -10.16165, 
    -10.05896, -9.956182, -9.853306, -9.750336, -9.647271, -9.544114, 
    -9.440862, -9.337517, -9.234077, -9.130546, -9.02692, -8.923202, 
    -8.81939, -8.715487, -8.61149, -8.507401, -8.403219, -8.298946, 
    -8.194581, -8.090123, -7.985575, -7.880935, -7.776203, -7.671381, 
    -7.566467, -7.461463, -7.356368, -7.251183, -7.145908, -7.040543, 
    -6.935087, -6.829543, -6.723908, -6.618185, -6.512372, -6.406472, 
    -6.300482, -6.194404, -6.088237, -5.981983, -5.87564, -5.769211, 
    -5.662694, -5.556089, -5.449399, -5.34262, -5.235756, -5.128806, 
    -5.021769, -4.914647, -4.807439, -4.700146, -4.592768, -4.485305, 
    -4.377758, -4.270125, -4.16241, -4.05461, -3.946726, -3.83876, -3.73071, 
    -3.622577, -3.514362, -3.406065, -3.297685, -3.189224, -3.080682, 
    -2.972058, -2.863353, -2.754568, -2.645702, -2.536756, -2.42773, 
    -2.318625, -2.20944, -2.100177, -1.990835, -1.881414, -1.771916, 
    -1.662339, -1.552685, -1.442955, -1.333147, -1.223262, -1.113302, 
    -1.003265, -0.893153, -0.7829654, -0.672703, -0.5623658, -0.4519544, 
    -0.3414689, -0.2309097, -0.1202771, -0.009571564, 0.1012067, 0.2120573, 
    0.32298, 0.4339743, 0.54504, 0.6561767, 0.767384, 0.8786616, 0.9900092, 
    1.101426, 1.212913, 1.324468, 1.436092, 1.547784, 1.659544, 1.771371, 
    1.883265, 1.995226, 2.107254, 2.219347, 2.331506, 2.44373, 2.556019, 
    2.668372, 2.78079, 2.893271, 3.005816, 3.118423, 3.231093, 3.343825, 
    3.456618, 3.569473, 3.682389, 3.795366, 3.908402, 4.021499, 4.134654, 
    4.247869, 4.361142, 4.474473, 4.587862, 4.701308, 4.81481, 4.92837, 
    5.041985, 5.155656, 5.269382, 5.383162, 5.496997, 5.610886, 5.724828, 
    5.838824, 5.952871, 6.066971, 6.181123, 6.295326, 6.409579, 6.523883, 
    6.638237, 6.75264, 6.867093, 6.981594, 7.096143, 7.210739, 7.325383, 
    7.440073, 7.554811, 7.669593, 7.784421, 7.899294, 8.014212, 8.129172, 
    8.244178, 8.359225, 8.474316, 8.589448, 8.704622, 8.819838, 8.935093, 
    9.050389, 9.165725, 9.2811, 9.396514, 9.511966, 9.627455, 9.742982, 
    9.858546, 9.974146, 10.08978, 10.20545, 10.32116, 10.4369, 10.55267, 
    10.66848, 10.78432, 10.90019, 11.0161, 11.13204, 11.248, 11.364, 
    11.48003, 11.59608, 11.71217, 11.82828, 11.94442, 12.06059, 12.17679, 
    12.29301, 12.40926, 12.52553, 12.64183, 12.75815, 12.87449, 12.99086, 
    13.10725, 13.22367, 13.3401, 13.45656, 13.57304, 13.68953, 13.80605, 
    13.92259, 14.03914, 14.15571, 14.2723, 14.38891, 14.50553, 14.62217, 
    14.73882, 14.85549, 14.97218, 15.08887, 15.20559, 15.32231, 15.43904, 
    15.55579, 15.67255, 15.78932, 15.9061, 16.02289, 16.13968, 16.25649, 
    16.37331, 16.49013, 16.60696, 16.72379, 16.84063, 16.95748, 17.07433, 
    17.19118, 17.30804, 17.42491, 17.54177, 17.65864, 17.77551, 17.89237, 
    18.00924, 18.12611, 18.24298, 18.35985, 18.47672, 18.59358, 18.71044, 
    18.8273, 18.94415, 19.061, 19.17785, 19.29469, 19.41152, 19.52835, 
    19.64517, 19.76199, 19.87879, 19.99559, 20.11238, 20.22915, 20.34592, 
    20.46268, 20.57942, 20.69616, 20.81288, 20.92959, 21.04628, 21.16296, 
    21.27963, 21.39628, 21.51292, 21.62954, 21.74614, 21.86273, 21.9793, 
    22.09585, 22.21238, 22.3289, 22.44539, 22.56186, 22.67832, 22.79475, 
    22.91116, 23.02755, 23.14391, 23.26025, 23.37657, 23.49287, 23.60913, 
    23.72538, 23.8416, 23.95779, 24.07395, 24.19009, 24.3062, 24.42228, 
    24.53833, 24.65435, 24.77034, 24.88631, 25.00224, 25.11814, 25.234, 
    25.34984, 25.46564, 25.58141, 25.69715, 25.81285, 25.92851, 26.04414, 
    26.15974, 26.2753, 26.39082, 26.5063, 26.62175, 26.73715, 26.85252, 
    26.96785, 27.08314, 27.19839, 27.3136, 27.42877, 27.54389, 27.65898, 
    27.77402, 27.88902, 28.00397, 28.11888, 28.23375, 28.34857, 28.46334, 
    28.57807, 28.69275, 28.80739, 28.92198, 29.03652, 29.15101, 29.26546, 
    29.37986, 29.4942, 29.6085, 29.72274, 29.83694, 29.95108, 30.06517, 
    30.17921, 30.2932, 30.40713, 30.52101, 30.63484, 30.74861, 30.86233, 
    30.97599, 31.0896, 31.20315, 31.31664, 31.43008, 31.54346, 31.65678, 
    31.77004, 31.88325, 31.9964, 32.10948, 32.22251, 32.33548, 32.44838, 
    32.56123, 32.67401, 32.78674, 32.89939, 33.01199, 33.12453, 33.237, 
    33.3494, 33.46175, 33.57403, 33.68624, 33.79839, 33.91047, 34.02249, 
    34.13444, 34.24632, 34.35814, 34.46989, 34.58157, 34.69318, 34.80473, 
    34.9162, 35.02761, 35.13895, 35.25021, 35.36141, 35.47253, 35.58359, 
    35.69457, 35.80548, 35.91632, 36.02709, 36.13778, 36.2484, 36.35895, 
    36.46943, 36.57983, 36.69015, 36.8004, 36.91058, 37.02068, 37.1307, 
    37.24065, 37.35052, 37.46032, 37.57004,
  -11.43549, -11.33381, -11.23203, -11.13015, -11.02818, -10.92612, 
    -10.82395, -10.72169, -10.61934, -10.51689, -10.41434, -10.3117, 
    -10.20897, -10.10614, -10.00321, -9.900189, -9.797074, -9.693865, 
    -9.590561, -9.487163, -9.383671, -9.280085, -9.176405, -9.072632, 
    -8.968765, -8.864805, -8.760752, -8.656606, -8.552366, -8.448034, 
    -8.34361, -8.239094, -8.134484, -8.029784, -7.924991, -7.820107, 
    -7.715131, -7.610064, -7.504905, -7.399656, -7.294315, -7.188885, 
    -7.083364, -6.977752, -6.872051, -6.76626, -6.660379, -6.554409, 
    -6.448349, -6.3422, -6.235963, -6.129637, -6.023223, -5.91672, -5.81013, 
    -5.703452, -5.596685, -5.489832, -5.382892, -5.275865, -5.168751, 
    -5.061551, -4.954265, -4.846893, -4.739435, -4.631891, -4.524263, 
    -4.416549, -4.308751, -4.200868, -4.092901, -3.98485, -3.876715, 
    -3.768497, -3.660195, -3.551811, -3.443344, -3.334795, -3.226163, 
    -3.117449, -3.008654, -2.899778, -2.79082, -2.681782, -2.572663, 
    -2.463464, -2.354185, -2.244827, -2.135389, -2.025872, -1.916277, 
    -1.806602, -1.69685, -1.58702, -1.477112, -1.367128, -1.257066, 
    -1.146927, -1.036712, -0.9264217, -0.8160552, -0.7056134, -0.5950966, 
    -0.484505, -0.3738391, -0.2630991, -0.1522854, -0.04139822, 0.06956197, 
    0.1805949, 0.2917002, 0.4028775, 0.5141266, 0.625447, 0.7368384, 
    0.8483005, 0.9598328, 1.071435, 1.183107, 1.294848, 1.406658, 1.518537, 
    1.630484, 1.742498, 1.85458, 1.966729, 2.078945, 2.191227, 2.303575, 
    2.415988, 2.528466, 2.64101, 2.753618, 2.866289, 2.979025, 3.091823, 
    3.204685, 3.317609, 3.430595, 3.543642, 3.656751, 3.769921, 3.883151, 
    3.996441, 4.109791, 4.2232, 4.336668, 4.450193, 4.563778, 4.677419, 
    4.791118, 4.904874, 5.018685, 5.132553, 5.246476, 5.360454, 5.474487, 
    5.588574, 5.702714, 5.816908, 5.931155, 6.045454, 6.159805, 6.274207, 
    6.388661, 6.503165, 6.617719, 6.732323, 6.846977, 6.961679, 7.076429, 
    7.191227, 7.306073, 7.420966, 7.535905, 7.650891, 7.765922, 7.880998, 
    7.996119, 8.111284, 8.226493, 8.341744, 8.45704, 8.572376, 8.687756, 
    8.803176, 8.918637, 9.034139, 9.14968, 9.265261, 9.38088, 9.496539, 
    9.612235, 9.727969, 9.84374, 9.959547, 10.07539, 10.19127, 10.30718, 
    10.42313, 10.53911, 10.65513, 10.77118, 10.88726, 11.00337, 11.11952, 
    11.23569, 11.3519, 11.46814, 11.5844, 11.7007, 11.81702, 11.93337, 
    12.04975, 12.16616, 12.28259, 12.39905, 12.51553, 12.63204, 12.74857, 
    12.86513, 12.98171, 13.09831, 13.21494, 13.33158, 13.44825, 13.56494, 
    13.68165, 13.79838, 13.91513, 14.03189, 14.14868, 14.26548, 14.3823, 
    14.49914, 14.61599, 14.73286, 14.84974, 14.96664, 15.08355, 15.20047, 
    15.31741, 15.43436, 15.55132, 15.66829, 15.78527, 15.90226, 16.01927, 
    16.13628, 16.2533, 16.37033, 16.48736, 16.6044, 16.72145, 16.83851, 
    16.95557, 17.07263, 17.1897, 17.30678, 17.42385, 17.54093, 17.65801, 
    17.77509, 17.89218, 18.00926, 18.12634, 18.24343, 18.36051, 18.47759, 
    18.59467, 18.71174, 18.82882, 18.94588, 19.06295, 19.18001, 19.29706, 
    19.41411, 19.53115, 19.64819, 19.76521, 19.88223, 19.99924, 20.11624, 
    20.23323, 20.35022, 20.46719, 20.58414, 20.70109, 20.81803, 20.93495, 
    21.05186, 21.16875, 21.28563, 21.4025, 21.51935, 21.63618, 21.75299, 
    21.86979, 21.98658, 22.10334, 22.22009, 22.33681, 22.45352, 22.5702, 
    22.68687, 22.80351, 22.92013, 23.03673, 23.15331, 23.26986, 23.38639, 
    23.5029, 23.61938, 23.73583, 23.85226, 23.96866, 24.08503, 24.20138, 
    24.3177, 24.43399, 24.55025, 24.66648, 24.78269, 24.89886, 25.015, 
    25.13111, 25.24718, 25.36323, 25.47924, 25.59521, 25.71115, 25.82706, 
    25.94294, 26.05877, 26.17458, 26.29034, 26.40607, 26.52176, 26.63741, 
    26.75303, 26.8686, 26.98413, 27.09963, 27.21508, 27.3305, 27.44587, 
    27.5612, 27.67649, 27.79173, 27.90694, 28.02209, 28.13721, 28.25228, 
    28.3673, 28.48228, 28.59721, 28.7121, 28.82693, 28.94173, 29.05647, 
    29.17116, 29.28581, 29.4004, 29.51495, 29.62945, 29.74389, 29.85829, 
    29.97263, 30.08692, 30.20116, 30.31534, 30.42948, 30.54355, 30.65758, 
    30.77155, 30.88546, 30.99932, 31.11312, 31.22687, 31.34056, 31.45419, 
    31.56777, 31.68129, 31.79474, 31.90814, 32.02148, 32.13477, 32.24799, 
    32.36115, 32.47424, 32.58728, 32.70026, 32.81317, 32.92603, 33.03881, 
    33.15154, 33.2642, 33.3768, 33.48933, 33.6018, 33.7142, 33.82654, 
    33.93881, 34.05101, 34.16315, 34.27523, 34.38723, 34.49916, 34.61103, 
    34.72283, 34.83456, 34.94622, 35.05782, 35.16933, 35.28079, 35.39217, 
    35.50348, 35.61472, 35.72588, 35.83698, 35.94799, 36.05894, 36.16982, 
    36.28062, 36.39135, 36.502, 36.61258, 36.72309, 36.83352, 36.94387, 
    37.05415, 37.16436, 37.27448, 37.38453, 37.4945, 37.6044,
  -11.48458, -11.38275, -11.28084, -11.17882, -11.07671, -10.9745, -10.8722, 
    -10.7698, -10.6673, -10.56471, -10.46202, -10.35924, -10.25636, 
    -10.15338, -10.05031, -9.947146, -9.843886, -9.740532, -9.637082, 
    -9.533537, -9.429898, -9.326165, -9.222338, -9.118417, -9.014401, 
    -8.910293, -8.80609, -8.701794, -8.597404, -8.492923, -8.388347, 
    -8.283679, -8.178919, -8.074065, -7.96912, -7.864082, -7.758953, 
    -7.653732, -7.548419, -7.443015, -7.33752, -7.231934, -7.126256, 
    -7.020489, -6.91463, -6.808682, -6.702644, -6.596516, -6.490297, 
    -6.38399, -6.277594, -6.171108, -6.064533, -5.95787, -5.851119, 
    -5.744279, -5.637352, -5.530336, -5.423234, -5.316044, -5.208766, 
    -5.101403, -4.993952, -4.886415, -4.778792, -4.671083, -4.563289, 
    -4.455409, -4.347445, -4.239395, -4.13126, -4.023041, -3.914738, 
    -3.806351, -3.697881, -3.589327, -3.48069, -3.37197, -3.263168, 
    -3.154283, -3.045317, -2.936269, -2.827139, -2.717928, -2.608636, 
    -2.499264, -2.389811, -2.280278, -2.170666, -2.060974, -1.951203, 
    -1.841353, -1.731425, -1.621418, -1.511334, -1.401171, -1.290932, 
    -1.180615, -1.070222, -0.9597527, -0.849207, -0.7385857, -0.6278889, 
    -0.517117, -0.4062704, -0.2953493, -0.1843541, -0.07328518, 0.03785719, 
    0.1490726, 0.2603609, 0.3717215, 0.4831541, 0.5946586, 0.7062343, 
    0.8178811, 0.9295986, 1.041386, 1.153244, 1.265171, 1.377168, 1.489233, 
    1.601367, 1.713569, 1.825839, 1.938176, 2.050581, 2.163051, 2.275589, 
    2.388191, 2.50086, 2.613594, 2.726392, 2.839255, 2.952181, 3.065171, 
    3.178225, 3.291341, 3.40452, 3.51776, 3.631062, 3.744425, 3.857849, 
    3.971334, 4.084877, 4.198482, 4.312144, 4.425866, 4.539646, 4.653483, 
    4.767378, 4.88133, 4.995339, 5.109404, 5.223525, 5.3377, 5.451931, 
    5.566216, 5.680555, 5.794948, 5.909394, 6.023892, 6.138443, 6.253046, 
    6.3677, 6.482404, 6.597159, 6.711965, 6.826819, 6.941723, 7.056675, 
    7.171676, 7.286724, 7.401819, 7.516962, 7.63215, 7.747385, 7.862664, 
    7.977989, 8.093358, 8.208772, 8.324228, 8.439728, 8.555269, 8.670854, 
    8.78648, 8.902146, 9.017854, 9.133601, 9.249389, 9.365215, 9.48108, 
    9.596983, 9.712924, 9.828902, 9.944917, 10.06097, 10.17706, 10.29318, 
    10.40933, 10.52552, 10.64175, 10.75801, 10.8743, 10.99062, 11.10697, 
    11.22336, 11.33978, 11.45622, 11.5727, 11.6892, 11.80574, 11.9223, 
    12.03889, 12.15551, 12.27215, 12.38882, 12.50551, 12.62223, 12.73898, 
    12.85575, 12.97254, 13.08935, 13.20619, 13.32305, 13.43993, 13.55683, 
    13.67375, 13.7907, 13.90766, 14.02464, 14.14163, 14.25865, 14.37568, 
    14.49273, 14.60979, 14.72688, 14.84397, 14.96108, 15.07821, 15.19534, 
    15.31249, 15.42966, 15.54683, 15.66402, 15.78121, 15.89842, 16.01564, 
    16.13286, 16.2501, 16.36734, 16.48459, 16.60185, 16.71911, 16.83638, 
    16.95366, 17.07093, 17.18822, 17.3055, 17.4228, 17.54009, 17.65738, 
    17.77468, 17.89198, 18.00928, 18.12658, 18.24387, 18.36117, 18.47847, 
    18.59576, 18.71305, 18.83034, 18.94762, 19.0649, 19.18217, 19.29944, 
    19.4167, 19.53396, 19.65121, 19.76845, 19.88568, 20.0029, 20.12012, 
    20.23733, 20.35452, 20.4717, 20.58888, 20.70604, 20.82319, 20.94032, 
    21.05744, 21.17455, 21.29165, 21.40872, 21.52579, 21.64283, 21.75986, 
    21.87687, 21.99387, 22.11085, 22.2278, 22.34474, 22.46166, 22.57856, 
    22.69544, 22.81229, 22.92913, 23.04594, 23.16273, 23.27949, 23.39623, 
    23.51295, 23.62964, 23.7463, 23.86294, 23.97956, 24.09614, 24.2127, 
    24.32923, 24.44573, 24.5622, 24.67864, 24.79505, 24.91143, 25.02778, 
    25.1441, 25.26039, 25.37664, 25.49286, 25.60904, 25.72519, 25.84131, 
    25.95739, 26.07344, 26.18945, 26.30542, 26.42135, 26.53725, 26.65311, 
    26.76893, 26.88471, 27.00045, 27.11615, 27.23181, 27.34743, 27.46301, 
    27.57855, 27.69404, 27.80949, 27.92489, 28.04026, 28.15557, 28.27085, 
    28.38607, 28.50126, 28.61639, 28.73148, 28.84652, 28.96151, 29.07646, 
    29.19135, 29.3062, 29.421, 29.53574, 29.65044, 29.76509, 29.87968, 
    29.99422, 30.10871, 30.22315, 30.33754, 30.45187, 30.56614, 30.68036, 
    30.79453, 30.90864, 31.0227, 31.1367, 31.25064, 31.36453, 31.47836, 
    31.59213, 31.70584, 31.81949, 31.93309, 32.04662, 32.1601, 32.27351, 
    32.38686, 32.50016, 32.61339, 32.72655, 32.83966, 32.95271, 33.06569, 
    33.1786, 33.29145, 33.40424, 33.51697, 33.62962, 33.74222, 33.85474, 
    33.96721, 34.0796, 34.19193, 34.30418, 34.41637, 34.5285, 34.64055, 
    34.75254, 34.86446, 34.9763, 35.08808, 35.19978, 35.31142, 35.42299, 
    35.53448, 35.6459, 35.75725, 35.86853, 35.97973, 36.09086, 36.20192, 
    36.3129, 36.42381, 36.53465, 36.6454, 36.75609, 36.8667, 36.97723, 
    37.08769, 37.19807, 37.30838, 37.4186, 37.52875, 37.63882,
  -11.53374, -11.43177, -11.32972, -11.22756, -11.12531, -11.02296, 
    -10.92052, -10.81797, -10.71534, -10.6126, -10.50977, -10.40684, 
    -10.30382, -10.2007, -10.09749, -9.994179, -9.890773, -9.787272, 
    -9.683677, -9.579986, -9.4762, -9.37232, -9.268345, -9.164275, -9.060112, 
    -8.955853, -8.851501, -8.747056, -8.642516, -8.537884, -8.433157, 
    -8.328338, -8.223425, -8.11842, -8.013322, -7.908131, -7.802848, 
    -7.697473, -7.592006, -7.486447, -7.380797, -7.275055, -7.169222, 
    -7.063298, -6.957283, -6.851177, -6.744981, -6.638694, -6.532318, 
    -6.425851, -6.319295, -6.21265, -6.105915, -5.999092, -5.892179, 
    -5.785178, -5.678089, -5.570911, -5.463645, -5.356292, -5.248852, 
    -5.141324, -5.033709, -4.926008, -4.81822, -4.710345, -4.602385, 
    -4.494339, -4.386207, -4.277989, -4.169687, -4.061301, -3.952829, 
    -3.844274, -3.735634, -3.62691, -3.518103, -3.409213, -3.30024, 
    -3.191184, -3.082046, -2.972826, -2.863524, -2.75414, -2.644675, 
    -2.535129, -2.425502, -2.315795, -2.206008, -2.096141, -1.986194, 
    -1.876168, -1.766064, -1.65588, -1.545619, -1.435279, -1.324862, 
    -1.214367, -1.103795, -0.9931462, -0.8824212, -0.77162, -0.6607431, 
    -0.5497906, -0.4387631, -0.3276607, -0.2164838, -0.1052328, 0.006091967, 
    0.1174902, 0.2289616, 0.3405057, 0.4521223, 0.563811, 0.6755714, 
    0.7874032, 0.8993059, 1.011279, 1.123323, 1.235437, 1.34762, 1.459873, 
    1.572194, 1.684584, 1.797042, 1.909568, 2.022161, 2.134821, 2.247548, 
    2.36034, 2.473199, 2.586123, 2.699113, 2.812166, 2.925285, 3.038467, 
    3.151712, 3.265021, 3.378392, 3.491826, 3.605322, 3.718879, 3.832497, 
    3.946176, 4.059915, 4.173713, 4.287572, 4.401489, 4.515465, 4.629499, 
    4.74359, 4.857739, 4.971945, 5.086208, 5.200526, 5.3149, 5.429329, 
    5.543813, 5.658351, 5.772943, 5.887589, 6.002287, 6.117038, 6.231841, 
    6.346695, 6.461601, 6.576557, 6.691564, 6.80662, 6.921726, 7.03688, 
    7.152084, 7.267334, 7.382633, 7.497979, 7.613371, 7.728809, 7.844293, 
    7.959822, 8.075396, 8.191013, 8.306675, 8.422379, 8.538127, 8.653917, 
    8.769749, 8.885621, 9.001535, 9.11749, 9.233483, 9.349517, 9.465589, 
    9.581699, 9.697848, 9.814034, 9.930257, 10.04652, 10.16281, 10.27914, 
    10.39551, 10.51191, 10.62834, 10.74481, 10.86131, 10.97784, 11.0944, 
    11.211, 11.32763, 11.44428, 11.56097, 11.67769, 11.79443, 11.9112, 
    12.028, 12.14483, 12.26169, 12.37857, 12.49547, 12.61241, 12.72936, 
    12.84634, 12.96335, 13.08037, 13.19742, 13.3145, 13.43159, 13.5487, 
    13.66584, 13.78299, 13.90017, 14.01736, 14.13457, 14.2518, 14.36905, 
    14.48631, 14.60359, 14.72088, 14.83819, 14.95552, 15.07285, 15.19021, 
    15.30757, 15.42495, 15.54234, 15.65974, 15.77715, 15.89457, 16.012, 
    16.12944, 16.24689, 16.36435, 16.48181, 16.59929, 16.71676, 16.83425, 
    16.95174, 17.06923, 17.18673, 17.30423, 17.42174, 17.53925, 17.65676, 
    17.77427, 17.89178, 18.00929, 18.12681, 18.24432, 18.36183, 18.47934, 
    18.59685, 18.71436, 18.83186, 18.94936, 19.06685, 19.18434, 19.30182, 
    19.4193, 19.53677, 19.65423, 19.77169, 19.88914, 20.00657, 20.124, 
    20.24142, 20.35883, 20.47623, 20.59362, 20.71099, 20.82836, 20.94571, 
    21.06304, 21.18037, 21.29767, 21.41496, 21.53224, 21.6495, 21.76674, 
    21.88397, 22.00118, 22.11837, 22.23554, 22.35269, 22.46982, 22.58694, 
    22.70402, 22.82109, 22.93814, 23.05516, 23.17216, 23.28914, 23.40609, 
    23.52302, 23.63992, 23.7568, 23.87365, 23.99047, 24.10727, 24.22404, 
    24.34078, 24.45749, 24.57417, 24.69082, 24.80745, 24.92404, 25.0406, 
    25.15712, 25.27362, 25.39008, 25.50651, 25.6229, 25.73926, 25.85559, 
    25.97188, 26.08813, 26.20435, 26.32053, 26.43667, 26.55277, 26.66884, 
    26.78487, 26.90086, 27.0168, 27.13271, 27.24858, 27.3644, 27.48018, 
    27.59593, 27.71162, 27.82728, 27.94289, 28.05846, 28.17398, 28.28946, 
    28.40489, 28.52027, 28.63561, 28.7509, 28.86614, 28.98134, 29.09649, 
    29.21158, 29.32663, 29.44163, 29.55658, 29.67148, 29.78632, 29.90112, 
    30.01586, 30.13055, 30.24519, 30.35977, 30.4743, 30.58878, 30.7032, 
    30.81756, 30.93187, 31.04612, 31.16032, 31.27446, 31.38854, 31.50257, 
    31.61654, 31.73044, 31.84429, 31.95808, 32.07181, 32.18548, 32.29909, 
    32.41264, 32.52612, 32.63955, 32.75291, 32.86621, 32.97944, 33.09261, 
    33.20572, 33.31876, 33.43174, 33.54466, 33.65751, 33.77029, 33.883, 
    33.99566, 34.10824, 34.22075, 34.3332, 34.44558, 34.55789, 34.67013, 
    34.7823, 34.89441, 35.00644, 35.1184, 35.23029, 35.34211, 35.45386, 
    35.56554, 35.67714, 35.78868, 35.90014, 36.01152, 36.12284, 36.23407, 
    36.34524, 36.45633, 36.56735, 36.67829, 36.78915, 36.89994, 37.01065, 
    37.12129, 37.23185, 37.34233, 37.45274, 37.56306, 37.67331,
  -11.58297, -11.48087, -11.37867, -11.27638, -11.17399, -11.0715, -10.96891, 
    -10.86623, -10.76345, -10.66057, -10.5576, -10.45453, -10.35136, 
    -10.2481, -10.14474, -10.04128, -9.937735, -9.834088, -9.730346, 
    -9.626509, -9.522576, -9.418549, -9.314425, -9.210208, -9.105896, 
    -9.001489, -8.896988, -8.792392, -8.687702, -8.582919, -8.478042, 
    -8.37307, -8.268005, -8.162848, -8.057597, -7.952253, -7.846817, 
    -7.741288, -7.635666, -7.529953, -7.424147, -7.318249, -7.21226, 
    -7.106179, -7.000007, -6.893744, -6.78739, -6.680945, -6.57441, 
    -6.467784, -6.361069, -6.254263, -6.147368, -6.040384, -5.933311, 
    -5.826148, -5.718896, -5.611557, -5.504128, -5.396612, -5.289008, 
    -5.181315, -5.073536, -4.96567, -4.857717, -4.749676, -4.64155, 
    -4.533337, -4.425038, -4.316654, -4.208184, -4.099629, -3.990989, 
    -3.882264, -3.773455, -3.664562, -3.555585, -3.446524, -3.33738, 
    -3.228153, -3.118842, -3.00945, -2.899975, -2.790418, -2.68078, -2.57106, 
    -2.461259, -2.351378, -2.241416, -2.131373, -2.02125, -1.911049, 
    -1.800767, -1.690407, -1.579968, -1.46945, -1.358855, -1.248182, 
    -1.137431, -1.026603, -0.9156982, -0.8047169, -0.6936595, -0.5825263, 
    -0.4713176, -0.3600336, -0.2486748, -0.1372415, -0.02573407, 0.08584723, 
    0.197502, 0.30923, 0.4210307, 0.5329039, 0.6448492, 0.7568662, 0.8689546, 
    0.9811141, 1.093344, 1.205645, 1.318015, 1.430455, 1.542964, 1.655542, 
    1.768188, 1.880903, 1.993685, 2.106535, 2.219451, 2.332434, 2.445484, 
    2.558599, 2.671779, 2.785025, 2.898335, 3.011709, 3.125147, 3.238649, 
    3.352213, 3.465841, 3.57953, 3.693281, 3.807094, 3.920967, 4.034901, 
    4.148896, 4.262949, 4.377063, 4.491235, 4.605466, 4.719755, 4.834101, 
    4.948504, 5.062964, 5.177481, 5.292054, 5.406682, 5.521364, 5.636102, 
    5.750894, 5.865739, 5.980638, 6.095589, 6.210592, 6.325648, 6.440755, 
    6.555912, 6.671121, 6.78638, 6.901688, 7.017045, 7.132451, 7.247905, 
    7.363407, 7.478956, 7.594552, 7.710195, 7.825883, 7.941617, 8.057395, 
    8.173218, 8.289084, 8.404995, 8.520948, 8.636945, 8.752982, 8.869061, 
    8.985183, 9.101343, 9.217545, 9.333785, 9.450066, 9.566383, 9.68274, 
    9.799134, 9.915565, 10.03203, 10.14854, 10.26508, 10.38165, 10.49826, 
    10.6149, 10.73158, 10.84829, 10.96503, 11.08181, 11.19861, 11.31545, 
    11.43232, 11.54922, 11.66614, 11.7831, 11.90008, 12.0171, 12.13414, 
    12.2512, 12.36829, 12.48541, 12.60256, 12.71973, 12.83692, 12.95414, 
    13.07138, 13.18864, 13.30592, 13.42323, 13.54056, 13.65791, 13.77527, 
    13.89266, 14.01007, 14.12749, 14.24494, 14.3624, 14.47987, 14.59737, 
    14.71488, 14.8324, 14.94994, 15.06749, 15.18506, 15.30264, 15.42023, 
    15.53783, 15.65545, 15.77307, 15.89071, 16.00836, 16.12601, 16.24368, 
    16.36135, 16.47903, 16.59672, 16.71441, 16.83211, 16.94981, 17.06752, 
    17.18524, 17.30296, 17.42068, 17.5384, 17.65613, 17.77385, 17.89158, 
    18.00931, 18.12704, 18.24477, 18.3625, 18.48022, 18.59794, 18.71567, 
    18.83338, 18.9511, 19.06881, 19.18651, 19.30421, 19.4219, 19.53959, 
    19.65726, 19.77494, 19.8926, 20.01025, 20.1279, 20.24553, 20.36316, 
    20.48077, 20.59837, 20.71596, 20.83354, 20.95111, 21.06866, 21.18619, 
    21.30371, 21.42122, 21.53871, 21.65619, 21.77364, 21.89108, 22.0085, 
    22.12591, 22.24329, 22.36066, 22.478, 22.59533, 22.71263, 22.82991, 
    22.94717, 23.06441, 23.18162, 23.29881, 23.41597, 23.53311, 23.65023, 
    23.76732, 23.88438, 24.00142, 24.11842, 24.2354, 24.35236, 24.46928, 
    24.58617, 24.70303, 24.81987, 24.93667, 25.05344, 25.17017, 25.28688, 
    25.40355, 25.52019, 25.63679, 25.75336, 25.86989, 25.98639, 26.10285, 
    26.21928, 26.33567, 26.45202, 26.56833, 26.6846, 26.80084, 26.91703, 
    27.03319, 27.1493, 27.26538, 27.38141, 27.4974, 27.61334, 27.72925, 
    27.84511, 27.96092, 28.07669, 28.19242, 28.3081, 28.42374, 28.53933, 
    28.65487, 28.77036, 28.88581, 29.00121, 29.11656, 29.23186, 29.34711, 
    29.46231, 29.57746, 29.69256, 29.8076, 29.9226, 30.03754, 30.15243, 
    30.26727, 30.38205, 30.49678, 30.61145, 30.72607, 30.84064, 30.95514, 
    31.0696, 31.18399, 31.29833, 31.41261, 31.52683, 31.64099, 31.7551, 
    31.86914, 31.98313, 32.09705, 32.21091, 32.32472, 32.43846, 32.55214, 
    32.66576, 32.77931, 32.8928, 33.00623, 33.11959, 33.23289, 33.34613, 
    33.4593, 33.5724, 33.68544, 33.79842, 33.91132, 34.02416, 34.13693, 
    34.24963, 34.36227, 34.47484, 34.58734, 34.69976, 34.81213, 34.92441, 
    35.03663, 35.14878, 35.26086, 35.37286, 35.4848, 35.59666, 35.70845, 
    35.82016, 35.93181, 36.04338, 36.15487, 36.2663, 36.37764, 36.48891, 
    36.60011, 36.71123, 36.82228, 36.93325, 37.04414, 37.15496, 37.26569, 
    37.37635, 37.48694, 37.59744, 37.70787,
  -11.63228, -11.53004, -11.4277, -11.32527, -11.22274, -11.12011, -11.01738, 
    -10.91456, -10.81163, -10.70861, -10.6055, -10.50229, -10.39898, 
    -10.29557, -10.19207, -10.08847, -9.984771, -9.880979, -9.777091, 
    -9.673107, -9.569027, -9.464852, -9.360581, -9.256216, -9.151754, 
    -9.047199, -8.942548, -8.837803, -8.732963, -8.628028, -8.523, -8.417877, 
    -8.31266, -8.20735, -8.101946, -7.996449, -7.890859, -7.785176, 
    -7.679399, -7.573531, -7.46757, -7.361516, -7.255371, -7.149133, 
    -7.042804, -6.936383, -6.829872, -6.723269, -6.616574, -6.50979, 
    -6.402915, -6.295949, -6.188894, -6.081748, -5.974514, -5.867189, 
    -5.759776, -5.652273, -5.544682, -5.437002, -5.329234, -5.221378, 
    -5.113434, -5.005403, -4.897284, -4.789077, -4.680785, -4.572405, 
    -4.463939, -4.355387, -4.246749, -4.138026, -4.029217, -3.920324, 
    -3.811345, -3.702282, -3.593134, -3.483902, -3.374587, -3.265188, 
    -3.155706, -3.046141, -2.936494, -2.826764, -2.716952, -2.607058, 
    -2.497083, -2.387026, -2.276889, -2.166671, -2.056372, -1.945994, 
    -1.835536, -1.724998, -1.614382, -1.503686, -1.392912, -1.28206, 
    -1.17113, -1.060123, -0.9490383, -0.8378768, -0.7266387, -0.6153245, 
    -0.5039343, -0.3924686, -0.2809276, -0.1693117, -0.05762133, 0.05414328, 
    0.1659818, 0.2778938, 0.3898789, 0.5019369, 0.6140673, 0.7262699, 
    0.8385442, 0.9508899, 1.063307, 1.175794, 1.288352, 1.400979, 1.513677, 
    1.626443, 1.739278, 1.852182, 1.965153, 2.078193, 2.191299, 2.304473, 
    2.417713, 2.531019, 2.644391, 2.757829, 2.871331, 2.984898, 3.098529, 
    3.212224, 3.325982, 3.439803, 3.553686, 3.667632, 3.781639, 3.895708, 
    4.009838, 4.124028, 4.238278, 4.352587, 4.466956, 4.581384, 4.69587, 
    4.810414, 4.925015, 5.039674, 5.154389, 5.26916, 5.383987, 5.498869, 
    5.613807, 5.728798, 5.843844, 5.958943, 6.074095, 6.1893, 6.304557, 
    6.419866, 6.535225, 6.650636, 6.766097, 6.881608, 6.997168, 7.112778, 
    7.228435, 7.344141, 7.459894, 7.575695, 7.691541, 7.807435, 7.923373, 
    8.039357, 8.155385, 8.271458, 8.387574, 8.503734, 8.619936, 8.736181, 
    8.852468, 8.968795, 9.085163, 9.201572, 9.318021, 9.434508, 9.551035, 
    9.667601, 9.784203, 9.900843, 10.01752, 10.13423, 10.25098, 10.36777, 
    10.48458, 10.60144, 10.71833, 10.83525, 10.9522, 11.06918, 11.1862, 
    11.30325, 11.42033, 11.53744, 11.65458, 11.77174, 11.88894, 12.00616, 
    12.12342, 12.24069, 12.358, 12.47533, 12.59269, 12.71007, 12.82748, 
    12.94491, 13.06236, 13.17984, 13.29733, 13.41485, 13.5324, 13.64996, 
    13.76754, 13.88514, 14.00276, 14.1204, 14.23806, 14.35573, 14.47342, 
    14.59113, 14.70886, 14.8266, 14.94435, 15.06212, 15.1799, 15.29769, 
    15.4155, 15.53332, 15.65115, 15.76899, 15.88684, 16.00471, 16.12258, 
    16.24046, 16.35834, 16.47624, 16.59414, 16.71205, 16.82997, 16.94789, 
    17.06581, 17.18374, 17.30168, 17.41961, 17.53755, 17.65549, 17.77344, 
    17.89138, 18.00933, 18.12727, 18.24522, 18.36316, 18.4811, 18.59904, 
    18.71698, 18.83491, 18.95284, 19.07077, 19.18869, 19.3066, 19.42451, 
    19.54241, 19.66031, 19.77819, 19.89607, 20.01394, 20.1318, 20.24965, 
    20.36749, 20.48532, 20.60314, 20.72094, 20.83873, 20.95651, 21.07428, 
    21.19203, 21.30977, 21.42749, 21.54519, 21.66288, 21.78055, 21.89821, 
    22.01584, 22.13346, 22.25106, 22.36864, 22.4862, 22.60374, 22.72125, 
    22.83875, 22.95622, 23.07367, 23.1911, 23.3085, 23.42588, 23.54323, 
    23.66056, 23.77786, 23.89513, 24.01238, 24.1296, 24.24679, 24.36396, 
    24.48109, 24.59819, 24.71527, 24.83231, 24.94932, 25.0663, 25.18325, 
    25.30017, 25.41705, 25.5339, 25.65071, 25.76749, 25.88423, 26.00094, 
    26.11761, 26.23425, 26.35084, 26.4674, 26.58392, 26.7004, 26.81684, 
    26.93325, 27.04961, 27.16593, 27.28221, 27.39845, 27.51464, 27.6308, 
    27.74691, 27.86297, 27.97899, 28.09497, 28.2109, 28.32679, 28.44263, 
    28.55842, 28.67417, 28.78986, 28.90551, 29.02111, 29.13667, 29.25217, 
    29.36762, 29.48303, 29.59838, 29.71368, 29.82893, 29.94412, 30.05927, 
    30.17436, 30.28939, 30.40438, 30.51931, 30.63418, 30.749, 30.86376, 
    30.97847, 31.09312, 31.20771, 31.32224, 31.43672, 31.55114, 31.6655, 
    31.7798, 31.89404, 32.00822, 32.12234, 32.2364, 32.3504, 32.46433, 
    32.57821, 32.69202, 32.80577, 32.91945, 33.03307, 33.14663, 33.26012, 
    33.37355, 33.48691, 33.6002, 33.71343, 33.8266, 33.93969, 34.05272, 
    34.16568, 34.27858, 34.3914, 34.50415, 34.61684, 34.72946, 34.842, 
    34.95448, 35.06689, 35.17922, 35.29148, 35.40368, 35.51579, 35.62784, 
    35.73981, 35.85172, 35.96354, 36.07529, 36.18697, 36.29858, 36.41011, 
    36.52156, 36.63294, 36.74424, 36.85546, 36.96661, 37.07769, 37.18868, 
    37.2996, 37.41044, 37.5212, 37.63189, 37.74249,
  -11.68167, -11.57929, -11.47681, -11.37424, -11.27157, -11.16879, 
    -11.06593, -10.96296, -10.8599, -10.75673, -10.65348, -10.55012, 
    -10.44667, -10.34311, -10.23947, -10.13572, -10.03188, -9.927944, 
    -9.823911, -9.71978, -9.615554, -9.511231, -9.406813, -9.302299, 
    -9.197689, -9.092983, -8.988183, -8.883287, -8.778297, -8.673212, 
    -8.568032, -8.462758, -8.357389, -8.251926, -8.14637, -8.040719, 
    -7.934975, -7.829138, -7.723207, -7.617183, -7.511066, -7.404857, 
    -7.298555, -7.192161, -7.085675, -6.979096, -6.872427, -6.765665, 
    -6.658812, -6.551868, -6.444833, -6.337708, -6.230492, -6.123185, 
    -6.015789, -5.908303, -5.800727, -5.693062, -5.585307, -5.477464, 
    -5.369532, -5.261511, -5.153403, -5.045206, -4.936922, -4.828549, 
    -4.72009, -4.611544, -4.502911, -4.394191, -4.285385, -4.176493, 
    -4.067515, -3.958452, -3.849304, -3.74007, -3.630752, -3.52135, 
    -3.411863, -3.302292, -3.192638, -3.082901, -2.97308, -2.863177, 
    -2.753191, -2.643123, -2.532973, -2.422741, -2.312428, -2.202034, 
    -2.09156, -1.981005, -1.87037, -1.759655, -1.64886, -1.537987, -1.427034, 
    -1.316003, -1.204894, -1.093707, -0.9824421, -0.8711001, -0.7596811, 
    -0.6481855, -0.5366136, -0.4249659, -0.3132425, -0.2014438, -0.08957019, 
    0.02237799, 0.1344004, 0.2464967, 0.3586666, 0.4709096, 0.5832255, 
    0.6956139, 0.8080743, 0.9206066, 1.03321, 1.145885, 1.25863, 1.371446, 
    1.484331, 1.597286, 1.710311, 1.823404, 1.936565, 2.049794, 2.163092, 
    2.276456, 2.389887, 2.503385, 2.616949, 2.730578, 2.844273, 2.958033, 
    3.071857, 3.185745, 3.299697, 3.413712, 3.52779, 3.641931, 3.756133, 
    3.870398, 3.984723, 4.099109, 4.213555, 4.328062, 4.442628, 4.557253, 
    4.671937, 4.786679, 4.901478, 5.016335, 5.131249, 5.24622, 5.361247, 
    5.476328, 5.591466, 5.706658, 5.821904, 5.937204, 6.052557, 6.167964, 
    6.283422, 6.398933, 6.514495, 6.630108, 6.745772, 6.861486, 6.97725, 
    7.093063, 7.208924, 7.324834, 7.440792, 7.556797, 7.672849, 7.788947, 
    7.905091, 8.02128, 8.137515, 8.253794, 8.370117, 8.486483, 8.602892, 
    8.719344, 8.835837, 8.952373, 9.068949, 9.185566, 9.302222, 9.418919, 
    9.535654, 9.652428, 9.769239, 9.886089, 10.00298, 10.1199, 10.23686, 
    10.35385, 10.47088, 10.58794, 10.70504, 10.82217, 10.93934, 11.05653, 
    11.17376, 11.29102, 11.40831, 11.52563, 11.64298, 11.76036, 11.87777, 
    11.99521, 12.11267, 12.23016, 12.34768, 12.46523, 12.5828, 12.70039, 
    12.81801, 12.93566, 13.05332, 13.17101, 13.28872, 13.40646, 13.52421, 
    13.64199, 13.75979, 13.8776, 13.99544, 14.11329, 14.23116, 14.34906, 
    14.46696, 14.58488, 14.70282, 14.82078, 14.93875, 15.05673, 15.17473, 
    15.29274, 15.41076, 15.5288, 15.64684, 15.7649, 15.88297, 16.00105, 
    16.11913, 16.23723, 16.35533, 16.47344, 16.59156, 16.70969, 16.82782, 
    16.94596, 17.0641, 17.18225, 17.3004, 17.41855, 17.53671, 17.65486, 
    17.77302, 17.89118, 18.00935, 18.12751, 18.24567, 18.36383, 18.48199, 
    18.60014, 18.71829, 18.83644, 18.95459, 19.07273, 19.19087, 19.309, 
    19.42712, 19.54524, 19.66335, 19.78145, 19.89955, 20.01763, 20.13571, 
    20.25378, 20.37183, 20.48988, 20.60791, 20.72593, 20.84394, 20.96193, 
    21.07992, 21.19788, 21.31583, 21.43377, 21.55169, 21.66959, 21.78748, 
    21.90535, 22.0232, 22.14104, 22.25885, 22.37664, 22.49441, 22.61217, 
    22.7299, 22.8476, 22.96529, 23.08295, 23.2006, 23.31821, 23.4358, 
    23.55337, 23.67091, 23.78842, 23.90591, 24.02337, 24.1408, 24.25821, 
    24.37558, 24.49293, 24.61024, 24.72753, 24.84478, 24.96201, 25.0792, 
    25.19636, 25.31348, 25.43058, 25.54763, 25.66466, 25.78165, 25.8986, 
    26.01552, 26.1324, 26.24924, 26.36605, 26.48281, 26.59954, 26.71623, 
    26.83288, 26.94949, 27.06606, 27.18259, 27.29908, 27.41553, 27.53193, 
    27.64829, 27.7646, 27.88087, 27.9971, 28.11328, 28.22942, 28.34551, 
    28.46156, 28.57755, 28.6935, 28.80941, 28.92526, 29.04107, 29.15682, 
    29.27253, 29.38818, 29.50379, 29.61934, 29.73484, 29.8503, 29.96569, 
    30.08104, 30.19633, 30.31157, 30.42675, 30.54188, 30.65695, 30.77197, 
    30.88693, 31.00184, 31.11669, 31.23148, 31.34621, 31.46088, 31.5755, 
    31.69006, 31.80455, 31.91899, 32.03337, 32.14768, 32.26194, 32.37613, 
    32.49026, 32.60433, 32.71833, 32.83228, 32.94615, 33.05997, 33.17372, 
    33.2874, 33.40102, 33.51457, 33.62806, 33.74148, 33.85484, 33.96812, 
    34.08134, 34.19449, 34.30757, 34.42059, 34.53353, 34.6464, 34.75921, 
    34.87194, 34.98461, 35.0972, 35.20972, 35.32217, 35.43455, 35.54685, 
    35.65908, 35.77124, 35.88332, 35.99533, 36.10727, 36.21914, 36.33092, 
    36.44263, 36.55427, 36.66583, 36.77731, 36.88872, 37.00005, 37.1113, 
    37.22247, 37.33357, 37.44459, 37.55553, 37.66639, 37.77717,
  -11.73113, -11.62861, -11.526, -11.42328, -11.32047, -11.21756, -11.11455, 
    -11.01144, -10.90823, -10.80493, -10.70153, -10.59803, -10.49443, 
    -10.39074, -10.28695, -10.18306, -10.07907, -9.974987, -9.870807, 
    -9.766529, -9.662156, -9.557686, -9.453119, -9.348457, -9.243698, 
    -9.138844, -9.033895, -8.928848, -8.823708, -8.718472, -8.61314, 
    -8.507714, -8.402193, -8.296578, -8.190868, -8.085064, -7.979167, 
    -7.873175, -7.767089, -7.66091, -7.554637, -7.448272, -7.341814, 
    -7.235263, -7.128619, -7.021883, -6.915055, -6.808135, -6.701123, 
    -6.594019, -6.486825, -6.379539, -6.272162, -6.164695, -6.057137, 
    -5.949489, -5.84175, -5.733922, -5.626005, -5.517998, -5.409902, 
    -5.301716, -5.193443, -5.085081, -4.97663, -4.868092, -4.759466, 
    -4.650753, -4.541953, -4.433065, -4.32409, -4.21503, -4.105883, -3.99665, 
    -3.887332, -3.777928, -3.668439, -3.558866, -3.449208, -3.339465, 
    -3.229638, -3.119728, -3.009734, -2.899657, -2.789497, -2.679255, 
    -2.56893, -2.458523, -2.348035, -2.237465, -2.126814, -2.016082, 
    -1.90527, -1.794377, -1.683405, -1.572353, -1.461221, -1.350011, 
    -1.238722, -1.127355, -1.01591, -0.9043871, -0.792787, -0.6811098, 
    -0.569356, -0.4575259, -0.3456199, -0.2336381, -0.1215811, -0.009449041, 
    0.1027576, 0.2150385, 0.3273933, 0.4398217, 0.5523232, 0.6648977, 
    0.7775446, 0.8902636, 1.003054, 1.115917, 1.22885, 1.341854, 1.454928, 
    1.568072, 1.681286, 1.794568, 1.90792, 2.02134, 2.134827, 2.248383, 
    2.362005, 2.475695, 2.589451, 2.703273, 2.817161, 2.931113, 3.045131, 
    3.159213, 3.273359, 3.387569, 3.501842, 3.616178, 3.730576, 3.845036, 
    3.959557, 4.07414, 4.188783, 4.303486, 4.41825, 4.533072, 4.647954, 
    4.762895, 4.877893, 4.992949, 5.108062, 5.223232, 5.338459, 5.453741, 
    5.569078, 5.684471, 5.799918, 5.91542, 6.030974, 6.146583, 6.262244, 
    6.377957, 6.493721, 6.609538, 6.725405, 6.841322, 6.95729, 7.073307, 
    7.189373, 7.305487, 7.42165, 7.53786, 7.654117, 7.770421, 7.886771, 
    8.003166, 8.119607, 8.236093, 8.352622, 8.469195, 8.585812, 8.702472, 
    8.819173, 8.935916, 9.0527, 9.169525, 9.286391, 9.403296, 9.520241, 
    9.637223, 9.754245, 9.871304, 9.9884, 10.10553, 10.2227, 10.33991, 
    10.45715, 10.57442, 10.69173, 10.80907, 10.92645, 11.04386, 11.1613, 
    11.27877, 11.39627, 11.5138, 11.63137, 11.74896, 11.86658, 11.98423, 
    12.10191, 12.21961, 12.33734, 12.4551, 12.57289, 12.69069, 12.80853, 
    12.92638, 13.04427, 13.16217, 13.2801, 13.39805, 13.51602, 13.63401, 
    13.75202, 13.87005, 13.9881, 14.10617, 14.22426, 14.34236, 14.46048, 
    14.57862, 14.69678, 14.81495, 14.93313, 15.05133, 15.16955, 15.28777, 
    15.40601, 15.52426, 15.64252, 15.7608, 15.87908, 15.99738, 16.11568, 
    16.23399, 16.35231, 16.47064, 16.58898, 16.70732, 16.82567, 16.94402, 
    17.06238, 17.18074, 17.29911, 17.41748, 17.53585, 17.65423, 17.77261, 
    17.89098, 18.00936, 18.12774, 18.24612, 18.3645, 18.48287, 18.60124, 
    18.71961, 18.83798, 18.95634, 19.0747, 19.19305, 19.3114, 19.42974, 
    19.54808, 19.6664, 19.78472, 19.90303, 20.02134, 20.13963, 20.25791, 
    20.37618, 20.49444, 20.61269, 20.73093, 20.84916, 20.96737, 21.08556, 
    21.20375, 21.32191, 21.44007, 21.5582, 21.67632, 21.79442, 21.91251, 
    22.03057, 22.14862, 22.26665, 22.38466, 22.50265, 22.62061, 22.73856, 
    22.85648, 22.97438, 23.09226, 23.21011, 23.32794, 23.44575, 23.56353, 
    23.68128, 23.79901, 23.91671, 24.03438, 24.15203, 24.26965, 24.38723, 
    24.50479, 24.62232, 24.73982, 24.85728, 24.97472, 25.09212, 25.20949, 
    25.32683, 25.44413, 25.5614, 25.67864, 25.79584, 25.913, 26.03012, 
    26.14721, 26.26427, 26.38128, 26.49826, 26.6152, 26.7321, 26.84896, 
    26.96578, 27.08255, 27.19929, 27.31598, 27.43264, 27.54925, 27.66581, 
    27.78234, 27.89882, 28.01525, 28.13164, 28.24798, 28.36428, 28.48053, 
    28.59673, 28.71288, 28.82899, 28.94505, 29.06106, 29.17702, 29.29293, 
    29.40879, 29.52459, 29.64035, 29.75606, 29.87171, 29.98731, 30.10285, 
    30.21835, 30.33379, 30.44917, 30.5645, 30.67977, 30.79499, 30.91015, 
    31.02526, 31.1403, 31.25529, 31.37022, 31.48509, 31.59991, 31.71466, 
    31.82936, 31.94399, 32.05856, 32.17307, 32.28753, 32.40191, 32.51624, 
    32.6305, 32.7447, 32.85884, 32.97291, 33.08692, 33.20086, 33.31474, 
    33.42855, 33.54229, 33.65597, 33.76958, 33.88313, 33.9966, 34.11002, 
    34.22335, 34.33663, 34.44983, 34.56296, 34.67603, 34.78902, 34.90194, 
    35.01479, 35.12757, 35.24028, 35.35291, 35.46548, 35.57797, 35.69038, 
    35.80273, 35.915, 36.02719, 36.13931, 36.25136, 36.36333, 36.47522, 
    36.58704, 36.69878, 36.81044, 36.92204, 37.03354, 37.14498, 37.25633, 
    37.36761, 37.47881, 37.58992, 37.70097, 37.81192,
  -11.78067, -11.67801, -11.57526, -11.4724, -11.36945, -11.2664, -11.16325, 
    -11.06, -10.95665, -10.8532, -10.74966, -10.64602, -10.54228, -10.43844, 
    -10.3345, -10.23047, -10.12633, -10.02211, -9.917779, -9.813354, 
    -9.708835, -9.604217, -9.499502, -9.394691, -9.289784, -9.18478, 
    -9.07968, -8.974485, -8.869194, -8.763806, -8.658324, -8.552746, 
    -8.447073, -8.341305, -8.235442, -8.129484, -8.023433, -7.917286, 
    -7.811046, -7.704711, -7.598283, -7.491762, -7.385147, -7.278439, 
    -7.171638, -7.064744, -6.957757, -6.850678, -6.743508, -6.636245, 
    -6.52889, -6.421444, -6.313906, -6.206277, -6.098558, -5.990747, 
    -5.882847, -5.774856, -5.666775, -5.558604, -5.450344, -5.341994, 
    -5.233555, -5.125027, -5.016411, -4.907707, -4.798914, -4.690033, 
    -4.581065, -4.47201, -4.362867, -4.253637, -4.144321, -4.034919, 
    -3.925431, -3.815856, -3.706196, -3.596451, -3.486621, -3.376706, 
    -3.266707, -3.156624, -3.046457, -2.936206, -2.825872, -2.715455, 
    -2.604955, -2.494373, -2.383708, -2.272962, -2.162134, -2.051225, 
    -1.940236, -1.829165, -1.718015, -1.606784, -1.495474, -1.384084, 
    -1.272615, -1.161068, -1.049442, -0.9377382, -0.8259567, -0.7140978, 
    -0.6021618, -0.4901492, -0.3780601, -0.2658951, -0.1536543, -0.04133821, 
    0.07105289, 0.1835186, 0.2960587, 0.4086726, 0.5213602, 0.6341209, 
    0.7469546, 0.8598607, 0.9728389, 1.085889, 1.19901, 1.312203, 1.425466, 
    1.538799, 1.652202, 1.765675, 1.879217, 1.992828, 2.106507, 2.220253, 
    2.334068, 2.447949, 2.561898, 2.675913, 2.789993, 2.90414, 3.018351, 
    3.132627, 3.246968, 3.361372, 3.475841, 3.590372, 3.704966, 3.819622, 
    3.93434, 4.049119, 4.16396, 4.27886, 4.393821, 4.508842, 4.623922, 
    4.739061, 4.854259, 4.969514, 5.084827, 5.200197, 5.315623, 5.431106, 
    5.546645, 5.662238, 5.777887, 5.89359, 6.009347, 6.125157, 6.241021, 
    6.356936, 6.472904, 6.588924, 6.704995, 6.821116, 6.937288, 7.053509, 
    7.16978, 7.286099, 7.402467, 7.518883, 7.635345, 7.751855, 7.868412, 
    7.985013, 8.101661, 8.218353, 8.335091, 8.451871, 8.568695, 8.685562, 
    8.802472, 8.919424, 9.036417, 9.153451, 9.270525, 9.38764, 9.504793, 
    9.621986, 9.739218, 9.856486, 9.973793, 10.09114, 10.20852, 10.32593, 
    10.44338, 10.56087, 10.67839, 10.79594, 10.91353, 11.03115, 11.1488, 
    11.26649, 11.3842, 11.50195, 11.61972, 11.73753, 11.85536, 11.97323, 
    12.09112, 12.20904, 12.32698, 12.44495, 12.56295, 12.68097, 12.79902, 
    12.91709, 13.03519, 13.15331, 13.27145, 13.38962, 13.5078, 13.62601, 
    13.74423, 13.86248, 13.98075, 14.09903, 14.21733, 14.33566, 14.45399, 
    14.57235, 14.69072, 14.8091, 14.92751, 15.04592, 15.16435, 15.28279, 
    15.40125, 15.51972, 15.6382, 15.75669, 15.87519, 15.9937, 16.11222, 
    16.23075, 16.34929, 16.46783, 16.58639, 16.70495, 16.82351, 16.94208, 
    17.06066, 17.17924, 17.29782, 17.41641, 17.535, 17.65359, 17.77219, 
    17.89078, 18.00938, 18.12798, 18.24657, 18.36517, 18.48376, 18.60235, 
    18.72093, 18.83952, 18.9581, 19.07667, 19.19524, 19.31381, 19.43237, 
    19.55092, 19.66946, 19.788, 19.90653, 20.02505, 20.14356, 20.26206, 
    20.38054, 20.49902, 20.61749, 20.73594, 20.85438, 20.97281, 21.09122, 
    21.20962, 21.32801, 21.44637, 21.56473, 21.68306, 21.80138, 21.91968, 
    22.03796, 22.15623, 22.27447, 22.39269, 22.5109, 22.62908, 22.74724, 
    22.86538, 22.98349, 23.10158, 23.21965, 23.3377, 23.45572, 23.57371, 
    23.69168, 23.80962, 23.92753, 24.04542, 24.16328, 24.28111, 24.39891, 
    24.51668, 24.63442, 24.75213, 24.86981, 24.98746, 25.10507, 25.22265, 
    25.3402, 25.45772, 25.5752, 25.69264, 25.81005, 25.92743, 26.04477, 
    26.16207, 26.27933, 26.39655, 26.51374, 26.63089, 26.748, 26.86506, 
    26.98209, 27.09908, 27.21602, 27.33293, 27.44979, 27.5666, 27.68338, 
    27.80011, 27.91679, 28.03343, 28.15003, 28.26658, 28.38308, 28.49954, 
    28.61594, 28.7323, 28.84862, 28.96488, 29.08109, 29.19726, 29.31337, 
    29.42943, 29.54544, 29.6614, 29.77731, 29.89317, 30.00897, 30.12472, 
    30.24041, 30.35605, 30.47164, 30.58717, 30.70264, 30.81806, 30.93342, 
    31.04872, 31.16397, 31.27916, 31.39429, 31.50936, 31.62437, 31.73932, 
    31.85421, 31.96904, 32.08381, 32.19852, 32.31317, 32.42775, 32.54227, 
    32.65673, 32.77112, 32.88545, 32.99972, 33.11392, 33.22806, 33.34213, 
    33.45613, 33.57007, 33.68394, 33.79774, 33.91148, 34.02515, 34.13875, 
    34.25228, 34.36574, 34.47913, 34.59246, 34.70571, 34.81889, 34.932, 
    35.04504, 35.158, 35.2709, 35.38372, 35.49647, 35.60915, 35.72175, 
    35.83428, 35.94673, 36.05911, 36.17141, 36.28364, 36.3958, 36.50787, 
    36.61987, 36.7318, 36.84364, 36.95541, 37.0671, 37.17872, 37.29025, 
    37.40171, 37.51309, 37.62439, 37.7356, 37.84674,
  -11.83029, -11.72749, -11.6246, -11.5216, -11.41851, -11.31532, -11.21202, 
    -11.10863, -11.00514, -10.90156, -10.79787, -10.69408, -10.5902, 
    -10.48621, -10.38213, -10.27795, -10.17368, -10.0693, -9.964828, 
    -9.860257, -9.755589, -9.650825, -9.545962, -9.441003, -9.335946, 
    -9.230793, -9.125544, -9.020198, -8.914756, -8.809217, -8.703584, 
    -8.597854, -8.492028, -8.386107, -8.280091, -8.173981, -8.067774, 
    -7.961473, -7.855078, -7.748589, -7.642004, -7.535327, -7.428555, 
    -7.32169, -7.214731, -7.107679, -7.000535, -6.893297, -6.785967, 
    -6.678544, -6.571029, -6.463422, -6.355724, -6.247934, -6.140052, 
    -6.03208, -5.924016, -5.815862, -5.707617, -5.599283, -5.490858, 
    -5.382343, -5.273739, -5.165046, -5.056264, -4.947393, -4.838433, 
    -4.729385, -4.620249, -4.511025, -4.401714, -4.292316, -4.18283, 
    -4.073258, -3.963599, -3.853854, -3.744023, -3.634107, -3.524105, 
    -3.414017, -3.303845, -3.193589, -3.083248, -2.972823, -2.862315, 
    -2.751723, -2.641048, -2.53029, -2.419449, -2.308527, -2.197522, 
    -2.086436, -1.975268, -1.86402, -1.752691, -1.641281, -1.529792, 
    -1.418222, -1.306574, -1.194846, -1.083039, -0.971154, -0.8591908, 
    -0.7471499, -0.6350315, -0.522836, -0.4105638, -0.2982151, -0.1857904, 
    -0.07328991, 0.03928592, 0.1519368, 0.2646623, 0.3774621, 0.490336, 
    0.6032833, 0.716304, 0.8293975, 0.9425635, 1.055802, 1.169111, 1.282493, 
    1.395945, 1.509468, 1.623061, 1.736724, 1.850457, 1.964258, 2.078129, 
    2.192067, 2.306074, 2.420148, 2.534289, 2.648497, 2.762771, 2.877111, 
    2.991517, 3.105987, 3.220523, 3.335122, 3.449786, 3.564513, 3.679303, 
    3.794156, 3.90907, 4.024047, 4.139085, 4.254183, 4.369343, 4.484562, 
    4.599841, 4.715178, 4.830575, 4.94603, 5.061543, 5.177113, 5.29274, 
    5.408424, 5.524164, 5.639959, 5.755809, 5.871714, 5.987673, 6.103686, 
    6.219753, 6.335872, 6.452044, 6.568267, 6.684542, 6.800867, 6.917243, 
    7.03367, 7.150146, 7.26667, 7.383244, 7.499865, 7.616534, 7.733251, 
    7.850013, 7.966822, 8.083677, 8.200577, 8.317521, 8.43451, 8.551542, 
    8.668617, 8.785736, 8.902896, 9.020099, 9.137341, 9.254625, 9.371949, 
    9.489313, 9.606716, 9.724157, 9.841638, 9.959154, 10.07671, 10.1943, 
    10.31193, 10.42959, 10.54729, 10.66502, 10.78279, 10.90059, 11.01842, 
    11.13628, 11.25418, 11.37211, 11.49007, 11.60806, 11.72607, 11.84412, 
    11.9622, 12.0803, 12.19844, 12.3166, 12.43478, 12.553, 12.67123, 12.7895, 
    12.90778, 13.02609, 13.14443, 13.26279, 13.38116, 13.49957, 13.61799, 
    13.73643, 13.85489, 13.97338, 14.09188, 14.2104, 14.32893, 14.44749, 
    14.56606, 14.68465, 14.80325, 14.92187, 15.0405, 15.15915, 15.27781, 
    15.39648, 15.51516, 15.63386, 15.75257, 15.87129, 15.99002, 16.10875, 
    16.2275, 16.34626, 16.46502, 16.58379, 16.70257, 16.82135, 16.94014, 
    17.05893, 17.17773, 17.29653, 17.41534, 17.53415, 17.65296, 17.77177, 
    17.89058, 18.0094, 18.12821, 18.24702, 18.36584, 18.48465, 18.60345, 
    18.72226, 18.84106, 18.95986, 19.07865, 19.19744, 19.31622, 19.435, 
    19.55377, 19.67253, 19.79128, 19.91003, 20.02877, 20.14749, 20.26621, 
    20.38492, 20.50361, 20.62229, 20.74096, 20.85962, 20.97827, 21.0969, 
    21.21551, 21.33411, 21.4527, 21.57127, 21.68982, 21.80835, 21.92687, 
    22.04537, 22.16385, 22.28231, 22.40075, 22.51917, 22.63756, 22.75594, 
    22.87429, 22.99262, 23.11093, 23.22921, 23.34747, 23.46571, 23.58391, 
    23.7021, 23.82025, 23.93838, 24.05648, 24.17455, 24.2926, 24.41061, 
    24.52859, 24.64655, 24.76447, 24.88236, 25.00023, 25.11805, 25.23585, 
    25.35361, 25.47133, 25.58903, 25.70668, 25.8243, 25.94189, 26.05944, 
    26.17695, 26.29442, 26.41186, 26.52925, 26.64661, 26.76393, 26.88121, 
    26.99844, 27.11564, 27.23279, 27.34991, 27.46697, 27.584, 27.70098, 
    27.81792, 27.93481, 28.05166, 28.16846, 28.28522, 28.40192, 28.51859, 
    28.6352, 28.75177, 28.86828, 28.98475, 29.10117, 29.21754, 29.33385, 
    29.45012, 29.56634, 29.6825, 29.79861, 29.91467, 30.03067, 30.14662, 
    30.26252, 30.37836, 30.49415, 30.60988, 30.72555, 30.84117, 30.95673, 
    31.07224, 31.18768, 31.30307, 31.4184, 31.53367, 31.64888, 31.76403, 
    31.87912, 31.99414, 32.10911, 32.22402, 32.33886, 32.45364, 32.56836, 
    32.68301, 32.7976, 32.91212, 33.02658, 33.14098, 33.25531, 33.36958, 
    33.48377, 33.5979, 33.71196, 33.82596, 33.93989, 34.05375, 34.16754, 
    34.28126, 34.39491, 34.5085, 34.62201, 34.73545, 34.84882, 34.96212, 
    35.07534, 35.1885, 35.30158, 35.41459, 35.52752, 35.64038, 35.75317, 
    35.86589, 35.97853, 36.09109, 36.20358, 36.31599, 36.42833, 36.54059, 
    36.65277, 36.76488, 36.87691, 36.98886, 37.10073, 37.21252, 37.32424, 
    37.43587, 37.54743, 37.65891, 37.77031, 37.88162,
  -11.87998, -11.77705, -11.67401, -11.57088, -11.46764, -11.36431, 
    -11.26088, -11.15735, -11.05371, -10.94998, -10.84615, -10.74222, 
    -10.6382, -10.53407, -10.42984, -10.32552, -10.2211, -10.11657, 
    -10.01195, -9.907237, -9.802422, -9.697509, -9.592499, -9.487391, 
    -9.382186, -9.276883, -9.171484, -9.065988, -8.960395, -8.854706, 
    -8.74892, -8.643038, -8.53706, -8.430986, -8.324817, -8.218553, 
    -8.112192, -8.005736, -7.899186, -7.792541, -7.685801, -7.578967, 
    -7.472039, -7.365016, -7.2579, -7.15069, -7.043387, -6.93599, -6.828501, 
    -6.720918, -6.613243, -6.505476, -6.397616, -6.289664, -6.181621, 
    -6.073486, -5.96526, -5.856942, -5.748534, -5.640035, -5.531446, 
    -5.422766, -5.313997, -5.205138, -5.096189, -4.987151, -4.878025, 
    -4.768809, -4.659505, -4.550113, -4.440633, -4.331065, -4.22141, 
    -4.111668, -4.001839, -3.891923, -3.78192, -3.671832, -3.561658, 
    -3.451398, -3.341053, -3.230623, -3.120109, -3.00951, -2.898826, 
    -2.788059, -2.677209, -2.566275, -2.455258, -2.344159, -2.232977, 
    -2.121714, -2.010368, -1.898942, -1.787434, -1.675845, -1.564176, 
    -1.452427, -1.340598, -1.228689, -1.116701, -1.004635, -0.8924897, 
    -0.7802664, -0.6679654, -0.5555868, -0.4431311, -0.3305986, -0.2179896, 
    -0.1053045, 0.007456293, 0.1202925, 0.2332038, 0.3461898, 0.4592502, 
    0.5723845, 0.6855924, 0.7988735, 0.9122276, 1.025654, 1.139153, 1.252723, 
    1.366365, 1.480078, 1.593861, 1.707715, 1.821638, 1.935631, 2.049693, 
    2.163824, 2.278023, 2.392289, 2.506624, 2.621025, 2.735493, 2.850027, 
    2.964627, 3.079293, 3.194023, 3.308818, 3.423678, 3.538601, 3.653587, 
    3.768637, 3.883749, 3.998923, 4.114159, 4.229455, 4.344813, 4.460231, 
    4.575709, 4.691246, 4.806843, 4.922498, 5.038211, 5.153982, 5.26981, 
    5.385695, 5.501636, 5.617633, 5.733685, 5.849792, 5.965955, 6.08217, 
    6.19844, 6.314763, 6.431138, 6.547566, 6.664045, 6.780575, 6.897157, 
    7.013788, 7.130469, 7.2472, 7.363979, 7.480807, 7.597682, 7.714606, 
    7.831575, 7.948592, 8.065654, 8.182761, 8.299914, 8.417111, 8.534352, 
    8.651636, 8.768964, 8.886333, 9.003744, 9.121198, 9.238691, 9.356225, 
    9.4738, 9.591413, 9.709065, 9.826756, 9.944485, 10.06225, 10.18005, 
    10.29789, 10.41577, 10.53368, 10.65162, 10.7696, 10.88761, 11.00566, 
    11.12373, 11.24184, 11.35999, 11.47816, 11.59636, 11.71459, 11.83286, 
    11.95115, 12.06947, 12.18781, 12.30619, 12.42459, 12.54302, 12.66147, 
    12.77995, 12.89845, 13.01698, 13.13553, 13.2541, 13.3727, 13.49131, 
    13.60995, 13.72861, 13.84729, 13.96599, 14.08471, 14.20344, 14.3222, 
    14.44097, 14.55976, 14.67856, 14.79738, 14.91622, 15.03507, 15.15393, 
    15.27281, 15.3917, 15.5106, 15.62951, 15.74844, 15.86738, 15.98632, 
    16.10528, 16.22425, 16.34322, 16.4622, 16.58119, 16.70018, 16.81919, 
    16.93819, 17.0572, 17.17622, 17.29524, 17.41426, 17.53329, 17.65232, 
    17.77135, 17.89038, 18.00941, 18.12845, 18.24748, 18.36651, 18.48554, 
    18.60456, 18.72359, 18.84261, 18.96162, 19.08063, 19.19964, 19.31864, 
    19.43764, 19.55662, 19.6756, 19.79457, 19.91354, 20.03249, 20.15144, 
    20.27037, 20.3893, 20.50821, 20.62711, 20.746, 20.86487, 20.98374, 
    21.10258, 21.22142, 21.34023, 21.45904, 21.57782, 21.69659, 21.81534, 
    21.93407, 22.05279, 22.17149, 22.29016, 22.40882, 22.52745, 22.64606, 
    22.76466, 22.88323, 23.00177, 23.12029, 23.23879, 23.35727, 23.47572, 
    23.59414, 23.71254, 23.83091, 23.94925, 24.06757, 24.18585, 24.30411, 
    24.42234, 24.54054, 24.6587, 24.77684, 24.89495, 25.01302, 25.13106, 
    25.24907, 25.36704, 25.48498, 25.60288, 25.72075, 25.83858, 25.95638, 
    26.07414, 26.19186, 26.30955, 26.42719, 26.5448, 26.66237, 26.7799, 
    26.89738, 27.01483, 27.13224, 27.2496, 27.36692, 27.4842, 27.60143, 
    27.71862, 27.83577, 27.95287, 28.06992, 28.18693, 28.30389, 28.42081, 
    28.53768, 28.6545, 28.77127, 28.88799, 29.00467, 29.12129, 29.23786, 
    29.35438, 29.47086, 29.58727, 29.70364, 29.81996, 29.93622, 30.05242, 
    30.16858, 30.28468, 30.40072, 30.51671, 30.63264, 30.74852, 30.86434, 
    30.9801, 31.0958, 31.21145, 31.32703, 31.44256, 31.55803, 31.67344, 
    31.78879, 31.90407, 32.0193, 32.13446, 32.24957, 32.3646, 32.47958, 
    32.59449, 32.70934, 32.82413, 32.93885, 33.0535, 33.16809, 33.28262, 
    33.39708, 33.51147, 33.62579, 33.74005, 33.85423, 33.96835, 34.08241, 
    34.19639, 34.3103, 34.42414, 34.53791, 34.65162, 34.76525, 34.87881, 
    34.99229, 35.10571, 35.21905, 35.33232, 35.44552, 35.55864, 35.67169, 
    35.78466, 35.89756, 36.01039, 36.12313, 36.23581, 36.3484, 36.46093, 
    36.57337, 36.68573, 36.79802, 36.91024, 37.02237, 37.13442, 37.2464, 
    37.35829, 37.47011, 37.58184, 37.6935, 37.80508, 37.91657,
  -11.92975, -11.82668, -11.72351, -11.62023, -11.51686, -11.41339, 
    -11.30981, -11.20614, -11.10236, -10.99849, -10.89452, -10.79044, 
    -10.68627, -10.582, -10.47763, -10.37316, -10.26859, -10.16392, 
    -10.05916, -9.954294, -9.849332, -9.744271, -9.639112, -9.533856, 
    -9.428502, -9.32305, -9.217502, -9.111855, -9.006111, -8.90027, 
    -8.794333, -8.688299, -8.582169, -8.475943, -8.369619, -8.263201, 
    -8.156686, -8.050076, -7.94337, -7.83657, -7.729674, -7.622684, 
    -7.515598, -7.408418, -7.301145, -7.193776, -7.086314, -6.978759, 
    -6.871109, -6.763367, -6.655532, -6.547604, -6.439582, -6.331469, 
    -6.223264, -6.114966, -6.006577, -5.898096, -5.789524, -5.680861, 
    -5.572107, -5.463262, -5.354327, -5.245302, -5.136188, -5.026983, 
    -4.917689, -4.808306, -4.698833, -4.589273, -4.479624, -4.369887, 
    -4.260062, -4.150149, -4.040149, -3.930062, -3.819889, -3.709628, 
    -3.599282, -3.488849, -3.378331, -3.267728, -3.157039, -3.046266, 
    -2.935407, -2.824465, -2.713439, -2.602329, -2.491136, -2.37986, 
    -2.268501, -2.157059, -2.045536, -1.933931, -1.822244, -1.710476, 
    -1.598627, -1.486697, -1.374688, -1.262598, -1.150429, -1.038181, 
    -0.9258537, -0.8134479, -0.7009639, -0.588402, -0.4757626, -0.363046, 
    -0.2502525, -0.1373825, -0.02443641, 0.0885855, 0.2016828, 0.3148553, 
    0.4281024, 0.5414239, 0.6548194, 0.7682884, 0.8818308, 0.995446, 
    1.109134, 1.222894, 1.336725, 1.450628, 1.564602, 1.678647, 1.792761, 
    1.906946, 2.0212, 2.135523, 2.249914, 2.364374, 2.478902, 2.593497, 
    2.708159, 2.822888, 2.937682, 3.052543, 3.167469, 3.28246, 3.397516, 
    3.512635, 3.627819, 3.743065, 3.858375, 3.973747, 4.08918, 4.204676, 
    4.320232, 4.435849, 4.551527, 4.667264, 4.78306, 4.898916, 5.014829, 
    5.130801, 5.24683, 5.362917, 5.47906, 5.595259, 5.711514, 5.827825, 
    5.94419, 6.060609, 6.177083, 6.293609, 6.410189, 6.526821, 6.643505, 
    6.76024, 6.877027, 6.993864, 7.110751, 7.227688, 7.344674, 7.461708, 
    7.578791, 7.695921, 7.813098, 7.930322, 8.047592, 8.164908, 8.282269, 
    8.399674, 8.517124, 8.634618, 8.752154, 8.869734, 8.987355, 9.105019, 
    9.222723, 9.340467, 9.458252, 9.576077, 9.69394, 9.811842, 9.929782, 
    10.04776, 10.16577, 10.28382, 10.40191, 10.52003, 10.63819, 10.75638, 
    10.87461, 10.99287, 11.11116, 11.22948, 11.34784, 11.46623, 11.58464, 
    11.70309, 11.82157, 11.94007, 12.05861, 12.17717, 12.29576, 12.41438, 
    12.53302, 12.65169, 12.77038, 12.8891, 13.00784, 13.12661, 13.2454, 
    13.36421, 13.48304, 13.6019, 13.72077, 13.83967, 13.95858, 14.07752, 
    14.19647, 14.31544, 14.43443, 14.55344, 14.67246, 14.7915, 14.91055, 
    15.02962, 15.1487, 15.2678, 15.38691, 15.50603, 15.62516, 15.7443, 
    15.86346, 15.98262, 16.1018, 16.22098, 16.34017, 16.45937, 16.57858, 
    16.69779, 16.81701, 16.93624, 17.05547, 17.17471, 17.29395, 17.41319, 
    17.53243, 17.65168, 17.77093, 17.89018, 18.00943, 18.12868, 18.24793, 
    18.36718, 18.48643, 18.60567, 18.72492, 18.84416, 18.96339, 19.08262, 
    19.20185, 19.32106, 19.44028, 19.55948, 19.67868, 19.79787, 19.91706, 
    20.03623, 20.15539, 20.27454, 20.39369, 20.51282, 20.63194, 20.75104, 
    20.87014, 20.98922, 21.10828, 21.22733, 21.34637, 21.46539, 21.58439, 
    21.70338, 21.82235, 21.9413, 22.06023, 22.17914, 22.29803, 22.4169, 
    22.53576, 22.65459, 22.7734, 22.89218, 23.01094, 23.12968, 23.2484, 
    23.36709, 23.48575, 23.60439, 23.723, 23.84159, 23.96015, 24.07867, 
    24.19718, 24.31565, 24.43409, 24.5525, 24.67089, 24.78924, 24.90755, 
    25.02584, 25.14409, 25.26231, 25.3805, 25.49865, 25.61677, 25.73485, 
    25.8529, 25.97091, 26.08888, 26.20681, 26.32471, 26.44256, 26.56038, 
    26.67816, 26.7959, 26.9136, 27.03125, 27.14887, 27.26644, 27.38397, 
    27.50146, 27.6189, 27.7363, 27.85365, 27.97096, 28.08822, 28.20544, 
    28.32261, 28.43973, 28.55681, 28.67384, 28.79081, 28.90774, 29.02462, 
    29.14145, 29.25823, 29.37496, 29.49163, 29.60826, 29.72483, 29.84134, 
    29.95781, 30.07422, 30.19058, 30.30688, 30.42313, 30.53932, 30.65545, 
    30.77153, 30.88755, 31.00351, 31.11942, 31.23526, 31.35105, 31.46678, 
    31.58244, 31.69805, 31.8136, 31.92908, 32.04451, 32.15987, 32.27517, 
    32.39041, 32.50558, 32.62069, 32.73573, 32.85072, 32.96563, 33.08048, 
    33.19527, 33.30998, 33.42463, 33.53922, 33.65374, 33.76818, 33.88256, 
    33.99688, 34.11112, 34.2253, 34.3394, 34.45343, 34.56739, 34.68129, 
    34.7951, 34.90886, 35.02253, 35.13614, 35.24966, 35.36312, 35.47651, 
    35.58982, 35.70305, 35.81621, 35.9293, 36.04231, 36.15524, 36.2681, 
    36.38088, 36.49359, 36.60621, 36.71876, 36.83123, 36.94363, 37.05594, 
    37.16818, 37.28033, 37.39241, 37.50441, 37.61633, 37.72816, 37.83992, 
    37.95159,
  -11.97961, -11.87639, -11.77308, -11.66967, -11.56615, -11.46254, 
    -11.35882, -11.25501, -11.15109, -11.04707, -10.94296, -10.83874, 
    -10.73443, -10.63001, -10.52549, -10.42088, -10.31617, -10.21135, 
    -10.10644, -10.00143, -9.89632, -9.791112, -9.685805, -9.5804, -9.474896, 
    -9.369295, -9.263597, -9.1578, -9.051905, -8.945913, -8.839824, 
    -8.733638, -8.627355, -8.520975, -8.414499, -8.307926, -8.201258, 
    -8.094493, -7.987632, -7.880675, -7.773623, -7.666476, -7.559234, 
    -7.451897, -7.344465, -7.236938, -7.129318, -7.021603, -6.913794, 
    -6.805892, -6.697896, -6.589807, -6.481625, -6.373349, -6.264981, 
    -6.156521, -6.047969, -5.939325, -5.830589, -5.721761, -5.612842, 
    -5.503832, -5.394732, -5.285541, -5.176259, -5.066887, -4.957426, 
    -4.847875, -4.738235, -4.628505, -4.518687, -4.408781, -4.298786, 
    -4.188703, -4.078532, -3.968274, -3.857928, -3.747496, -3.636977, 
    -3.526371, -3.41568, -3.304902, -3.19404, -3.083091, -2.972058, 
    -2.860941, -2.749738, -2.638452, -2.527082, -2.415629, -2.304093, 
    -2.192473, -2.080771, -1.968987, -1.857121, -1.745174, -1.633145, 
    -1.521035, -1.408845, -1.296574, -1.184223, -1.071793, -0.9592832, 
    -0.8466946, -0.7340274, -0.621282, -0.5084586, -0.3955576, -0.2825794, 
    -0.1695242, -0.05639258, 0.05681526, 0.1700989, 0.2834581, 0.3968923, 
    0.5104012, 0.6239846, 0.7376419, 0.8513728, 0.965177, 1.079054, 1.193004, 
    1.307025, 1.421119, 1.535284, 1.649519, 1.763826, 1.878202, 1.992648, 
    2.107164, 2.221748, 2.336402, 2.451123, 2.565912, 2.680769, 2.795692, 
    2.910682, 3.025738, 3.14086, 3.256047, 3.371299, 3.486616, 3.601996, 
    3.71744, 3.832948, 3.948518, 4.06415, 4.179844, 4.2956, 4.411417, 
    4.527294, 4.643231, 4.759228, 4.875284, 4.991399, 5.107572, 5.223803, 
    5.340091, 5.456437, 5.572839, 5.689297, 5.80581, 5.922379, 6.039002, 
    6.155679, 6.27241, 6.389194, 6.506031, 6.622921, 6.739861, 6.856854, 
    6.973897, 7.090991, 7.208134, 7.325326, 7.442568, 7.559858, 7.677196, 
    7.794581, 7.912013, 8.029491, 8.147017, 8.264586, 8.382201, 8.49986, 
    8.617563, 8.73531, 8.853099, 8.97093, 9.088804, 9.206719, 9.324675, 
    9.442671, 9.560707, 9.678782, 9.796896, 9.915048, 10.03324, 10.15146, 
    10.26973, 10.38803, 10.50636, 10.62473, 10.74314, 10.86158, 10.98005, 
    11.09856, 11.21709, 11.33566, 11.45427, 11.5729, 11.69156, 11.81025, 
    11.92897, 12.04772, 12.1665, 12.28531, 12.40414, 12.523, 12.64188, 
    12.76079, 12.87973, 12.99869, 13.11767, 13.23667, 13.3557, 13.47475, 
    13.59383, 13.71292, 13.83203, 13.95117, 14.07032, 14.18949, 14.30868, 
    14.42788, 14.54711, 14.66635, 14.7856, 14.90488, 15.02416, 15.14346, 
    15.26278, 15.3821, 15.50144, 15.62079, 15.74016, 15.85953, 15.97891, 
    16.09831, 16.21771, 16.33712, 16.45654, 16.57597, 16.6954, 16.81484, 
    16.93428, 17.05373, 17.17319, 17.29265, 17.41211, 17.53157, 17.65104, 
    17.77051, 17.88998, 18.00945, 18.12892, 18.24839, 18.36786, 18.48732, 
    18.60679, 18.72625, 18.84571, 18.96516, 19.08461, 19.20406, 19.32349, 
    19.44293, 19.56235, 19.68177, 19.80118, 19.92058, 20.03997, 20.15935, 
    20.27873, 20.39809, 20.51744, 20.63677, 20.7561, 20.87541, 20.99471, 
    21.11399, 21.23326, 21.35251, 21.47175, 21.59097, 21.71018, 21.82936, 
    21.94853, 22.06768, 22.18681, 22.30592, 22.42501, 22.54408, 22.66313, 
    22.78215, 22.90115, 23.02013, 23.13909, 23.25802, 23.37693, 23.49581, 
    23.61466, 23.73349, 23.85229, 23.97106, 24.08981, 24.20852, 24.32721, 
    24.44587, 24.5645, 24.68309, 24.80166, 24.92019, 25.03869, 25.15716, 
    25.27559, 25.39399, 25.51236, 25.63069, 25.74898, 25.86724, 25.98546, 
    26.10365, 26.22179, 26.3399, 26.45797, 26.576, 26.69399, 26.81194, 
    26.92984, 27.04771, 27.16554, 27.28332, 27.40106, 27.51875, 27.63641, 
    27.75401, 27.87158, 27.98909, 28.10657, 28.22399, 28.34137, 28.4587, 
    28.57598, 28.69321, 28.8104, 28.92754, 29.04462, 29.16166, 29.27864, 
    29.39557, 29.51245, 29.62928, 29.74606, 29.86278, 29.97945, 30.09606, 
    30.21262, 30.32913, 30.44558, 30.56197, 30.67831, 30.79459, 30.91081, 
    31.02697, 31.14308, 31.25912, 31.37511, 31.49104, 31.60691, 31.72272, 
    31.83846, 31.95415, 32.06977, 32.18533, 32.30083, 32.41626, 32.53163, 
    32.64693, 32.76218, 32.87735, 32.99247, 33.10751, 33.22249, 33.33741, 
    33.45225, 33.56703, 33.68174, 33.79638, 33.91095, 34.02546, 34.1399, 
    34.25426, 34.36856, 34.48278, 34.59694, 34.71102, 34.82503, 34.93896, 
    35.05283, 35.16662, 35.28034, 35.39399, 35.50756, 35.62106, 35.73448, 
    35.84782, 35.9611, 36.0743, 36.18741, 36.30046, 36.41342, 36.52631, 
    36.63912, 36.75185, 36.86451, 36.97709, 37.08958, 37.202, 37.31434, 
    37.4266, 37.53877, 37.65087, 37.76289, 37.87482, 37.98668,
  -12.02954, -11.92619, -11.82273, -11.71918, -11.61553, -11.51177, 
    -11.40791, -11.30396, -11.1999, -11.09574, -10.99148, -10.88712, 
    -10.78266, -10.6781, -10.57344, -10.46868, -10.36382, -10.25886, 
    -10.1538, -10.04865, -9.943387, -9.838031, -9.732576, -9.627022, 
    -9.52137, -9.415619, -9.30977, -9.203822, -9.097777, -8.991633, 
    -8.885393, -8.779055, -8.672619, -8.566086, -8.459456, -8.35273, 
    -8.245906, -8.138987, -8.03197, -7.924858, -7.81765, -7.710346, 
    -7.602947, -7.495452, -7.387862, -7.280177, -7.172398, -7.064524, 
    -6.956555, -6.848493, -6.740336, -6.632086, -6.523742, -6.415305, 
    -6.306775, -6.198152, -6.089436, -5.980628, -5.871728, -5.762736, 
    -5.653652, -5.544477, -5.43521, -5.325853, -5.216404, -5.106866, 
    -4.997237, -4.887518, -4.777709, -4.667811, -4.557823, -4.447747, 
    -4.337582, -4.227328, -4.116986, -4.006557, -3.896039, -3.785435, 
    -3.674743, -3.563964, -3.453099, -3.342148, -3.231111, -3.119987, 
    -3.008779, -2.897486, -2.786108, -2.674645, -2.563098, -2.451468, 
    -2.339753, -2.227956, -2.116075, -2.004112, -1.892067, -1.779939, 
    -1.66773, -1.55544, -1.443068, -1.330616, -1.218084, -1.105471, 
    -0.9927788, -0.8800071, -0.7671565, -0.6542272, -0.5412195, -0.4281339, 
    -0.3149706, -0.2017301, -0.08841263, 0.02498142, 0.1384517, 0.2519978, 
    0.3656194, 0.4793161, 0.5930876, 0.7069334, 0.8208532, 0.9348467, 
    1.048913, 1.163053, 1.277265, 1.391549, 1.505905, 1.620332, 1.734831, 
    1.849399, 1.964038, 2.078747, 2.193525, 2.308372, 2.423287, 2.53827, 
    2.653322, 2.76844, 2.883626, 2.998878, 3.114196, 3.229579, 3.345028, 
    3.460542, 3.57612, 3.691762, 3.807467, 3.923236, 4.039067, 4.154961, 
    4.270916, 4.386932, 4.503009, 4.619147, 4.735345, 4.851602, 4.967918, 
    5.084293, 5.200727, 5.317217, 5.433765, 5.55037, 5.667031, 5.783748, 
    5.900521, 6.017348, 6.13423, 6.251166, 6.368155, 6.485197, 6.602292, 
    6.719439, 6.836637, 6.953887, 7.071187, 7.188538, 7.305937, 7.423387, 
    7.540884, 7.65843, 7.776023, 7.893664, 8.011352, 8.129086, 8.246864, 
    8.364689, 8.482557, 8.600471, 8.718428, 8.836428, 8.95447, 9.072555, 
    9.190681, 9.308847, 9.427055, 9.545303, 9.66359, 9.781917, 9.900281, 
    10.01868, 10.13712, 10.2556, 10.37411, 10.49266, 10.61125, 10.72987, 
    10.84852, 10.96721, 11.08593, 11.20468, 11.32346, 11.44228, 11.56113, 
    11.68, 11.79891, 11.91785, 12.03681, 12.15581, 12.27483, 12.39388, 
    12.51295, 12.63205, 12.75118, 12.87033, 12.98951, 13.10871, 13.22793, 
    13.34718, 13.46645, 13.58574, 13.70505, 13.82438, 13.94373, 14.0631, 
    14.18249, 14.3019, 14.42132, 14.54076, 14.66022, 14.7797, 14.89919, 
    15.01869, 15.13821, 15.25774, 15.37729, 15.49685, 15.61642, 15.736, 
    15.85559, 15.9752, 16.09481, 16.21443, 16.33406, 16.4537, 16.57335, 
    16.693, 16.81266, 16.93232, 17.05199, 17.17167, 17.29135, 17.41103, 
    17.53071, 17.6504, 17.77009, 17.88978, 18.00947, 18.12916, 18.24885, 
    18.36853, 18.48822, 18.6079, 18.72759, 18.84727, 18.96694, 19.08661, 
    19.20627, 19.32593, 19.44558, 19.56523, 19.68486, 19.80449, 19.92411, 
    20.04372, 20.16333, 20.28292, 20.4025, 20.52207, 20.64162, 20.76117, 
    20.8807, 21.00021, 21.11972, 21.2392, 21.35868, 21.47813, 21.59757, 
    21.717, 21.8364, 21.95579, 22.07515, 22.1945, 22.31383, 22.43314, 
    22.55242, 22.67169, 22.79093, 22.91015, 23.02934, 23.14852, 23.26766, 
    23.38679, 23.50588, 23.62496, 23.744, 23.86302, 23.98201, 24.10097, 
    24.2199, 24.3388, 24.45768, 24.57652, 24.69533, 24.81411, 24.93286, 
    25.05157, 25.17025, 25.2889, 25.40751, 25.52609, 25.64464, 25.76314, 
    25.88161, 26.00005, 26.11844, 26.2368, 26.35512, 26.4734, 26.59165, 
    26.70985, 26.82801, 26.94613, 27.06421, 27.18224, 27.30023, 27.41818, 
    27.53609, 27.65395, 27.77177, 27.88954, 28.00727, 28.12495, 28.24258, 
    28.36017, 28.47771, 28.5952, 28.71264, 28.83003, 28.94737, 29.06466, 
    29.18191, 29.2991, 29.41623, 29.53332, 29.65035, 29.76734, 29.88426, 
    30.00114, 30.11795, 30.23472, 30.35143, 30.46808, 30.58467, 30.70121, 
    30.8177, 30.93412, 31.05049, 31.16679, 31.28304, 31.39923, 31.51536, 
    31.63142, 31.74743, 31.86338, 31.97926, 32.09508, 32.21084, 32.32653, 
    32.44217, 32.55774, 32.67324, 32.78868, 32.90405, 33.01936, 33.1346, 
    33.24977, 33.36488, 33.47992, 33.59489, 33.7098, 33.82463, 33.9394, 
    34.0541, 34.16873, 34.28329, 34.39777, 34.51219, 34.62653, 34.74081, 
    34.85501, 34.96914, 35.08319, 35.19717, 35.31108, 35.42492, 35.53867, 
    35.65236, 35.76597, 35.8795, 35.99296, 36.10634, 36.21965, 36.33288, 
    36.44603, 36.5591, 36.6721, 36.78501, 36.89785, 37.01061, 37.12329, 
    37.23589, 37.34841, 37.46085, 37.57321, 37.68549, 37.79768, 37.9098, 
    38.02183,
  -12.07955, -11.97606, -11.87247, -11.76877, -11.66498, -11.56108, 
    -11.45708, -11.35298, -11.24878, -11.14448, -11.04008, -10.93558, 
    -10.83097, -10.72627, -10.62146, -10.51656, -10.41155, -10.30645, 
    -10.20124, -10.09594, -9.990534, -9.88503, -9.779426, -9.673723, 
    -9.567922, -9.462021, -9.356022, -9.249924, -9.143727, -9.037433, 
    -8.93104, -8.82455, -8.717961, -8.611275, -8.504492, -8.397611, 
    -8.290632, -8.183558, -8.076386, -7.969118, -7.861754, -7.754293, 
    -7.646737, -7.539084, -7.431336, -7.323493, -7.215554, -7.107521, 
    -6.999393, -6.89117, -6.782852, -6.674441, -6.565936, -6.457336, 
    -6.348644, -6.239858, -6.130979, -6.022007, -5.912942, -5.803786, 
    -5.694537, -5.585196, -5.475763, -5.36624, -5.256624, -5.146918, 
    -5.037122, -4.927235, -4.817257, -4.70719, -4.597033, -4.486786, 
    -4.376451, -4.266026, -4.155514, -4.044912, -3.934223, -3.823446, 
    -3.712581, -3.601629, -3.49059, -3.379465, -3.268253, -3.156955, 
    -3.045571, -2.934102, -2.822547, -2.710908, -2.599184, -2.487375, 
    -2.375483, -2.263507, -2.151448, -2.039306, -1.927081, -1.814773, 
    -1.702384, -1.589912, -1.477359, -1.364726, -1.252011, -1.139216, 
    -1.026341, -0.9133858, -0.8003514, -0.687238, -0.5740459, -0.4607753, 
    -0.3474268, -0.2340005, -0.120497, -0.006916431, 0.1067407, 0.2204741, 
    0.3342833, 0.4481681, 0.5621279, 0.6761626, 0.7902716, 0.9044546, 
    1.018711, 1.133041, 1.247444, 1.361919, 1.476467, 1.591086, 1.705776, 
    1.820537, 1.935369, 2.050271, 2.165243, 2.280283, 2.395393, 2.510572, 
    2.625818, 2.741132, 2.856513, 2.971961, 3.087476, 3.203056, 3.318702, 
    3.434414, 3.550189, 3.66603, 3.781934, 3.897901, 4.013931, 4.130024, 
    4.24618, 4.362396, 4.478674, 4.595012, 4.711411, 4.82787, 4.944388, 
    5.060965, 5.177601, 5.294294, 5.411046, 5.527853, 5.644719, 5.76164, 
    5.878616, 5.995648, 6.112735, 6.229876, 6.34707, 6.464318, 6.581619, 
    6.698972, 6.816377, 6.933834, 7.051341, 7.168899, 7.286506, 7.404163, 
    7.521869, 7.639624, 7.757426, 7.875276, 7.993172, 8.111115, 8.229104, 
    8.347138, 8.465218, 8.583341, 8.701509, 8.819719, 8.937973, 9.056269, 
    9.174606, 9.292986, 9.411406, 9.529865, 9.648365, 9.766904, 9.885482, 
    10.0041, 10.12275, 10.24144, 10.36017, 10.47893, 10.59773, 10.71656, 
    10.83543, 10.95433, 11.07327, 11.19223, 11.31123, 11.43027, 11.54933, 
    11.66842, 11.78755, 11.9067, 12.02588, 12.14509, 12.26433, 12.38359, 
    12.50289, 12.6222, 12.74155, 12.86092, 12.98031, 13.09973, 13.21917, 
    13.33863, 13.45812, 13.57763, 13.69716, 13.81671, 13.93627, 14.05586, 
    14.17547, 14.2951, 14.41474, 14.5344, 14.65408, 14.77377, 14.89348, 
    15.01321, 15.13295, 15.2527, 15.37246, 15.49224, 15.61203, 15.73183, 
    15.85165, 15.97147, 16.0913, 16.21115, 16.331, 16.45085, 16.57072, 
    16.69059, 16.81047, 16.93036, 17.05025, 17.17014, 17.29004, 17.40994, 
    17.52985, 17.64976, 17.76966, 17.88957, 18.00948, 18.12939, 18.2493, 
    18.36921, 18.48912, 18.60902, 18.72893, 18.84882, 18.96872, 19.08861, 
    19.20849, 19.32837, 19.44824, 19.56811, 19.68796, 19.80781, 19.92765, 
    20.04749, 20.1673, 20.28712, 20.40692, 20.5267, 20.64648, 20.76624, 
    20.886, 21.00573, 21.12545, 21.24516, 21.36485, 21.48453, 21.60419, 
    21.72383, 21.84345, 21.96305, 22.08264, 22.20221, 22.32175, 22.44128, 
    22.56078, 22.68027, 22.79973, 22.91916, 23.03858, 23.15797, 23.27733, 
    23.39667, 23.51599, 23.63527, 23.75454, 23.87377, 23.99297, 24.11215, 
    24.2313, 24.35042, 24.46951, 24.58857, 24.70759, 24.82659, 24.94555, 
    25.06448, 25.18337, 25.30224, 25.42106, 25.53986, 25.65862, 25.77734, 
    25.89602, 26.01467, 26.13328, 26.25185, 26.37038, 26.48888, 26.60733, 
    26.72574, 26.84412, 26.96245, 27.08074, 27.19898, 27.31719, 27.43535, 
    27.55346, 27.67154, 27.78956, 27.90755, 28.02548, 28.14337, 28.26121, 
    28.37901, 28.49675, 28.61445, 28.7321, 28.8497, 28.96725, 29.08475, 
    29.2022, 29.3196, 29.43694, 29.55423, 29.67147, 29.78866, 29.90579, 
    30.02287, 30.13989, 30.25686, 30.37377, 30.49063, 30.60743, 30.72417, 
    30.84085, 30.95748, 31.07405, 31.19056, 31.307, 31.4234, 31.53972, 
    31.65599, 31.7722, 31.88834, 32.00443, 32.12045, 32.2364, 32.3523, 
    32.46813, 32.58389, 32.6996, 32.81523, 32.9308, 33.04631, 33.16174, 
    33.27711, 33.39242, 33.50765, 33.62282, 33.73792, 33.85295, 33.96791, 
    34.0828, 34.19762, 34.31237, 34.42705, 34.54166, 34.65619, 34.77066, 
    34.88505, 34.99937, 35.11361, 35.22778, 35.34188, 35.4559, 35.56985, 
    35.68372, 35.79752, 35.91124, 36.02489, 36.13846, 36.25195, 36.36536, 
    36.4787, 36.59196, 36.70514, 36.81824, 36.93126, 37.0442, 37.15706, 
    37.26985, 37.38255, 37.49517, 37.60771, 37.72017, 37.83254, 37.94484, 
    38.05705,
  -12.12964, -12.02601, -11.92228, -11.81845, -11.71451, -11.61047, 
    -11.50633, -11.40209, -11.29775, -11.19331, -11.08876, -10.98411, 
    -10.87937, -10.77452, -10.66957, -10.56452, -10.45937, -10.35412, 
    -10.24876, -10.14331, -10.03776, -9.932107, -9.826355, -9.720504, 
    -9.614552, -9.508503, -9.402353, -9.296104, -9.189757, -9.083311, 
    -8.976767, -8.870123, -8.763382, -8.656543, -8.549605, -8.442571, 
    -8.335438, -8.228208, -8.120881, -8.013456, -7.905936, -7.798318, 
    -7.690605, -7.582794, -7.474888, -7.366886, -7.258789, -7.150596, 
    -7.042307, -6.933924, -6.825446, -6.716873, -6.608206, -6.499444, 
    -6.390589, -6.28164, -6.172597, -6.063462, -5.954233, -5.844912, 
    -5.735497, -5.62599, -5.516392, -5.406701, -5.296919, -5.187046, 
    -5.077081, -4.967025, -4.856879, -4.746643, -4.636316, -4.525899, 
    -4.415393, -4.304798, -4.194114, -4.083341, -3.972479, -3.861529, 
    -3.750491, -3.639366, -3.528153, -3.416853, -3.305466, -3.193993, 
    -3.082433, -2.970788, -2.859057, -2.747241, -2.635339, -2.523353, 
    -2.411283, -2.299128, -2.18689, -2.074568, -1.962163, -1.849675, 
    -1.737105, -1.624453, -1.511719, -1.398903, -1.286006, -1.173028, 
    -1.05997, -0.946831, -0.8336127, -0.7203149, -0.606938, -0.4934823, 
    -0.3799481, -0.2663359, -0.152646, -0.0388787, 0.07496558, 0.1888865, 
    0.3028837, 0.4169568, 0.5311053, 0.6453291, 0.7596276, 0.8740005, 
    0.9884474, 1.102968, 1.217562, 1.332228, 1.446968, 1.561779, 1.676662, 
    1.791616, 1.906641, 2.021736, 2.136902, 2.252137, 2.367442, 2.482815, 
    2.598257, 2.713767, 2.829344, 2.944988, 3.0607, 3.176477, 3.292321, 
    3.40823, 3.524204, 3.640243, 3.756346, 3.872513, 3.988743, 4.105035, 
    4.221391, 4.337808, 4.454287, 4.570827, 4.687427, 4.804087, 4.920808, 
    5.037587, 5.154426, 5.271322, 5.388277, 5.505289, 5.622357, 5.739483, 
    5.856664, 5.973901, 6.091193, 6.208539, 6.32594, 6.443394, 6.560901, 
    6.678461, 6.796073, 6.913737, 7.031452, 7.149217, 7.267033, 7.384898, 
    7.502813, 7.620776, 7.738787, 7.856846, 7.974953, 8.093105, 8.211305, 
    8.329549, 8.447839, 8.566174, 8.684552, 8.802975, 8.921439, 9.039948, 
    9.158497, 9.277088, 9.39572, 9.514394, 9.633106, 9.751859, 9.870649, 
    9.989479, 10.10835, 10.22725, 10.34619, 10.46517, 10.58418, 10.70323, 
    10.82231, 10.94143, 11.06058, 11.17976, 11.29898, 11.41823, 11.53751, 
    11.65681, 11.77615, 11.89552, 12.01492, 12.13435, 12.25381, 12.37329, 
    12.4928, 12.61233, 12.73189, 12.85148, 12.97109, 13.09073, 13.21039, 
    13.33007, 13.44977, 13.5695, 13.68925, 13.80902, 13.9288, 14.04861, 
    14.16844, 14.28829, 14.40815, 14.52803, 14.64793, 14.76784, 14.88777, 
    15.00771, 15.12767, 15.24764, 15.36763, 15.48763, 15.60764, 15.72766, 
    15.84769, 15.96774, 16.08779, 16.20785, 16.32792, 16.448, 16.56809, 
    16.68818, 16.80828, 16.92839, 17.0485, 17.16861, 17.28873, 17.40886, 
    17.52898, 17.64911, 17.76924, 17.88937, 18.0095, 18.12963, 18.24976, 
    18.36989, 18.49002, 18.61015, 18.73027, 18.85039, 18.9705, 19.09061, 
    19.21072, 19.33082, 19.45091, 19.57099, 19.69107, 19.81114, 19.9312, 
    20.05125, 20.1713, 20.29133, 20.41135, 20.53135, 20.65135, 20.77134, 
    20.89131, 21.01126, 21.1312, 21.25113, 21.37104, 21.49093, 21.61081, 
    21.73067, 21.85052, 21.97034, 22.09015, 22.20993, 22.32969, 22.44944, 
    22.56916, 22.68886, 22.80854, 22.9282, 23.04783, 23.16744, 23.28702, 
    23.40658, 23.52611, 23.64561, 23.76509, 23.88454, 24.00397, 24.12336, 
    24.24273, 24.36206, 24.48137, 24.60064, 24.71988, 24.83909, 24.95827, 
    25.07742, 25.19653, 25.3156, 25.43465, 25.55365, 25.67263, 25.79156, 
    25.91046, 26.02932, 26.14814, 26.26693, 26.38568, 26.50438, 26.62305, 
    26.74167, 26.86026, 26.9788, 27.0973, 27.21576, 27.33418, 27.45255, 
    27.57088, 27.68916, 27.8074, 27.92559, 28.04373, 28.16183, 28.27988, 
    28.39789, 28.51584, 28.63375, 28.75161, 28.86942, 28.98717, 29.10488, 
    29.22253, 29.34014, 29.45769, 29.57519, 29.69263, 29.81003, 29.92736, 
    30.04465, 30.16188, 30.27905, 30.39616, 30.51323, 30.63023, 30.74717, 
    30.86406, 30.98089, 31.09766, 31.21437, 31.33102, 31.44761, 31.56414, 
    31.68061, 31.79702, 31.91336, 32.02965, 32.14587, 32.26202, 32.37812, 
    32.49414, 32.61011, 32.72601, 32.84184, 32.95761, 33.07331, 33.18894, 
    33.30451, 33.42001, 33.53544, 33.6508, 33.76609, 33.88132, 33.99648, 
    34.11156, 34.22657, 34.34151, 34.45639, 34.57119, 34.68591, 34.80057, 
    34.91515, 35.02966, 35.1441, 35.25846, 35.37275, 35.48696, 35.60109, 
    35.71515, 35.82914, 35.94305, 36.05688, 36.17064, 36.28431, 36.39791, 
    36.51143, 36.62488, 36.73824, 36.85153, 36.96473, 37.07786, 37.19091, 
    37.30387, 37.41676, 37.52956, 37.64228, 37.75492, 37.86747, 37.97995, 
    38.09234,
  -12.17981, -12.07605, -11.97217, -11.8682, -11.76412, -11.65995, -11.55567, 
    -11.45128, -11.3468, -11.24221, -11.13752, -11.03273, -10.92784, 
    -10.82285, -10.71775, -10.61256, -10.50726, -10.40186, -10.29636, 
    -10.19077, -10.08506, -9.979265, -9.873364, -9.767365, -9.661264, 
    -9.555064, -9.448764, -9.342365, -9.235867, -9.129269, -9.022572, 
    -8.915776, -8.808882, -8.701889, -8.594798, -8.487609, -8.380322, 
    -8.272937, -8.165454, -8.057874, -7.950196, -7.842422, -7.73455, 
    -7.626583, -7.518518, -7.410357, -7.302101, -7.193748, -7.085299, 
    -6.976756, -6.868116, -6.759382, -6.650553, -6.541629, -6.432611, 
    -6.323499, -6.214293, -6.104993, -5.9956, -5.886113, -5.776533, 
    -5.666861, -5.557096, -5.447238, -5.337289, -5.227248, -5.117115, 
    -5.006891, -4.896576, -4.78617, -4.675673, -4.565087, -4.45441, 
    -4.343644, -4.232788, -4.121842, -4.010808, -3.899686, -3.788474, 
    -3.677175, -3.565788, -3.454314, -3.342752, -3.231103, -3.119368, 
    -3.007546, -2.895638, -2.783645, -2.671566, -2.559402, -2.447153, 
    -2.334819, -2.222402, -2.1099, -1.997315, -1.884647, -1.771896, 
    -1.659062, -1.546146, -1.433148, -1.320068, -1.206907, -1.093666, 
    -0.9803433, -0.8669407, -0.7534583, -0.6398963, -0.5262551, -0.4125352, 
    -0.2987367, -0.1848601, -0.0709058, 0.04312592, 0.1572347, 0.2714201, 
    0.3856817, 0.5000194, 0.6144325, 0.7289208, 0.8434839, 0.9581214, 
    1.072833, 1.187618, 1.302476, 1.417408, 1.532411, 1.647487, 1.762634, 
    1.877853, 1.993142, 2.108502, 2.223932, 2.339432, 2.455, 2.570638, 
    2.686344, 2.802118, 2.917959, 3.033867, 3.149843, 3.265884, 3.381991, 
    3.498164, 3.614402, 3.730704, 3.84707, 3.9635, 4.079993, 4.196549, 
    4.313167, 4.429847, 4.546588, 4.663391, 4.780253, 4.897176, 5.014159, 
    5.1312, 5.248301, 5.365459, 5.482675, 5.599948, 5.717278, 5.834665, 
    5.952107, 6.069604, 6.187157, 6.304764, 6.422424, 6.540138, 6.657906, 
    6.775725, 6.893596, 7.011519, 7.129493, 7.247517, 7.365591, 7.483715, 
    7.601887, 7.720108, 7.838377, 7.956693, 8.075056, 8.193466, 8.311921, 
    8.430423, 8.548968, 8.667559, 8.786192, 8.90487, 9.02359, 9.142352, 
    9.261156, 9.380001, 9.498887, 9.617813, 9.736779, 9.855784, 9.974828, 
    10.09391, 10.21303, 10.33218, 10.45138, 10.5706, 10.68987, 10.80917, 
    10.9285, 11.04786, 11.16726, 11.2867, 11.40616, 11.52565, 11.64518, 
    11.76474, 11.88432, 12.00394, 12.12358, 12.24326, 12.36296, 12.48269, 
    12.60244, 12.72222, 12.84202, 12.96185, 13.08171, 13.20159, 13.32149, 
    13.44141, 13.56136, 13.68132, 13.80131, 13.92132, 14.04135, 14.16139, 
    14.28146, 14.40154, 14.52164, 14.64176, 14.76189, 14.88204, 15.0022, 
    15.12238, 15.24258, 15.36278, 15.483, 15.60323, 15.72348, 15.84373, 
    15.96399, 16.08427, 16.20455, 16.32484, 16.44514, 16.56545, 16.68576, 
    16.80609, 16.92641, 17.04675, 17.16708, 17.28742, 17.40777, 17.52811, 
    17.64846, 17.76881, 17.88917, 18.00952, 18.12987, 18.25022, 18.37057, 
    18.49092, 18.61127, 18.73161, 18.85195, 18.97229, 19.09262, 19.21295, 
    19.33327, 19.45358, 19.57389, 19.69419, 19.81448, 19.93476, 20.05503, 
    20.17529, 20.29555, 20.41579, 20.53602, 20.65623, 20.77644, 20.89663, 
    21.0168, 21.13697, 21.25711, 21.37724, 21.49736, 21.61746, 21.73754, 
    21.8576, 21.97764, 22.09767, 22.21767, 22.33766, 22.45762, 22.57756, 
    22.69748, 22.81738, 22.93725, 23.0571, 23.17693, 23.29673, 23.41651, 
    23.53625, 23.65598, 23.77567, 23.89534, 24.01498, 24.13459, 24.25418, 
    24.37373, 24.49325, 24.61274, 24.7322, 24.85163, 24.97102, 25.09038, 
    25.20971, 25.329, 25.44826, 25.56748, 25.68667, 25.80582, 25.92493, 
    26.04401, 26.16304, 26.28204, 26.401, 26.51992, 26.6388, 26.75764, 
    26.87644, 26.99519, 27.11391, 27.23258, 27.3512, 27.46979, 27.58833, 
    27.70682, 27.82527, 27.94367, 28.06203, 28.18033, 28.2986, 28.41681, 
    28.53498, 28.65309, 28.77116, 28.88917, 29.00714, 29.12505, 29.24292, 
    29.36073, 29.47849, 29.59619, 29.71384, 29.83144, 29.94899, 30.06647, 
    30.18391, 30.30128, 30.41861, 30.53587, 30.65308, 30.77023, 30.88732, 
    31.00435, 31.12132, 31.23824, 31.35509, 31.47188, 31.58861, 31.70528, 
    31.82189, 31.93844, 32.05492, 32.17134, 32.2877, 32.40399, 32.52022, 
    32.63638, 32.75248, 32.86851, 32.98447, 33.10037, 33.2162, 33.33196, 
    33.44766, 33.56329, 33.67884, 33.79433, 33.90975, 34.0251, 34.14038, 
    34.25558, 34.37072, 34.48579, 34.60078, 34.7157, 34.83054, 34.94532, 
    35.06002, 35.17464, 35.2892, 35.40367, 35.51807, 35.6324, 35.74665, 
    35.86082, 35.97492, 36.08894, 36.20288, 36.31674, 36.43053, 36.54424, 
    36.65786, 36.77142, 36.88488, 36.99828, 37.11158, 37.22481, 37.33796, 
    37.45103, 37.56401, 37.67691, 37.78974, 37.90247, 38.01513, 38.1277,
  -12.23007, -12.12616, -12.02215, -11.91804, -11.81382, -11.7095, -11.60508, 
    -11.50055, -11.39593, -11.2912, -11.18637, -11.08143, -10.9764, 
    -10.87126, -10.76602, -10.66068, -10.55523, -10.44969, -10.34405, 
    -10.2383, -10.13245, -10.0265, -9.920455, -9.814305, -9.708055, 
    -9.601706, -9.495255, -9.388705, -9.282056, -9.175306, -9.068458, 
    -8.96151, -8.854462, -8.747315, -8.640071, -8.532727, -8.425285, 
    -8.317744, -8.210106, -8.10237, -7.994536, -7.886604, -7.778575, 
    -7.67045, -7.562227, -7.453907, -7.345491, -7.236978, -7.12837, 
    -7.019665, -6.910865, -6.801969, -6.692978, -6.583892, -6.474711, 
    -6.365435, -6.256065, -6.146601, -6.037043, -5.927391, -5.817646, 
    -5.707808, -5.597876, -5.487852, -5.377735, -5.267526, -5.157225, 
    -5.046832, -4.936348, -4.825772, -4.715106, -4.604349, -4.493501, 
    -4.382563, -4.271535, -4.160418, -4.049211, -3.937915, -3.826531, 
    -3.715057, -3.603496, -3.491847, -3.38011, -3.268285, -3.156374, 
    -3.044375, -2.932291, -2.82012, -2.707863, -2.595521, -2.483093, 
    -2.370581, -2.257983, -2.145302, -2.032537, -1.919688, -1.806755, 
    -1.69374, -1.580642, -1.467461, -1.354199, -1.240855, -1.127429, 
    -1.013923, -0.9003359, -0.7866685, -0.6729212, -0.5590944, -0.4451883, 
    -0.3312033, -0.2171398, -0.1029981, 0.01122129, 0.1255182, 0.2398921, 
    0.3543427, 0.4688696, 0.5834724, 0.6981508, 0.8129043, 0.9277326, 
    1.042635, 1.157612, 1.272662, 1.387786, 1.502982, 1.618251, 1.733592, 
    1.849005, 1.964488, 2.080043, 2.195668, 2.311363, 2.427127, 2.542961, 
    2.658863, 2.774834, 2.890872, 3.006978, 3.123151, 3.239391, 3.355697, 
    3.472069, 3.588506, 3.705007, 3.821573, 3.938204, 4.054897, 4.171654, 
    4.288474, 4.405355, 4.522298, 4.639303, 4.756369, 4.873495, 4.99068, 
    5.107925, 5.225229, 5.342592, 5.460012, 5.577491, 5.695026, 5.812618, 
    5.930265, 6.047969, 6.165728, 6.283541, 6.401409, 6.51933, 6.637305, 
    6.755332, 6.873411, 6.991542, 7.109725, 7.227958, 7.346241, 7.464574, 
    7.582956, 7.701387, 7.819866, 7.938393, 8.056967, 8.175588, 8.294254, 
    8.412967, 8.531725, 8.650527, 8.769373, 8.888263, 9.007195, 9.126171, 
    9.245189, 9.364247, 9.483347, 9.602487, 9.721666, 9.840886, 9.960144, 
    10.07944, 10.19877, 10.31814, 10.43755, 10.557, 10.67648, 10.79599, 
    10.91554, 11.03512, 11.15474, 11.27438, 11.39406, 11.51378, 11.63352, 
    11.7533, 11.8731, 11.99293, 12.1128, 12.23269, 12.3526, 12.47255, 
    12.59252, 12.71252, 12.83255, 12.95259, 13.07267, 13.19276, 13.31288, 
    13.43303, 13.55319, 13.67338, 13.79359, 13.91381, 14.03406, 14.15433, 
    14.27461, 14.39492, 14.51524, 14.63558, 14.75593, 14.8763, 14.99669, 
    15.11708, 15.2375, 15.35793, 15.47836, 15.59882, 15.71928, 15.83976, 
    15.96024, 16.08074, 16.20124, 16.32176, 16.44228, 16.56281, 16.68334, 
    16.80389, 16.92443, 17.04499, 17.16555, 17.28611, 17.40668, 17.52724, 
    17.64782, 17.76839, 17.88896, 18.00954, 18.13011, 18.25068, 18.37126, 
    18.49183, 18.6124, 18.73296, 18.85353, 18.97408, 19.09464, 19.21518, 
    19.33572, 19.45626, 19.57679, 19.69731, 19.81782, 19.93832, 20.05882, 
    20.1793, 20.29977, 20.42024, 20.54069, 20.66113, 20.78155, 20.90196, 
    21.02236, 21.14274, 21.26311, 21.38346, 21.5038, 21.62411, 21.74442, 
    21.8647, 21.98496, 22.10521, 22.22543, 22.34563, 22.46582, 22.58598, 
    22.70612, 22.82623, 22.94633, 23.0664, 23.18644, 23.30646, 23.42646, 
    23.54642, 23.66637, 23.78628, 23.90617, 24.02602, 24.14585, 24.26565, 
    24.38542, 24.50516, 24.62487, 24.74454, 24.86419, 24.9838, 25.10337, 
    25.22292, 25.34243, 25.4619, 25.58134, 25.70074, 25.82011, 25.93943, 
    26.05872, 26.17797, 26.29719, 26.41636, 26.5355, 26.65459, 26.77364, 
    26.89265, 27.01162, 27.13055, 27.24943, 27.36827, 27.48706, 27.60581, 
    27.72452, 27.84318, 27.96179, 28.08036, 28.19888, 28.31735, 28.43577, 
    28.55415, 28.67247, 28.79075, 28.90897, 29.02715, 29.14527, 29.26334, 
    29.38136, 29.49933, 29.61724, 29.7351, 29.8529, 29.97065, 30.08835, 
    30.20599, 30.32357, 30.4411, 30.55857, 30.67598, 30.79333, 30.91063, 
    31.02786, 31.14504, 31.26215, 31.37921, 31.4962, 31.61314, 31.73001, 
    31.84682, 31.96357, 32.08025, 32.19687, 32.31343, 32.42992, 32.54634, 
    32.6627, 32.779, 32.89523, 33.01139, 33.12749, 33.24352, 33.35947, 
    33.47537, 33.59119, 33.70694, 33.82263, 33.93824, 34.05378, 34.16926, 
    34.28466, 34.39999, 34.51524, 34.63043, 34.74554, 34.86058, 34.97554, 
    35.09044, 35.20525, 35.32, 35.43466, 35.54925, 35.66376, 35.77821, 
    35.89257, 36.00685, 36.12106, 36.23519, 36.34924, 36.46321, 36.57711, 
    36.69092, 36.80465, 36.91831, 37.03188, 37.14538, 37.25879, 37.37212, 
    37.48537, 37.59854, 37.71162, 37.82462, 37.93755, 38.05038, 38.16313,
  -12.2804, -12.17636, -12.07221, -11.96795, -11.8636, -11.75914, -11.65457, 
    -11.54991, -11.44514, -11.34026, -11.23529, -11.13021, -11.02503, 
    -10.91975, -10.81437, -10.70888, -10.60329, -10.4976, -10.39181, 
    -10.28591, -10.17992, -10.07382, -9.967626, -9.861327, -9.754928, 
    -9.648428, -9.541827, -9.435126, -9.328325, -9.221424, -9.114424, 
    -9.007322, -8.900122, -8.792822, -8.685423, -8.577925, -8.470328, 
    -8.362633, -8.254838, -8.146946, -8.038955, -7.930866, -7.82268, 
    -7.714396, -7.606014, -7.497535, -7.38896, -7.280287, -7.171518, 
    -7.062653, -6.953691, -6.844634, -6.735481, -6.626232, -6.516888, 
    -6.407449, -6.297915, -6.188286, -6.078563, -5.968746, -5.858835, 
    -5.748831, -5.638732, -5.528541, -5.418257, -5.30788, -5.197411, 
    -5.086849, -4.976195, -4.86545, -4.754613, -4.643685, -4.532667, 
    -4.421557, -4.310358, -4.199068, -4.087688, -3.976219, -3.864661, 
    -3.753013, -3.641277, -3.529453, -3.41754, -3.30554, -3.193452, 
    -3.081277, -2.969015, -2.856667, -2.744232, -2.631711, -2.519105, 
    -2.406413, -2.293636, -2.180774, -2.067828, -1.954798, -1.841684, 
    -1.728487, -1.615207, -1.501844, -1.388398, -1.274871, -1.161261, 
    -1.04757, -0.9337986, -0.8199461, -0.7060133, -0.5920004, -0.4779079, 
    -0.3637361, -0.2494854, -0.1351562, -0.02074871, 0.09373656, 0.2082993, 
    0.3229391, 0.4376556, 0.5524484, 0.6673172, 0.7822614, 0.8972809, 
    1.012375, 1.127544, 1.242787, 1.358103, 1.473492, 1.588955, 1.704489, 
    1.820096, 1.935774, 2.051524, 2.167344, 2.283234, 2.399195, 2.515225, 
    2.631324, 2.747492, 2.863728, 2.980032, 3.096403, 3.212842, 3.329346, 
    3.445917, 3.562554, 3.679255, 3.796022, 3.912853, 4.029747, 4.146706, 
    4.263727, 4.380811, 4.497956, 4.615163, 4.732432, 4.849761, 4.967151, 
    5.084599, 5.202108, 5.319675, 5.437301, 5.554984, 5.672725, 5.790522, 
    5.908376, 6.026287, 6.144252, 6.262272, 6.380347, 6.498476, 6.616659, 
    6.734894, 6.853182, 6.971522, 7.089913, 7.208355, 7.326849, 7.445391, 
    7.563983, 7.682625, 7.801315, 7.920053, 8.038837, 8.15767, 8.276548, 
    8.395473, 8.514442, 8.633457, 8.752517, 8.871619, 8.990765, 9.109954, 
    9.229185, 9.348457, 9.467771, 9.587126, 9.70652, 9.825953, 9.945427, 
    10.06494, 10.18449, 10.30407, 10.4237, 10.54336, 10.66305, 10.78278, 
    10.90255, 11.02235, 11.14218, 11.26205, 11.38194, 11.50187, 11.62183, 
    11.74183, 11.86185, 11.9819, 12.10198, 12.22209, 12.34223, 12.46239, 
    12.58258, 12.7028, 12.82304, 12.94331, 13.06361, 13.18392, 13.30426, 
    13.42463, 13.54501, 13.66542, 13.78584, 13.90629, 14.02676, 14.14725, 
    14.26775, 14.38828, 14.50882, 14.62938, 14.74995, 14.87055, 14.99115, 
    15.11177, 15.23241, 15.35306, 15.47372, 15.59439, 15.71508, 15.83577, 
    15.95648, 16.0772, 16.19793, 16.31866, 16.43941, 16.56016, 16.68092, 
    16.80168, 16.92245, 17.04323, 17.16401, 17.28479, 17.40558, 17.52637, 
    17.64717, 17.76796, 17.88876, 18.00955, 18.13035, 18.25115, 18.37194, 
    18.49273, 18.61353, 18.73431, 18.8551, 18.97588, 19.09665, 19.21742, 
    19.33819, 19.45894, 19.57969, 19.70044, 19.82117, 19.9419, 20.06261, 
    20.18332, 20.30401, 20.4247, 20.54537, 20.66603, 20.78667, 20.90731, 
    21.02793, 21.14853, 21.26912, 21.38969, 21.51025, 21.63079, 21.75131, 
    21.87181, 21.9923, 22.11276, 22.23321, 22.35363, 22.47404, 22.59442, 
    22.71478, 22.83511, 22.95543, 23.07571, 23.19598, 23.31622, 23.43643, 
    23.55662, 23.67678, 23.79691, 23.91702, 24.03709, 24.15714, 24.27716, 
    24.39714, 24.5171, 24.63702, 24.75692, 24.87678, 24.9966, 25.1164, 
    25.23616, 25.35588, 25.47557, 25.59523, 25.71485, 25.83443, 25.95397, 
    26.07347, 26.19294, 26.31237, 26.43176, 26.55111, 26.67041, 26.78968, 
    26.9089, 27.02809, 27.14722, 27.26632, 27.38537, 27.50438, 27.62334, 
    27.74226, 27.86113, 27.97996, 28.09873, 28.21746, 28.33615, 28.45478, 
    28.57336, 28.6919, 28.81038, 28.92882, 29.0472, 29.16553, 29.28381, 
    29.40204, 29.52021, 29.63833, 29.7564, 29.87441, 29.99237, 30.11027, 
    30.22812, 30.3459, 30.46364, 30.58131, 30.69893, 30.81648, 30.93398, 
    31.05142, 31.1688, 31.28612, 31.40338, 31.52058, 31.63771, 31.75479, 
    31.8718, 31.98875, 32.10563, 32.22245, 32.33921, 32.4559, 32.57253, 
    32.68909, 32.80558, 32.92201, 33.03837, 33.15466, 33.27089, 33.38705, 
    33.50314, 33.61915, 33.7351, 33.85098, 33.96679, 34.08253, 34.1982, 
    34.31379, 34.42931, 34.54477, 34.66014, 34.77545, 34.89068, 35.00584, 
    35.12092, 35.23593, 35.35086, 35.46571, 35.5805, 35.6952, 35.80983, 
    35.92438, 36.03885, 36.15325, 36.26756, 36.3818, 36.49596, 36.61004, 
    36.72404, 36.83796, 36.9518, 37.06556, 37.17924, 37.29284, 37.40635, 
    37.51978, 37.63313, 37.7464, 37.85958, 37.97268, 38.0857, 38.19863,
  -12.33082, -12.22663, -12.12234, -12.01795, -11.91345, -11.80885, 
    -11.70415, -11.59934, -11.49443, -11.38941, -11.2843, -11.17907, 
    -11.07375, -10.96832, -10.86279, -10.75716, -10.65143, -10.54559, 
    -10.43965, -10.33361, -10.22747, -10.12122, -10.01488, -9.90843, 
    -9.801882, -9.695231, -9.588481, -9.481629, -9.374677, -9.267624, 
    -9.16047, -9.053217, -8.945863, -8.838409, -8.730856, -8.623203, 
    -8.515451, -8.4076, -8.29965, -8.191602, -8.083454, -7.975208, -7.866863, 
    -7.758421, -7.649881, -7.541243, -7.432508, -7.323676, -7.214746, 
    -7.10572, -6.996597, -6.887378, -6.778062, -6.668651, -6.559144, 
    -6.449541, -6.339843, -6.23005, -6.120162, -6.010179, -5.900102, 
    -5.789931, -5.679666, -5.569307, -5.458856, -5.34831, -5.237672, 
    -5.126942, -5.016119, -4.905203, -4.794196, -4.683097, -4.571908, 
    -4.460627, -4.349255, -4.237792, -4.12624, -4.014597, -3.902865, 
    -3.791043, -3.679132, -3.567132, -3.455044, -3.342868, -3.230604, 
    -3.118252, -3.005812, -2.893286, -2.780673, -2.667973, -2.555188, 
    -2.442316, -2.32936, -2.216317, -2.103191, -1.989979, -1.876684, 
    -1.763304, -1.649842, -1.536296, -1.422667, -1.308955, -1.195162, 
    -1.081286, -0.9673294, -0.8532915, -0.7391727, -0.6249736, -0.5106944, 
    -0.3963356, -0.2818974, -0.1673802, -0.05278451, 0.06188945, 0.1766413, 
    0.2914706, 0.4063769, 0.52136, 0.6364195, 0.7515548, 0.8667658, 
    0.9820519, 1.097413, 1.212848, 1.328357, 1.44394, 1.559596, 1.675325, 
    1.791126, 1.907, 2.022944, 2.13896, 2.255047, 2.371204, 2.487431, 
    2.603727, 2.720092, 2.836526, 2.953028, 3.069598, 3.186235, 3.302939, 
    3.41971, 3.536546, 3.653449, 3.770416, 3.887448, 4.004544, 4.121704, 
    4.238927, 4.356213, 4.473561, 4.590971, 4.708443, 4.825976, 4.94357, 
    5.061223, 5.178936, 5.296708, 5.414539, 5.532428, 5.650374, 5.768379, 
    5.886439, 6.004556, 6.122729, 6.240956, 6.359239, 6.477576, 6.595967, 
    6.714411, 6.832908, 6.951457, 7.070057, 7.18871, 7.307413, 7.426166, 
    7.544969, 7.663821, 7.782722, 7.901671, 8.020668, 8.139712, 8.258802, 
    8.377939, 8.497122, 8.616349, 8.735621, 8.854938, 8.974298, 9.0937, 
    9.213145, 9.332632, 9.45216, 9.57173, 9.691339, 9.810987, 9.930676, 
    10.0504, 10.17017, 10.28997, 10.40981, 10.52969, 10.6496, 10.76955, 
    10.88953, 11.00955, 11.1296, 11.24968, 11.36979, 11.48994, 11.61012, 
    11.73033, 11.85057, 11.97084, 12.09114, 12.21147, 12.33183, 12.45221, 
    12.57262, 12.69306, 12.81352, 12.93401, 13.05452, 13.17506, 13.29562, 
    13.4162, 13.53681, 13.65744, 13.77808, 13.89875, 14.01944, 14.14015, 
    14.26088, 14.38162, 14.50239, 14.62317, 14.74397, 14.86478, 14.98561, 
    15.10645, 15.22731, 15.34818, 15.46906, 15.58996, 15.71087, 15.83178, 
    15.95271, 16.07365, 16.1946, 16.31556, 16.43653, 16.5575, 16.67848, 
    16.79947, 16.92046, 17.04146, 17.16247, 17.28347, 17.40448, 17.5255, 
    17.64651, 17.76753, 17.88855, 18.00957, 18.13059, 18.25161, 18.37263, 
    18.49364, 18.61466, 18.73567, 18.85668, 18.97768, 19.09868, 19.21967, 
    19.34066, 19.46164, 19.58261, 19.70357, 19.82453, 19.94548, 20.06642, 
    20.18734, 20.30826, 20.42917, 20.55006, 20.67094, 20.79181, 20.91267, 
    21.03351, 21.15433, 21.27514, 21.39594, 21.51672, 21.63748, 21.75822, 
    21.87894, 21.99965, 22.12033, 22.241, 22.36165, 22.48227, 22.60287, 
    22.72345, 22.84401, 22.96454, 23.08505, 23.20553, 23.32599, 23.44643, 
    23.56683, 23.68721, 23.80756, 23.92789, 24.04818, 24.16845, 24.28868, 
    24.40889, 24.52906, 24.64921, 24.76932, 24.8894, 25.00944, 25.12945, 
    25.24943, 25.36937, 25.48928, 25.60915, 25.72898, 25.84878, 25.96854, 
    26.08826, 26.20794, 26.32759, 26.44719, 26.56675, 26.68627, 26.80575, 
    26.92519, 27.04459, 27.16394, 27.28325, 27.40251, 27.52173, 27.64091, 
    27.76004, 27.87912, 27.99816, 28.11715, 28.23609, 28.35498, 28.47383, 
    28.59262, 28.71137, 28.83006, 28.94871, 29.0673, 29.18584, 29.30433, 
    29.42276, 29.54115, 29.65948, 29.77775, 29.89597, 30.01413, 30.13224, 
    30.25029, 30.36829, 30.48622, 30.6041, 30.72193, 30.83969, 30.95739, 
    31.07504, 31.19262, 31.31014, 31.4276, 31.54501, 31.66234, 31.77962, 
    31.89683, 32.01398, 32.13107, 32.24809, 32.36505, 32.48194, 32.59877, 
    32.71553, 32.83222, 32.94884, 33.06541, 33.1819, 33.29832, 33.41467, 
    33.53096, 33.64717, 33.76332, 33.8794, 33.9954, 34.11134, 34.2272, 
    34.34299, 34.4587, 34.57435, 34.68992, 34.80542, 34.92084, 35.03619, 
    35.15146, 35.26666, 35.38179, 35.49683, 35.6118, 35.7267, 35.84151, 
    35.95626, 36.07092, 36.1855, 36.30001, 36.41443, 36.52878, 36.64304, 
    36.75723, 36.87133, 36.98536, 37.0993, 37.21317, 37.32695, 37.44065, 
    37.55426, 37.6678, 37.78125, 37.89461, 38.00789, 38.12109, 38.2342,
  -12.38132, -12.277, -12.17257, -12.06803, -11.9634, -11.85865, -11.75381, 
    -11.64886, -11.5438, -11.43865, -11.33338, -11.22802, -11.12255, 
    -11.01698, -10.91131, -10.80553, -10.69965, -10.59366, -10.48758, 
    -10.38139, -10.2751, -10.16871, -10.06221, -9.955616, -9.848917, 
    -9.742117, -9.635216, -9.528213, -9.421109, -9.313904, -9.206598, 
    -9.099192, -8.991685, -8.884078, -8.77637, -8.668563, -8.560656, 
    -8.452649, -8.344543, -8.236338, -8.128033, -8.019629, -7.911128, 
    -7.802527, -7.693828, -7.585031, -7.476136, -7.367144, -7.258053, 
    -7.148866, -7.039582, -6.930201, -6.820723, -6.711148, -6.601478, 
    -6.491711, -6.381849, -6.271891, -6.161838, -6.05169, -5.941447, 
    -5.831109, -5.720677, -5.610151, -5.499531, -5.388818, -5.278011, 
    -5.167111, -5.056118, -4.945033, -4.833856, -4.722586, -4.611224, 
    -4.499771, -4.388227, -4.276592, -4.164866, -4.05305, -3.941143, 
    -3.829147, -3.717061, -3.604886, -3.492622, -3.38027, -3.267828, 
    -3.155299, -3.042682, -2.929978, -2.817186, -2.704308, -2.591343, 
    -2.478292, -2.365155, -2.251932, -2.138624, -2.025231, -1.911754, 
    -1.798192, -1.684546, -1.570817, -1.457004, -1.343109, -1.229131, 
    -1.115071, -1.000929, -0.8867049, -0.7724001, -0.6580144, -0.5435483, 
    -0.4290021, -0.3143761, -0.1996708, -0.08488651, 0.02997643, 0.1449176, 
    0.2599367, 0.3750333, 0.490207, 0.6054574, 0.7207841, 0.8361868, 
    0.9516651, 1.067219, 1.182847, 1.298549, 1.414326, 1.530176, 1.646099, 
    1.762096, 1.878164, 1.994304, 2.110516, 2.226799, 2.343153, 2.459577, 
    2.576071, 2.692634, 2.809266, 2.925967, 3.042736, 3.159572, 3.276476, 
    3.393446, 3.510483, 3.627586, 3.744754, 3.861987, 3.979285, 4.096647, 
    4.214073, 4.331562, 4.449113, 4.566727, 4.684402, 4.802139, 4.919937, 
    5.037795, 5.155714, 5.273691, 5.391727, 5.509822, 5.627975, 5.746186, 
    5.864453, 5.982778, 6.101158, 6.219594, 6.338084, 6.45663, 6.575229, 
    6.693882, 6.812589, 6.931347, 7.050158, 7.16902, 7.287934, 7.406898, 
    7.525912, 7.644975, 7.764088, 7.883248, 8.002458, 8.121714, 8.241017, 
    8.360367, 8.479762, 8.599203, 8.718689, 8.838219, 8.957792, 9.07741, 
    9.197069, 9.316771, 9.436514, 9.556298, 9.676124, 9.795988, 9.915893, 
    10.03584, 10.15582, 10.27584, 10.39589, 10.51599, 10.63612, 10.75628, 
    10.87648, 10.99671, 11.11698, 11.23728, 11.35762, 11.47798, 11.59838, 
    11.71881, 11.83927, 11.95976, 12.08028, 12.20083, 12.3214, 12.44201, 
    12.56264, 12.6833, 12.80398, 12.92469, 13.04542, 13.16618, 13.28696, 
    13.40776, 13.52859, 13.64944, 13.77031, 13.8912, 14.01211, 14.13304, 
    14.25399, 14.37496, 14.49594, 14.61694, 14.73796, 14.859, 14.98005, 
    15.10111, 15.22219, 15.34329, 15.46439, 15.58551, 15.70664, 15.82778, 
    15.94894, 16.0701, 16.19127, 16.31245, 16.43364, 16.55484, 16.67604, 
    16.79725, 16.91847, 17.03969, 17.16092, 17.28215, 17.40339, 17.52462, 
    17.64586, 17.7671, 17.88835, 18.00959, 18.13083, 18.25208, 18.37332, 
    18.49456, 18.61579, 18.73703, 18.85826, 18.97948, 19.1007, 19.22192, 
    19.34313, 19.46433, 19.58553, 19.70672, 19.8279, 19.94907, 20.07023, 
    20.19138, 20.31252, 20.43365, 20.55477, 20.67587, 20.79696, 20.91804, 
    21.0391, 21.16015, 21.28118, 21.4022, 21.5232, 21.64418, 21.76515, 
    21.88609, 22.00702, 22.12793, 22.24881, 22.36968, 22.49052, 22.61135, 
    22.73215, 22.85293, 22.97368, 23.09441, 23.21511, 23.33579, 23.45645, 
    23.57707, 23.69767, 23.81824, 23.93879, 24.0593, 24.17978, 24.30024, 
    24.42067, 24.54106, 24.66142, 24.78175, 24.90204, 25.02231, 25.14254, 
    25.26273, 25.38289, 25.50301, 25.6231, 25.74315, 25.86316, 25.98314, 
    26.10308, 26.22297, 26.34283, 26.46265, 26.58243, 26.70217, 26.82186, 
    26.94151, 27.06112, 27.18069, 27.30021, 27.41969, 27.53913, 27.65852, 
    27.77786, 27.89715, 28.0164, 28.1356, 28.25476, 28.37386, 28.49292, 
    28.61192, 28.73088, 28.84978, 28.96864, 29.08744, 29.20619, 29.32489, 
    29.44353, 29.56213, 29.68066, 29.79914, 29.91757, 30.03594, 30.15426, 
    30.27252, 30.39072, 30.50886, 30.62695, 30.74498, 30.86294, 30.98085, 
    31.0987, 31.21649, 31.33422, 31.45188, 31.56949, 31.68703, 31.80451, 
    31.92192, 32.03927, 32.15656, 32.27378, 32.39094, 32.50803, 32.62506, 
    32.74202, 32.85891, 32.97574, 33.0925, 33.20919, 33.32581, 33.44236, 
    33.55885, 33.67526, 33.7916, 33.90787, 34.02407, 34.1402, 34.25626, 
    34.37224, 34.48816, 34.60399, 34.71976, 34.83545, 34.95107, 35.06661, 
    35.18207, 35.29746, 35.41278, 35.52802, 35.64318, 35.75826, 35.87327, 
    35.9882, 36.10305, 36.21782, 36.33251, 36.44713, 36.56166, 36.67611, 
    36.79049, 36.90478, 37.01899, 37.13312, 37.24717, 37.36113, 37.47501, 
    37.58881, 37.70253, 37.81616, 37.92971, 38.04317, 38.15655, 38.26985,
  -12.43191, -12.32744, -12.22287, -12.1182, -12.01342, -11.90854, -11.80355, 
    -11.69846, -11.59326, -11.48796, -11.38256, -11.27705, -11.17144, 
    -11.06572, -10.9599, -10.85398, -10.74795, -10.64182, -10.53559, 
    -10.42925, -10.32281, -10.21627, -10.10963, -10.00288, -9.896035, 
    -9.789085, -9.682033, -9.574879, -9.467624, -9.360267, -9.252809, 
    -9.145249, -9.037589, -8.929828, -8.821966, -8.714005, -8.605942, 
    -8.497779, -8.389517, -8.281155, -8.172693, -8.064133, -7.955472, 
    -7.846714, -7.737855, -7.628899, -7.519845, -7.410692, -7.301441, 
    -7.192092, -7.082646, -6.973103, -6.863462, -6.753725, -6.643891, 
    -6.53396, -6.423934, -6.313811, -6.203593, -6.093279, -5.98287, 
    -5.872365, -5.761766, -5.651073, -5.540285, -5.429403, -5.318427, 
    -5.207358, -5.096195, -4.98494, -4.873591, -4.76215, -4.650617, 
    -4.538992, -4.427276, -4.315467, -4.203568, -4.091578, -3.979497, 
    -3.867326, -3.755065, -3.642714, -3.530274, -3.417745, -3.305127, 
    -3.19242, -3.079625, -2.966743, -2.853772, -2.740715, -2.62757, 
    -2.514339, -2.401021, -2.287618, -2.174129, -2.060554, -1.946895, 
    -1.83315, -1.719321, -1.605409, -1.491412, -1.377333, -1.26317, 
    -1.148924, -1.034597, -0.9201871, -0.8056958, -0.6911233, -0.57647, 
    -0.4617361, -0.3469221, -0.2320284, -0.1170552, -0.002002946, 0.1131279, 
    0.2283371, 0.3436241, 0.4589887, 0.5744304, 0.6899489, 0.8055437, 
    0.9212144, 1.036961, 1.152782, 1.268679, 1.384649, 1.500694, 1.616812, 
    1.733003, 1.849267, 1.965603, 2.082012, 2.198491, 2.315042, 2.431664, 
    2.548355, 2.665117, 2.781947, 2.898847, 3.015815, 3.132851, 3.249955, 
    3.367126, 3.484363, 3.601667, 3.719037, 3.836472, 3.953972, 4.071536, 
    4.189165, 4.306857, 4.424612, 4.542429, 4.660309, 4.77825, 4.896253, 
    5.014316, 5.13244, 5.250623, 5.368865, 5.487167, 5.605527, 5.723944, 
    5.842419, 5.960951, 6.079539, 6.198183, 6.316883, 6.435637, 6.554446, 
    6.673308, 6.792224, 6.911193, 7.030214, 7.149287, 7.268411, 7.387586, 
    7.506812, 7.626087, 7.745411, 7.864785, 7.984206, 8.103675, 8.223191, 
    8.342754, 8.462363, 8.582018, 8.701718, 8.821463, 8.941251, 9.061082, 
    9.180957, 9.300874, 9.420833, 9.540833, 9.660873, 9.780954, 9.901075, 
    10.02123, 10.14143, 10.26167, 10.38194, 10.50225, 10.6226, 10.74298, 
    10.8634, 10.98385, 11.10434, 11.22486, 11.34541, 11.466, 11.58662, 
    11.70726, 11.82794, 11.94865, 12.06939, 12.19016, 12.31096, 12.43178, 
    12.55263, 12.67351, 12.79441, 12.91534, 13.0363, 13.15727, 13.27828, 
    13.3993, 13.52035, 13.64142, 13.76251, 13.88362, 14.00476, 14.12591, 
    14.24708, 14.36827, 14.48948, 14.6107, 14.73195, 14.8532, 14.97448, 
    15.09576, 15.21707, 15.33838, 15.45971, 15.58105, 15.70241, 15.82377, 
    15.94515, 16.06654, 16.18793, 16.30934, 16.43075, 16.55217, 16.6736, 
    16.79503, 16.91647, 17.03792, 17.15937, 17.28082, 17.40228, 17.52374, 
    17.64521, 17.76667, 17.88814, 18.00961, 18.13107, 18.25254, 18.37401, 
    18.49547, 18.61693, 18.73839, 18.85984, 18.98129, 19.10274, 19.22418, 
    19.34561, 19.46704, 19.58846, 19.70987, 19.83127, 19.95267, 20.07405, 
    20.19543, 20.31679, 20.43814, 20.55948, 20.68081, 20.80212, 20.92342, 
    21.04471, 21.16598, 21.28724, 21.40847, 21.5297, 21.6509, 21.77209, 
    21.89326, 22.01441, 22.13553, 22.25664, 22.37773, 22.4988, 22.61984, 
    22.74087, 22.86186, 22.98284, 23.10379, 23.22471, 23.34562, 23.46649, 
    23.58734, 23.70815, 23.82895, 23.94971, 24.07044, 24.19115, 24.31182, 
    24.43247, 24.55308, 24.67366, 24.79421, 24.91472, 25.0352, 25.15565, 
    25.27606, 25.39644, 25.51678, 25.63708, 25.75735, 25.87758, 25.99778, 
    26.11793, 26.23804, 26.35812, 26.47815, 26.59815, 26.7181, 26.83801, 
    26.95788, 27.0777, 27.19748, 27.31722, 27.43691, 27.55656, 27.67616, 
    27.79572, 27.91523, 28.03469, 28.1541, 28.27347, 28.39278, 28.51205, 
    28.63127, 28.75044, 28.86955, 28.98862, 29.10763, 29.22659, 29.3455, 
    29.46435, 29.58315, 29.7019, 29.82059, 29.93922, 30.0578, 30.17632, 
    30.29479, 30.4132, 30.53155, 30.64984, 30.76808, 30.88625, 31.00436, 
    31.12242, 31.24041, 31.35834, 31.47621, 31.59402, 31.71177, 31.82945, 
    31.94707, 32.06462, 32.18211, 32.29953, 32.41689, 32.53419, 32.65141, 
    32.76857, 32.88567, 33.00269, 33.11965, 33.23654, 33.35336, 33.47011, 
    33.58679, 33.7034, 33.81994, 33.93641, 34.0528, 34.16913, 34.28538, 
    34.40156, 34.51767, 34.6337, 34.74966, 34.86554, 34.98135, 35.09709, 
    35.21275, 35.32833, 35.44384, 35.55927, 35.67462, 35.78989, 35.90509, 
    36.02021, 36.13525, 36.25021, 36.36509, 36.47989, 36.59461, 36.70925, 
    36.82381, 36.93829, 37.05269, 37.167, 37.28123, 37.39538, 37.50945, 
    37.62343, 37.73733, 37.85115, 37.96488, 38.07853, 38.19209, 38.30556,
  -12.48257, -12.37797, -12.27326, -12.16845, -12.06353, -11.9585, -11.85338, 
    -11.74814, -11.6428, -11.53736, -11.43181, -11.32616, -11.2204, 
    -11.11454, -11.00858, -10.90251, -10.79634, -10.69006, -10.58368, 
    -10.4772, -10.37061, -10.26392, -10.15713, -10.05023, -9.943235, 
    -9.836136, -9.728932, -9.621628, -9.51422, -9.406712, -9.299101, 
    -9.191388, -9.083575, -8.97566, -8.867644, -8.759527, -8.651309, 
    -8.542991, -8.434572, -8.326054, -8.217435, -8.108717, -7.999898, 
    -7.890981, -7.781964, -7.672848, -7.563633, -7.45432, -7.344909, 
    -7.235399, -7.125791, -7.016085, -6.906282, -6.796381, -6.686384, 
    -6.576289, -6.466098, -6.355811, -6.245427, -6.134947, -6.024371, 
    -5.9137, -5.802934, -5.692072, -5.581116, -5.470066, -5.358921, 
    -5.247682, -5.13635, -5.024923, -4.913404, -4.801792, -4.690087, 
    -4.57829, -4.4664, -4.354419, -4.242346, -4.130182, -4.017926, -3.90558, 
    -3.793144, -3.680617, -3.568001, -3.455295, -3.342499, -3.229615, 
    -3.116642, -3.003581, -2.890432, -2.777195, -2.663871, -2.550459, 
    -2.436961, -2.323376, -2.209705, -2.095949, -1.982107, -1.86818, 
    -1.754168, -1.640071, -1.525891, -1.411626, -1.297279, -1.182848, 
    -1.068334, -0.9537382, -0.8390603, -0.7243007, -0.6094599, -0.4945381, 
    -0.3795358, -0.2644532, -0.1492909, -0.03404909, 0.08127177, 0.1966713, 
    0.3121492, 0.4277049, 0.5433382, 0.6590487, 0.7748358, 0.8906994, 
    1.006639, 1.122654, 1.238744, 1.354909, 1.471148, 1.587462, 1.703849, 
    1.820309, 1.936841, 2.053446, 2.170123, 2.286871, 2.40369, 2.52058, 
    2.63754, 2.75457, 2.871668, 2.988836, 3.106072, 3.223376, 3.340748, 
    3.458187, 3.575692, 3.693263, 3.8109, 3.928603, 4.04637, 4.164202, 
    4.282097, 4.400056, 4.518078, 4.636162, 4.754308, 4.872516, 4.990785, 
    5.109115, 5.227504, 5.345953, 5.464461, 5.583028, 5.701653, 5.820336, 
    5.939076, 6.057872, 6.176725, 6.295633, 6.414597, 6.533615, 6.652688, 
    6.771814, 6.890993, 7.010225, 7.129509, 7.248845, 7.368231, 7.487669, 
    7.607156, 7.726693, 7.846279, 7.965913, 8.085595, 8.205325, 8.325102, 
    8.444925, 8.564795, 8.684709, 8.804667, 8.924671, 9.044718, 9.164807, 
    9.284941, 9.405115, 9.525331, 9.645589, 9.765886, 9.886224, 10.0066, 
    10.12702, 10.24747, 10.36796, 10.48849, 10.60905, 10.72966, 10.85029, 
    10.97096, 11.09167, 11.21241, 11.33318, 11.45399, 11.57482, 11.69569, 
    11.81659, 11.93752, 12.05848, 12.17947, 12.30048, 12.42153, 12.5426, 
    12.6637, 12.78482, 12.90597, 13.02715, 13.14835, 13.26958, 13.39082, 
    13.51209, 13.63338, 13.7547, 13.87603, 13.99739, 14.11876, 14.24016, 
    14.36157, 14.483, 14.60445, 14.72591, 14.84739, 14.96889, 15.0904, 
    15.21193, 15.33347, 15.45502, 15.57659, 15.69817, 15.81976, 15.94135, 
    16.06297, 16.18459, 16.30621, 16.42785, 16.5495, 16.67115, 16.79281, 
    16.91447, 17.03614, 17.15782, 17.2795, 17.40118, 17.52287, 17.64455, 
    17.76624, 17.88793, 18.00962, 18.13132, 18.25301, 18.3747, 18.49638, 
    18.61807, 18.73975, 18.86143, 18.9831, 19.10477, 19.22644, 19.34809, 
    19.46975, 19.59139, 19.71303, 19.83465, 19.95627, 20.07788, 20.19948, 
    20.32107, 20.44264, 20.56421, 20.68576, 20.80729, 20.92882, 21.05033, 
    21.17182, 21.2933, 21.41476, 21.53621, 21.65764, 21.77905, 21.90044, 
    22.02181, 22.14316, 22.26449, 22.3858, 22.50709, 22.62836, 22.7496, 
    22.87082, 22.99202, 23.11319, 23.23434, 23.35546, 23.47655, 23.59762, 
    23.71866, 23.83967, 23.96066, 24.08161, 24.20254, 24.32343, 24.44429, 
    24.56513, 24.68593, 24.80669, 24.92743, 25.04813, 25.16879, 25.28942, 
    25.41002, 25.53058, 25.6511, 25.77159, 25.89203, 26.01244, 26.13281, 
    26.25315, 26.37344, 26.49369, 26.6139, 26.73407, 26.85419, 26.97428, 
    27.09431, 27.21431, 27.33426, 27.45417, 27.57403, 27.69385, 27.81362, 
    27.93334, 28.05301, 28.17264, 28.29222, 28.41175, 28.53123, 28.65066, 
    28.77004, 28.88936, 29.00864, 29.12786, 29.24703, 29.36615, 29.48522, 
    29.60423, 29.72318, 29.84208, 29.96092, 30.07971, 30.19844, 30.31712, 
    30.43573, 30.55429, 30.67279, 30.79123, 30.90961, 31.02793, 31.14619, 
    31.26439, 31.38252, 31.5006, 31.61861, 31.73656, 31.85444, 31.97226, 
    32.09002, 32.20771, 32.32534, 32.4429, 32.56039, 32.67782, 32.79519, 
    32.91248, 33.0297, 33.14686, 33.26395, 33.38097, 33.49791, 33.61479, 
    33.7316, 33.84834, 33.965, 34.0816, 34.19812, 34.31457, 34.43094, 
    34.54725, 34.66347, 34.77962, 34.8957, 35.01171, 35.12763, 35.24348, 
    35.35926, 35.47496, 35.59058, 35.70612, 35.82159, 35.93698, 36.05228, 
    36.16751, 36.28266, 36.39773, 36.51272, 36.62763, 36.74246, 36.8572, 
    36.97187, 37.08645, 37.20095, 37.31537, 37.42971, 37.54396, 37.65813, 
    37.77221, 37.88621, 38.00012, 38.11395, 38.22769, 38.34135,
  -12.53333, -12.42858, -12.32374, -12.21878, -12.11372, -12.00856, 
    -11.90329, -11.79791, -11.69243, -11.58684, -11.48115, -11.37535, 
    -11.26945, -11.16345, -11.05734, -10.95112, -10.84481, -10.73838, 
    -10.63186, -10.52523, -10.41849, -10.31165, -10.20471, -10.09767, 
    -9.99052, -9.883269, -9.775916, -9.66846, -9.560901, -9.453239, 
    -9.345476, -9.237611, -9.129643, -9.021575, -8.913404, -8.805132, 
    -8.696759, -8.588285, -8.479711, -8.371035, -8.262259, -8.153382, 
    -8.044406, -7.93533, -7.826154, -7.716878, -7.607504, -7.49803, 
    -7.388457, -7.278786, -7.169016, -7.059148, -6.949183, -6.839118, 
    -6.728957, -6.618698, -6.508342, -6.39789, -6.28734, -6.176694, 
    -6.065952, -5.955114, -5.84418, -5.733151, -5.622026, -5.510807, 
    -5.399493, -5.288085, -5.176582, -5.064985, -4.953295, -4.841511, 
    -4.729634, -4.617664, -4.505601, -4.393447, -4.2812, -4.168861, 
    -4.056432, -3.94391, -3.831298, -3.718596, -3.605803, -3.49292, 
    -3.379947, -3.266885, -3.153734, -3.040494, -2.927165, -2.813749, 
    -2.700244, -2.586652, -2.472973, -2.359207, -2.245354, -2.131416, 
    -2.017391, -1.90328, -1.789085, -1.674805, -1.56044, -1.44599, -1.331457, 
    -1.216841, -1.102141, -0.9873589, -0.872494, -0.757547, -0.6425184, 
    -0.5274084, -0.4122174, -0.2969459, -0.1815941, -0.06616242, 0.04934871, 
    0.1649389, 0.2806079, 0.3963551, 0.5121803, 0.6280831, 0.744063, 
    0.8601196, 0.9762527, 1.092462, 1.208746, 1.325106, 1.44154, 1.558049, 
    1.674632, 1.791288, 1.908017, 2.024819, 2.141693, 2.258639, 2.375656, 
    2.492745, 2.609903, 2.727132, 2.844431, 2.961799, 3.079235, 3.19674, 
    3.314313, 3.431953, 3.54966, 3.667434, 3.785273, 3.903178, 4.021149, 
    4.139184, 4.257284, 4.375447, 4.493673, 4.611962, 4.730314, 4.848727, 
    4.967202, 5.085738, 5.204334, 5.322989, 5.441705, 5.56048, 5.679313, 
    5.798203, 5.917152, 6.036157, 6.155219, 6.274337, 6.39351, 6.512738, 
    6.632021, 6.751358, 6.870748, 6.990191, 7.109686, 7.229234, 7.348833, 
    7.468482, 7.588182, 7.707932, 7.827731, 7.947579, 8.067475, 8.187419, 
    8.307409, 8.427447, 8.547531, 8.66766, 8.787834, 8.908053, 9.028316, 
    9.148622, 9.26897, 9.389361, 9.509794, 9.630269, 9.750784, 9.871338, 
    9.991933, 10.11257, 10.23324, 10.35395, 10.47469, 10.59548, 10.7163, 
    10.83715, 10.95804, 11.07897, 11.19993, 11.32092, 11.44194, 11.563, 
    11.68409, 11.80521, 11.92636, 12.04754, 12.16875, 12.28999, 12.41125, 
    12.53255, 12.65387, 12.77521, 12.89659, 13.01798, 13.13941, 13.26085, 
    13.38232, 13.50382, 13.62533, 13.74687, 13.86842, 13.99, 14.1116, 
    14.23322, 14.35485, 14.47651, 14.59818, 14.71987, 14.84157, 14.96329, 
    15.08503, 15.20678, 15.32854, 15.45032, 15.57211, 15.69391, 15.81573, 
    15.93755, 16.05939, 16.18123, 16.30308, 16.42495, 16.54682, 16.66869, 
    16.79058, 16.91247, 17.03436, 17.15626, 17.27816, 17.40007, 17.52198, 
    17.6439, 17.76581, 17.88773, 18.00964, 18.13156, 18.25348, 18.37539, 
    18.4973, 18.61921, 18.74112, 18.86302, 18.98492, 19.10682, 19.2287, 
    19.35059, 19.47246, 19.59433, 19.71619, 19.83805, 19.95989, 20.08172, 
    20.20354, 20.32536, 20.44715, 20.56894, 20.69072, 20.81248, 20.93423, 
    21.05596, 21.17768, 21.29938, 21.42107, 21.54274, 21.66439, 21.78602, 
    21.90763, 22.02923, 22.1508, 22.27236, 22.39389, 22.5154, 22.63689, 
    22.75836, 22.8798, 23.00122, 23.12262, 23.24398, 23.36533, 23.48664, 
    23.60793, 23.72919, 23.85043, 23.97163, 24.09281, 24.21395, 24.33507, 
    24.45615, 24.5772, 24.69822, 24.81921, 24.94016, 25.06108, 25.18197, 
    25.30282, 25.42363, 25.54441, 25.66515, 25.78585, 25.90652, 26.02715, 
    26.14773, 26.26828, 26.38879, 26.50926, 26.62968, 26.75007, 26.87041, 
    26.99071, 27.11097, 27.23118, 27.35135, 27.47147, 27.59154, 27.71157, 
    27.83156, 27.95149, 28.07138, 28.19122, 28.31101, 28.43076, 28.55045, 
    28.67009, 28.78968, 28.90922, 29.02871, 29.14814, 29.26752, 29.38685, 
    29.50612, 29.62535, 29.74451, 29.86362, 29.98267, 30.10167, 30.22061, 
    30.33949, 30.45831, 30.57708, 30.69578, 30.81443, 30.93302, 31.05154, 
    31.17001, 31.28841, 31.40675, 31.52503, 31.64325, 31.7614, 31.87949, 
    31.99752, 32.11548, 32.23337, 32.3512, 32.46896, 32.58666, 32.70429, 
    32.82185, 32.93935, 33.05677, 33.17413, 33.29142, 33.40863, 33.52578, 
    33.64286, 33.75986, 33.8768, 33.99366, 34.11045, 34.22717, 34.34381, 
    34.46038, 34.57688, 34.69331, 34.80965, 34.92593, 35.04212, 35.15825, 
    35.27429, 35.39025, 35.50615, 35.62196, 35.73769, 35.85335, 35.96893, 
    36.08443, 36.19985, 36.31519, 36.43044, 36.54562, 36.66072, 36.77573, 
    36.89067, 37.00552, 37.12029, 37.23498, 37.34958, 37.4641, 37.57854, 
    37.69289, 37.80716, 37.92134, 38.03543, 38.14944, 38.26337, 38.37721,
  -12.58416, -12.47928, -12.37429, -12.2692, -12.164, -12.05869, -11.95328, 
    -11.84776, -11.74214, -11.63641, -11.53057, -11.42463, -11.31859, 
    -11.21244, -11.10618, -10.99982, -10.89336, -10.78679, -10.68012, 
    -10.57334, -10.46646, -10.35947, -10.25238, -10.14519, -10.03789, 
    -9.930487, -9.822983, -9.715375, -9.607664, -9.499851, -9.391935, 
    -9.283916, -9.175796, -9.067573, -8.959248, -8.850821, -8.742292, 
    -8.633662, -8.524931, -8.416099, -8.307165, -8.198131, -8.088996, 
    -7.979761, -7.870426, -7.760991, -7.651456, -7.541821, -7.432088, 
    -7.322255, -7.212323, -7.102293, -6.992164, -6.881936, -6.771611, 
    -6.661188, -6.550667, -6.440049, -6.329334, -6.218522, -6.107613, 
    -5.996608, -5.885506, -5.774309, -5.663016, -5.551628, -5.440144, 
    -5.328566, -5.216892, -5.105124, -4.993263, -4.881308, -4.769258, 
    -4.657116, -4.54488, -4.432552, -4.320131, -4.207618, -4.095013, 
    -3.982317, -3.869529, -3.75665, -3.64368, -3.53062, -3.41747, -3.304229, 
    -3.1909, -3.077481, -2.963973, -2.850377, -2.736692, -2.622919, 
    -2.509059, -2.395111, -2.281076, -2.166955, -2.052747, -1.938454, 
    -1.824074, -1.70961, -1.59506, -1.480426, -1.365707, -1.250905, 
    -1.136019, -1.021049, -0.9059973, -0.7908627, -0.675646, -0.5603476, 
    -0.4449677, -0.3295068, -0.2139652, -0.09834338, 0.01735833, 0.1331395, 
    0.2489999, 0.3649389, 0.4809563, 0.5970517, 0.7132246, 0.8294747, 
    0.9458016, 1.062205, 1.178684, 1.295239, 1.411868, 1.528573, 1.645352, 
    1.762205, 1.879131, 1.99613, 2.113202, 2.230346, 2.347562, 2.464849, 
    2.582207, 2.699636, 2.817134, 2.934702, 3.052339, 3.170045, 3.287819, 
    3.405661, 3.523571, 3.641547, 3.759589, 3.877698, 3.995872, 4.114111, 
    4.232415, 4.350782, 4.469214, 4.587708, 4.706266, 4.824885, 4.943566, 
    5.062309, 5.181112, 5.299975, 5.418898, 5.53788, 5.656922, 5.776021, 
    5.895178, 6.014393, 6.133665, 6.252992, 6.372375, 6.491814, 6.611308, 
    6.730855, 6.850457, 6.970111, 7.089819, 7.209579, 7.32939, 7.449252, 
    7.569165, 7.689128, 7.809141, 7.929203, 8.049313, 8.169471, 8.289677, 
    8.409929, 8.530228, 8.650573, 8.770963, 8.891397, 9.011876, 9.132399, 
    9.252964, 9.373572, 9.494222, 9.614914, 9.735646, 9.856419, 9.977231, 
    10.09808, 10.21897, 10.3399, 10.46087, 10.58187, 10.70291, 10.82398, 
    10.94509, 11.06624, 11.18742, 11.30863, 11.42987, 11.55115, 11.67246, 
    11.7938, 11.91517, 12.03657, 12.158, 12.27946, 12.40095, 12.52247, 
    12.64401, 12.76558, 12.88717, 13.00879, 13.13044, 13.25211, 13.3738, 
    13.49552, 13.61726, 13.73902, 13.8608, 13.9826, 14.10442, 14.22626, 
    14.34812, 14.47, 14.5919, 14.71381, 14.83574, 14.95768, 15.07964, 
    15.20162, 15.32361, 15.44561, 15.56762, 15.68965, 15.81169, 15.93374, 
    16.0558, 16.17787, 16.29995, 16.42203, 16.54413, 16.66623, 16.78834, 
    16.91045, 17.03257, 17.1547, 17.27683, 17.39896, 17.5211, 17.64324, 
    17.76538, 17.88752, 18.00966, 18.1318, 18.25394, 18.37608, 18.49822, 
    18.62036, 18.74249, 18.86462, 18.98674, 19.10886, 19.23098, 19.35308, 
    19.47519, 19.59728, 19.71937, 19.84144, 19.96351, 20.08557, 20.20762, 
    20.32965, 20.45168, 20.57369, 20.69569, 20.81768, 20.93965, 21.06161, 
    21.18355, 21.30548, 21.42739, 21.54928, 21.67115, 21.79301, 21.91485, 
    22.03667, 22.15847, 22.28024, 22.402, 22.52374, 22.64545, 22.76714, 
    22.8888, 23.01044, 23.13206, 23.25365, 23.37522, 23.49676, 23.61827, 
    23.73975, 23.86121, 23.98263, 24.10403, 24.2254, 24.34673, 24.46803, 
    24.58931, 24.71055, 24.83175, 24.95293, 25.07407, 25.19517, 25.31624, 
    25.43727, 25.55827, 25.67923, 25.80015, 25.92104, 26.04188, 26.16269, 
    26.28345, 26.40418, 26.52487, 26.64551, 26.76611, 26.88667, 27.00718, 
    27.12766, 27.24809, 27.36847, 27.4888, 27.6091, 27.72934, 27.84954, 
    27.96969, 28.08979, 28.20985, 28.32985, 28.44981, 28.56971, 28.68957, 
    28.80937, 28.92912, 29.04882, 29.16847, 29.28806, 29.4076, 29.52708, 
    29.64651, 29.76589, 29.88521, 30.00447, 30.12367, 30.24282, 30.36191, 
    30.48094, 30.59992, 30.71883, 30.83768, 30.95648, 31.07521, 31.19388, 
    31.31249, 31.43104, 31.54952, 31.66795, 31.7863, 31.9046, 32.02283, 
    32.14099, 32.25909, 32.37712, 32.49509, 32.61298, 32.73082, 32.84858, 
    32.96627, 33.0839, 33.20146, 33.31894, 33.43636, 33.55371, 33.67099, 
    33.78819, 33.90532, 34.02238, 34.13937, 34.25628, 34.37313, 34.48989, 
    34.60659, 34.7232, 34.83974, 34.95621, 35.07261, 35.18892, 35.30516, 
    35.42132, 35.5374, 35.6534, 35.76933, 35.88518, 36.00095, 36.11664, 
    36.23225, 36.34777, 36.46323, 36.57859, 36.69388, 36.80908, 36.9242, 
    37.03924, 37.1542, 37.26907, 37.38386, 37.49857, 37.61319, 37.72772, 
    37.84217, 37.95654, 38.07082, 38.18501, 38.29912, 38.41314,
  -12.63509, -12.53006, -12.42494, -12.3197, -12.21436, -12.10891, -12.00336, 
    -11.8977, -11.79193, -11.68606, -11.58008, -11.474, -11.36781, -11.26152, 
    -11.15512, -11.04861, -10.942, -10.83528, -10.72846, -10.62154, 
    -10.51451, -10.40737, -10.30013, -10.19279, -10.08534, -9.977789, 
    -9.870133, -9.762375, -9.654512, -9.546546, -9.438478, -9.330306, 
    -9.222032, -9.113654, -9.005175, -8.896592, -8.787909, -8.679122, 
    -8.570234, -8.461245, -8.352154, -8.242962, -8.133669, -8.024275, 
    -7.91478, -7.805185, -7.69549, -7.585695, -7.4758, -7.365806, -7.255712, 
    -7.145518, -7.035226, -6.924835, -6.814346, -6.703758, -6.593072, 
    -6.482289, -6.371408, -6.260429, -6.149354, -6.038181, -5.926912, 
    -5.815547, -5.704085, -5.592527, -5.480874, -5.369125, -5.257282, 
    -5.145343, -5.03331, -4.921183, -4.808961, -4.696646, -4.584237, 
    -4.471735, -4.359139, -4.246452, -4.133672, -4.0208, -3.907836, -3.79478, 
    -3.681634, -3.568396, -3.455068, -3.34165, -3.228141, -3.114543, 
    -3.000855, -2.887079, -2.773214, -2.65926, -2.545218, -2.431088, 
    -2.316871, -2.202567, -2.088176, -1.973699, -1.859136, -1.744487, 
    -1.629752, -1.514932, -1.400028, -1.285039, -1.169967, -1.05481, 
    -0.9395708, -0.8242483, -0.7088432, -0.5933559, -0.4777868, -0.3621363, 
    -0.2464047, -0.1305924, -0.01469981, 0.1012727, 0.2173247, 0.3334559, 
    0.4496658, 0.5659541, 0.6823204, 0.7987642, 0.9152852, 1.031883, 
    1.148557, 1.265307, 1.382133, 1.499033, 1.616009, 1.733058, 1.850182, 
    1.967379, 2.084649, 2.201991, 2.319406, 2.436892, 2.55445, 2.672079, 
    2.789778, 2.907546, 3.025385, 3.143292, 3.261268, 3.379312, 3.497424, 
    3.615603, 3.733849, 3.852161, 3.970539, 4.088983, 4.207491, 4.326064, 
    4.444701, 4.563401, 4.682164, 4.80099, 4.919878, 5.038827, 5.157837, 
    5.276909, 5.39604, 5.515231, 5.63448, 5.753789, 5.873156, 5.99258, 
    6.112061, 6.231599, 6.351193, 6.470843, 6.590547, 6.710307, 6.83012, 
    6.949986, 7.069906, 7.189878, 7.309903, 7.429978, 7.550105, 7.670282, 
    7.790508, 7.910785, 8.031109, 8.151483, 8.271903, 8.392371, 8.512885, 
    8.633446, 8.754052, 8.874703, 8.995399, 9.116138, 9.23692, 9.357746, 
    9.478614, 9.599523, 9.720473, 9.841464, 9.962495, 10.08357, 10.20467, 
    10.32582, 10.44701, 10.56823, 10.68949, 10.81078, 10.93211, 11.05348, 
    11.17488, 11.29631, 11.41778, 11.53928, 11.66081, 11.78237, 11.90396, 
    12.02558, 12.14724, 12.26892, 12.39063, 12.51237, 12.63413, 12.75592, 
    12.87774, 12.99959, 13.12145, 13.24335, 13.36526, 13.4872, 13.60916, 
    13.73115, 13.85315, 13.97518, 14.09723, 14.21929, 14.34138, 14.46348, 
    14.5856, 14.70774, 14.82989, 14.95206, 15.07424, 15.19644, 15.31866, 
    15.44089, 15.56313, 15.68538, 15.80764, 15.92992, 16.0522, 16.1745, 
    16.2968, 16.41911, 16.54144, 16.66376, 16.7861, 16.90844, 17.03078, 
    17.15314, 17.27549, 17.39785, 17.52021, 17.64258, 17.76494, 17.88731, 
    18.00968, 18.13205, 18.25441, 18.37678, 18.49914, 18.62151, 18.74386, 
    18.86622, 18.98857, 19.11091, 19.23326, 19.35559, 19.47791, 19.60023, 
    19.72255, 19.84485, 19.96714, 20.08943, 20.2117, 20.33396, 20.45621, 
    20.57845, 20.70068, 20.82289, 20.94508, 21.06727, 21.18943, 21.31159, 
    21.43372, 21.55584, 21.67794, 21.80002, 21.92208, 22.04412, 22.16615, 
    22.28815, 22.41013, 22.53209, 22.65402, 22.77594, 22.89783, 23.01969, 
    23.14153, 23.26334, 23.38513, 23.50689, 23.62863, 23.75033, 23.87201, 
    23.99366, 24.11527, 24.23686, 24.35842, 24.47995, 24.60144, 24.7229, 
    24.84433, 24.96572, 25.08708, 25.20841, 25.32969, 25.45095, 25.57216, 
    25.69334, 25.81449, 25.93559, 26.05665, 26.17768, 26.29866, 26.41961, 
    26.54051, 26.66137, 26.78219, 26.90296, 27.0237, 27.14438, 27.26503, 
    27.38563, 27.50618, 27.62669, 27.74715, 27.86756, 27.98793, 28.10824, 
    28.22851, 28.34873, 28.4689, 28.58902, 28.70909, 28.8291, 28.94907, 
    29.06898, 29.18884, 29.30864, 29.42839, 29.54809, 29.66773, 29.78731, 
    29.90684, 30.02632, 30.14573, 30.26509, 30.38439, 30.50363, 30.62281, 
    30.74193, 30.86099, 30.97999, 31.09893, 31.21781, 31.33663, 31.45538, 
    31.57407, 31.6927, 31.81126, 31.92976, 32.04819, 32.16656, 32.28486, 
    32.4031, 32.52126, 32.63937, 32.7574, 32.87536, 32.99326, 33.11109, 
    33.22884, 33.34653, 33.46415, 33.5817, 33.69917, 33.81657, 33.93391, 
    34.05117, 34.16835, 34.28546, 34.4025, 34.51946, 34.63635, 34.75317, 
    34.8699, 34.98656, 35.10315, 35.21966, 35.33609, 35.45245, 35.56872, 
    35.68492, 35.80104, 35.91708, 36.03304, 36.14892, 36.26472, 36.38044, 
    36.49607, 36.61163, 36.7271, 36.84249, 36.95781, 37.07303, 37.18818, 
    37.30323, 37.41821, 37.5331, 37.64791, 37.76263, 37.87726, 37.99181, 
    38.10628, 38.22065, 38.33495, 38.44915,
  -12.68609, -12.58093, -12.47567, -12.37029, -12.26481, -12.15922, 
    -12.05353, -11.94772, -11.84181, -11.7358, -11.62968, -11.52345, 
    -11.41712, -11.31068, -11.20413, -11.09748, -10.99072, -10.88386, 
    -10.77689, -10.66982, -10.56264, -10.45536, -10.34797, -10.24047, 
    -10.13288, -10.02518, -9.917369, -9.809459, -9.701445, -9.593327, 
    -9.485105, -9.37678, -9.268352, -9.15982, -9.051186, -8.942448, 
    -8.833608, -8.724666, -8.615622, -8.506474, -8.397226, -8.287876, 
    -8.178425, -8.068871, -7.959218, -7.849463, -7.739607, -7.629651, 
    -7.519595, -7.409439, -7.299182, -7.188826, -7.078371, -6.967816, 
    -6.857163, -6.74641, -6.63556, -6.524611, -6.413563, -6.302418, 
    -6.191175, -6.079835, -5.968399, -5.856864, -5.745234, -5.633507, 
    -5.521684, -5.409765, -5.29775, -5.185641, -5.073436, -4.961136, 
    -4.848742, -4.736254, -4.623672, -4.510995, -4.398226, -4.285363, 
    -4.172408, -4.05936, -3.94622, -3.832988, -3.719664, -3.606249, 
    -3.492742, -3.379145, -3.265458, -3.15168, -3.037813, -2.923856, 
    -2.80981, -2.695675, -2.581452, -2.46714, -2.35274, -2.238253, -2.123679, 
    -2.009018, -1.89427, -1.779436, -1.664516, -1.549511, -1.434421, 
    -1.319245, -1.203986, -1.088642, -0.9732147, -0.857704, -0.7421103, 
    -0.6264339, -0.5106753, -0.3948349, -0.2789129, -0.1629099, -0.04682613, 
    0.06933797, 0.185582, 0.3019056, 0.4183084, 0.53479, 0.6513498, 
    0.7679878, 0.8847032, 1.001496, 1.118365, 1.235311, 1.352333, 1.46943, 
    1.586602, 1.703849, 1.82117, 1.938565, 2.056033, 2.173575, 2.291189, 
    2.408875, 2.526632, 2.644461, 2.762361, 2.880331, 2.99837, 3.11648, 
    3.234658, 3.352905, 3.47122, 3.589602, 3.708051, 3.826568, 3.94515, 
    4.063798, 4.182511, 4.30129, 4.420132, 4.539039, 4.658009, 4.777041, 
    4.896136, 5.015293, 5.134511, 5.25379, 5.37313, 5.492529, 5.611989, 
    5.731506, 5.851083, 5.970717, 6.090409, 6.210157, 6.329963, 6.449823, 
    6.56974, 6.689711, 6.809736, 6.929816, 7.049948, 7.170134, 7.290371, 
    7.41066, 7.531001, 7.651392, 7.771833, 7.892324, 8.012864, 8.133452, 
    8.254088, 8.374772, 8.495502, 8.61628, 8.737103, 8.85797, 8.978883, 
    9.099839, 9.22084, 9.341883, 9.462969, 9.584096, 9.705265, 9.826475, 
    9.947724, 10.06901, 10.19034, 10.31171, 10.43312, 10.55456, 10.67604, 
    10.79755, 10.9191, 11.04069, 11.16231, 11.28396, 11.40565, 11.52737, 
    11.64912, 11.77091, 11.89272, 12.01457, 12.13644, 12.25835, 12.38028, 
    12.50224, 12.62423, 12.74625, 12.86829, 12.99035, 13.11245, 13.23456, 
    13.3567, 13.47887, 13.60105, 13.72326, 13.84549, 13.96774, 14.09001, 
    14.2123, 14.33461, 14.45694, 14.57928, 14.70165, 14.82403, 14.94642, 
    15.06883, 15.19126, 15.3137, 15.43615, 15.55862, 15.6811, 15.80358, 
    15.92609, 16.0486, 16.17112, 16.29365, 16.41619, 16.53873, 16.66129, 
    16.78385, 16.90642, 17.02899, 17.15157, 17.27415, 17.39673, 17.51932, 
    17.64191, 17.76451, 17.8871, 18.0097, 18.13229, 18.25488, 18.37748, 
    18.50007, 18.62266, 18.74524, 18.86782, 18.9904, 19.11297, 19.23554, 
    19.3581, 19.48065, 19.6032, 19.72573, 19.84826, 19.97078, 20.09329, 
    20.21579, 20.33828, 20.46076, 20.58322, 20.70567, 20.82811, 20.95053, 
    21.07294, 21.19533, 21.31771, 21.44007, 21.56241, 21.68474, 21.80704, 
    21.92933, 22.0516, 22.17385, 22.29607, 22.41828, 22.54046, 22.66262, 
    22.78476, 22.90687, 23.02896, 23.15102, 23.27306, 23.39507, 23.51705, 
    23.63901, 23.76094, 23.88284, 24.00471, 24.12655, 24.24836, 24.37014, 
    24.49188, 24.6136, 24.73528, 24.85693, 24.97855, 25.10013, 25.22167, 
    25.34318, 25.46465, 25.58609, 25.70749, 25.82885, 25.95017, 26.07146, 
    26.1927, 26.3139, 26.43507, 26.55619, 26.67727, 26.7983, 26.9193, 
    27.04025, 27.16115, 27.28201, 27.40283, 27.5236, 27.64432, 27.765, 
    27.88563, 28.00621, 28.12674, 28.24722, 28.36765, 28.48804, 28.60837, 
    28.72865, 28.84888, 28.96906, 29.08918, 29.20925, 29.32927, 29.44923, 
    29.56914, 29.68899, 29.80879, 29.92853, 30.04821, 30.16784, 30.2874, 
    30.40691, 30.52636, 30.64575, 30.76508, 30.88435, 31.00356, 31.12271, 
    31.24179, 31.36082, 31.47977, 31.59867, 31.7175, 31.83627, 31.95498, 
    32.07361, 32.19218, 32.31069, 32.42913, 32.5475, 32.66581, 32.78404, 
    32.90221, 33.02031, 33.13834, 33.25629, 33.37418, 33.492, 33.60975, 
    33.72742, 33.84502, 33.96255, 34.08001, 34.19739, 34.3147, 34.43194, 
    34.5491, 34.66618, 34.78319, 34.90013, 35.01698, 35.13377, 35.25047, 
    35.36709, 35.48364, 35.60011, 35.7165, 35.83281, 35.94904, 36.06519, 
    36.18127, 36.29726, 36.41317, 36.52899, 36.64474, 36.7604, 36.87598, 
    36.99148, 37.10689, 37.22223, 37.33747, 37.45263, 37.56771, 37.6827, 
    37.79761, 37.91243, 38.02716, 38.14181, 38.25637, 38.37084, 38.48523,
  -12.73719, -12.63189, -12.52648, -12.42097, -12.31534, -12.20961, 
    -12.10378, -11.99783, -11.89178, -11.78562, -11.67936, -11.57299, 
    -11.46651, -11.35992, -11.25323, -11.14644, -11.03953, -10.93252, 
    -10.82541, -10.71819, -10.61086, -10.50343, -10.39589, -10.28825, 
    -10.1805, -10.07265, -9.96469, -9.856628, -9.748462, -9.640191, 
    -9.531816, -9.423338, -9.314755, -9.20607, -9.097281, -8.988388, 
    -8.879393, -8.770294, -8.661093, -8.551789, -8.442383, -8.332874, 
    -8.223265, -8.113552, -8.003738, -7.893824, -7.783808, -7.67369, 
    -7.563473, -7.453154, -7.342736, -7.232217, -7.121598, -7.01088, 
    -6.900062, -6.789145, -6.678128, -6.567013, -6.4558, -6.344488, 
    -6.233078, -6.121571, -6.009966, -5.898263, -5.786464, -5.674567, 
    -5.562574, -5.450485, -5.338299, -5.226018, -5.113642, -5.00117, 
    -4.888603, -4.775941, -4.663185, -4.550335, -4.437391, -4.324353, 
    -4.211222, -4.097998, -3.984681, -3.871272, -3.757771, -3.644178, 
    -3.530493, -3.416718, -3.302851, -3.188894, -3.074846, -2.960709, 
    -2.846482, -2.732165, -2.61776, -2.503266, -2.388684, -2.274013, 
    -2.159255, -2.04441, -1.929477, -1.814458, -1.699353, -1.584162, 
    -1.468885, -1.353523, -1.238077, -1.122545, -1.00693, -0.8912305, 
    -0.7754478, -0.6595821, -0.5436337, -0.427603, -0.3114904, -0.1952963, 
    -0.07902107, 0.03733493, 0.1537713, 0.2702877, 0.3868836, 0.5035587, 
    0.6203126, 0.7371449, 0.8540551, 0.9710429, 1.088108, 1.20525, 1.322468, 
    1.439762, 1.557131, 1.674576, 1.792095, 1.909688, 2.027355, 2.145096, 
    2.262909, 2.380795, 2.498753, 2.616783, 2.734884, 2.853055, 2.971297, 
    3.089608, 3.207989, 3.326438, 3.444957, 3.563543, 3.682196, 3.800917, 
    3.919704, 4.038557, 4.157476, 4.27646, 4.395509, 4.514622, 4.633799, 
    4.753038, 4.872341, 4.991705, 5.111132, 5.23062, 5.350168, 5.469777, 
    5.589446, 5.709173, 5.82896, 5.948805, 6.068707, 6.188667, 6.308683, 
    6.428756, 6.548884, 6.669068, 6.789306, 6.909598, 7.029944, 7.150343, 
    7.270794, 7.391298, 7.511853, 7.632459, 7.753115, 7.873821, 7.994576, 
    8.11538, 8.236233, 8.357133, 8.47808, 8.599073, 8.720113, 8.841199, 
    8.962329, 9.083503, 9.204721, 9.325983, 9.447288, 9.568634, 9.690022, 
    9.811451, 9.93292, 10.05443, 10.17598, 10.29756, 10.41919, 10.54085, 
    10.66255, 10.78429, 10.90606, 11.02787, 11.14971, 11.27159, 11.3935, 
    11.51544, 11.63741, 11.75942, 11.88146, 12.00353, 12.12562, 12.24775, 
    12.36991, 12.49209, 12.6143, 12.73654, 12.85881, 12.9811, 13.10342, 
    13.22576, 13.34812, 13.47051, 13.59292, 13.71535, 13.83781, 13.96029, 
    14.08278, 14.2053, 14.32783, 14.45039, 14.57296, 14.69555, 14.81815, 
    14.94077, 15.06341, 15.18606, 15.30873, 15.43141, 15.5541, 15.6768, 
    15.79952, 15.92225, 16.04498, 16.16773, 16.29049, 16.41325, 16.53603, 
    16.65881, 16.7816, 16.90439, 17.02719, 17.15, 17.2728, 17.39562, 
    17.51843, 17.64125, 17.76407, 17.88689, 18.00971, 18.13254, 18.25536, 
    18.37818, 18.50099, 18.62381, 18.74662, 18.86943, 18.99223, 19.11503, 
    19.23783, 19.36061, 19.48339, 19.60617, 19.72893, 19.85169, 19.97443, 
    20.09717, 20.21989, 20.34261, 20.46531, 20.588, 20.71068, 20.83334, 
    20.95599, 21.07863, 21.20124, 21.32385, 21.44643, 21.569, 21.69155, 
    21.81409, 21.9366, 22.05909, 22.18156, 22.30401, 22.42644, 22.54885, 
    22.67124, 22.7936, 22.91593, 23.03825, 23.16053, 23.28279, 23.40503, 
    23.52724, 23.64942, 23.77157, 23.89369, 24.01579, 24.13785, 24.25988, 
    24.38188, 24.50385, 24.62579, 24.74769, 24.86957, 24.9914, 25.1132, 
    25.23497, 25.3567, 25.4784, 25.60005, 25.72167, 25.84325, 25.96479, 
    26.0863, 26.20776, 26.32918, 26.45056, 26.5719, 26.6932, 26.81446, 
    26.93567, 27.05684, 27.17796, 27.29904, 27.42007, 27.54106, 27.66199, 
    27.78289, 27.90373, 28.02453, 28.14528, 28.26597, 28.38662, 28.50722, 
    28.62777, 28.74826, 28.86871, 28.9891, 29.10943, 29.22972, 29.34995, 
    29.47012, 29.59024, 29.7103, 29.83031, 29.95026, 30.07016, 30.18999, 
    30.30977, 30.42949, 30.54915, 30.66875, 30.78829, 30.90776, 31.02718, 
    31.14654, 31.26583, 31.38506, 31.50422, 31.62333, 31.74236, 31.86134, 
    31.98025, 32.09909, 32.21787, 32.33658, 32.45522, 32.5738, 32.6923, 
    32.81074, 32.92911, 33.04741, 33.16564, 33.2838, 33.40189, 33.51991, 
    33.63786, 33.75573, 33.87354, 33.99126, 34.10892, 34.2265, 34.34401, 
    34.46144, 34.5788, 34.69608, 34.81329, 34.93042, 35.04747, 35.16444, 
    35.28134, 35.39816, 35.5149, 35.63157, 35.74815, 35.86465, 35.98108, 
    36.09742, 36.21368, 36.32986, 36.44596, 36.56198, 36.67792, 36.79377, 
    36.90954, 37.02522, 37.14083, 37.25634, 37.37178, 37.48713, 37.60239, 
    37.71757, 37.83266, 37.94766, 38.06258, 38.17741, 38.29216, 38.40681, 
    38.52138,
  -12.78837, -12.68293, -12.57738, -12.47173, -12.36597, -12.26009, 
    -12.15412, -12.04803, -11.94184, -11.83554, -11.72913, -11.62261, 
    -11.51599, -11.40926, -11.30242, -11.19548, -11.08843, -10.98127, 
    -10.87401, -10.76664, -10.65917, -10.55159, -10.4439, -10.33611, 
    -10.22821, -10.1202, -10.0121, -9.903883, -9.795565, -9.687141, 
    -9.578614, -9.469982, -9.361246, -9.252405, -9.143461, -9.034413, 
    -8.925261, -8.816007, -8.706649, -8.597188, -8.487624, -8.377957, 
    -8.268188, -8.158317, -8.048344, -7.938269, -7.828092, -7.717813, 
    -7.607434, -7.496953, -7.386372, -7.27569, -7.164908, -7.054026, 
    -6.943043, -6.831961, -6.720779, -6.609499, -6.498119, -6.386641, 
    -6.275063, -6.163388, -6.051614, -5.939743, -5.827774, -5.715708, 
    -5.603545, -5.491285, -5.378929, -5.266476, -5.153927, -5.041283, 
    -4.928543, -4.815708, -4.702778, -4.589753, -4.476634, -4.363421, 
    -4.250114, -4.136714, -4.023221, -3.909635, -3.795956, -3.682185, 
    -3.568322, -3.454367, -3.340321, -3.226184, -3.111956, -2.997638, 
    -2.883229, -2.768731, -2.654143, -2.539467, -2.424701, -2.309847, 
    -2.194906, -2.079876, -1.964759, -1.849554, -1.734263, -1.618886, 
    -1.503423, -1.387874, -1.272239, -1.15652, -1.040716, -0.9248281, 
    -0.8088561, -0.6928008, -0.5766623, -0.4604411, -0.3441376, -0.2277521, 
    -0.1112851, 0.005263146, 0.1218922, 0.2386016, 0.355391, 0.4722599, 
    0.5892081, 0.7062351, 0.8233405, 0.9405239, 1.057785, 1.175123, 1.292538, 
    1.410029, 1.527596, 1.645238, 1.762956, 1.880748, 1.998614, 2.116554, 
    2.234568, 2.352654, 2.470813, 2.589043, 2.707345, 2.825718, 2.944162, 
    3.062676, 3.18126, 3.299913, 3.418635, 3.537425, 3.656283, 3.775208, 
    3.894201, 4.01326, 4.132384, 4.251575, 4.37083, 4.49015, 4.609534, 
    4.728981, 4.848492, 4.968065, 5.0877, 5.207397, 5.327154, 5.446973, 
    5.566851, 5.68679, 5.806787, 5.926842, 6.046956, 6.167127, 6.287356, 
    6.40764, 6.527981, 6.648377, 6.768829, 6.889335, 7.009894, 7.130507, 
    7.251173, 7.371891, 7.49266, 7.613481, 7.734353, 7.855275, 7.976246, 
    8.097266, 8.218335, 8.339452, 8.460616, 8.581827, 8.703085, 8.824388, 
    8.945736, 9.067128, 9.188565, 9.310046, 9.431569, 9.553135, 9.674743, 
    9.796391, 9.91808, 10.03981, 10.16158, 10.28339, 10.40523, 10.52712, 
    10.64904, 10.771, 10.89299, 11.01502, 11.13708, 11.25918, 11.38131, 
    11.50348, 11.62568, 11.74791, 11.87017, 11.99246, 12.11478, 12.23713, 
    12.35951, 12.48192, 12.60436, 12.72682, 12.84931, 12.97182, 13.09437, 
    13.21693, 13.33952, 13.46214, 13.58477, 13.70743, 13.83011, 13.95281, 
    14.07553, 14.19828, 14.32104, 14.44382, 14.56661, 14.68943, 14.81226, 
    14.93511, 15.05797, 15.18085, 15.30374, 15.42665, 15.54957, 15.6725, 
    15.79544, 15.9184, 16.04136, 16.16434, 16.28732, 16.41031, 16.53332, 
    16.65632, 16.77934, 16.90236, 17.02539, 17.14842, 17.27146, 17.3945, 
    17.51754, 17.64059, 17.76363, 17.88668, 18.00973, 18.13278, 18.25583, 
    18.37888, 18.50192, 18.62497, 18.748, 18.87104, 18.99407, 19.1171, 
    19.24012, 19.36313, 19.48614, 19.60914, 19.73213, 19.85512, 19.97809, 
    20.10106, 20.22401, 20.34695, 20.46988, 20.5928, 20.7157, 20.83859, 
    20.96147, 21.08433, 21.20717, 21.33, 21.45281, 21.57561, 21.69838, 
    21.82114, 21.94388, 22.0666, 22.1893, 22.31197, 22.43463, 22.55726, 
    22.67987, 22.80246, 22.92502, 23.04756, 23.17007, 23.29255, 23.41501, 
    23.53745, 23.65985, 23.78222, 23.90457, 24.02689, 24.14918, 24.27143, 
    24.39366, 24.51585, 24.63801, 24.76014, 24.88223, 25.00429, 25.12631, 
    25.2483, 25.37025, 25.49217, 25.61404, 25.73588, 25.85769, 25.97945, 
    26.10117, 26.22285, 26.3445, 26.4661, 26.58766, 26.70917, 26.83065, 
    26.95208, 27.07346, 27.1948, 27.3161, 27.43735, 27.55855, 27.67971, 
    27.80082, 27.92188, 28.04289, 28.16386, 28.28477, 28.40563, 28.52645, 
    28.64721, 28.76792, 28.88858, 29.00918, 29.12973, 29.25023, 29.37067, 
    29.49106, 29.61139, 29.73167, 29.85188, 29.97205, 30.09215, 30.2122, 
    30.33219, 30.45212, 30.57199, 30.69179, 30.81154, 30.93123, 31.05085, 
    31.17042, 31.28992, 31.40936, 31.52873, 31.64804, 31.76728, 31.88646, 
    32.00558, 32.12463, 32.24361, 32.36252, 32.48137, 32.60015, 32.71886, 
    32.8375, 32.95607, 33.07458, 33.19301, 33.31137, 33.42966, 33.54788, 
    33.66603, 33.7841, 33.90211, 34.02003, 34.13789, 34.25567, 34.37337, 
    34.491, 34.60856, 34.72604, 34.84344, 34.96077, 35.07802, 35.19519, 
    35.31228, 35.4293, 35.54623, 35.66309, 35.77987, 35.89656, 36.01318, 
    36.12971, 36.24617, 36.36254, 36.47883, 36.59504, 36.71117, 36.82721, 
    36.94316, 37.05904, 37.17483, 37.29053, 37.40616, 37.52169, 37.63714, 
    37.75251, 37.86778, 37.98298, 38.09808, 38.21309, 38.32802, 38.44286, 
    38.55761,
  -12.83964, -12.73406, -12.62837, -12.52258, -12.41667, -12.31066, 
    -12.20454, -12.09831, -11.99198, -11.88553, -11.77898, -11.67232, 
    -11.56555, -11.45868, -11.3517, -11.24461, -11.13741, -11.03011, 
    -10.9227, -10.81518, -10.70756, -10.59983, -10.49199, -10.38405, -10.276, 
    -10.16785, -10.05959, -9.951224, -9.842753, -9.734179, -9.625498, 
    -9.516712, -9.407822, -9.298826, -9.189728, -9.080523, -8.971216, 
    -8.861805, -8.75229, -8.642672, -8.532949, -8.423124, -8.313197, 
    -8.203166, -8.093033, -7.982798, -7.87246, -7.762021, -7.651479, 
    -7.540837, -7.430093, -7.319248, -7.208302, -7.097255, -6.986108, 
    -6.874861, -6.763514, -6.652067, -6.540521, -6.428875, -6.31713, 
    -6.205287, -6.093345, -5.981305, -5.869166, -5.75693, -5.644597, 
    -5.532166, -5.419639, -5.307014, -5.194293, -5.081476, -4.968563, 
    -4.855554, -4.74245, -4.629251, -4.515957, -4.402568, -4.289086, 
    -4.175509, -4.061839, -3.948075, -3.834219, -3.720269, -3.606227, 
    -3.492093, -3.377867, -3.26355, -3.149142, -3.034642, -2.920053, 
    -2.805372, -2.690603, -2.575743, -2.460794, -2.345757, -2.23063, 
    -2.115416, -2.000114, -1.884724, -1.769247, -1.653683, -1.538033, 
    -1.422297, -1.306474, -1.190567, -1.074574, -0.9584972, -0.8423358, 
    -0.7260905, -0.6097617, -0.4933496, -0.3768549, -0.2602777, -0.1436186, 
    -0.02687783, 0.08994412, 0.2068469, 0.3238301, 0.4408933, 0.5580361, 
    0.6752582, 0.792559, 0.9099382, 1.027395, 1.14493, 1.262542, 1.380231, 
    1.497995, 1.615836, 1.733752, 1.851744, 1.96981, 2.08795, 2.206163, 
    2.32445, 2.44281, 2.561242, 2.679746, 2.798321, 2.916968, 3.035685, 
    3.154472, 3.273329, 3.392254, 3.511249, 3.630312, 3.749442, 3.86864, 
    3.987905, 4.107236, 4.226633, 4.346095, 4.465622, 4.585214, 4.704869, 
    4.824588, 4.94437, 5.064214, 5.18412, 5.304088, 5.424116, 5.544205, 
    5.664354, 5.784562, 5.90483, 6.025155, 6.145538, 6.265979, 6.386476, 
    6.50703, 6.62764, 6.748304, 6.869024, 6.989798, 7.110625, 7.231505, 
    7.352438, 7.473423, 7.59446, 7.715547, 7.836685, 7.957873, 8.07911, 
    8.200396, 8.32173, 8.443111, 8.564541, 8.686016, 8.807537, 8.929104, 
    9.050715, 9.172372, 9.294071, 9.415814, 9.5376, 9.659427, 9.781296, 
    9.903206, 10.02516, 10.14715, 10.26917, 10.39124, 10.51335, 10.63549, 
    10.75767, 10.87989, 11.00214, 11.12442, 11.24675, 11.3691, 11.49149, 
    11.61391, 11.73636, 11.85885, 11.98136, 12.10391, 12.22648, 12.34909, 
    12.47172, 12.59438, 12.71707, 12.83979, 12.96253, 13.08529, 13.20809, 
    13.3309, 13.45374, 13.5766, 13.69949, 13.82239, 13.94532, 14.06827, 
    14.19124, 14.31422, 14.43723, 14.56025, 14.6833, 14.80635, 14.92943, 
    15.05252, 15.17562, 15.29875, 15.42188, 15.54502, 15.66818, 15.79136, 
    15.91454, 16.03773, 16.16093, 16.28415, 16.40737, 16.5306, 16.65383, 
    16.77708, 16.90033, 17.02358, 17.14684, 17.27011, 17.39337, 17.51665, 
    17.63992, 17.7632, 17.88647, 18.00975, 18.13303, 18.25631, 18.37958, 
    18.50285, 18.62613, 18.74939, 18.87266, 18.99592, 19.11917, 19.24242, 
    19.36566, 19.4889, 19.61213, 19.73535, 19.85856, 19.98176, 20.10495, 
    20.22813, 20.3513, 20.47445, 20.5976, 20.72073, 20.84385, 20.96695, 
    21.09004, 21.21311, 21.33617, 21.45921, 21.58223, 21.70523, 21.82822, 
    21.95118, 22.07413, 22.19705, 22.31995, 22.44283, 22.56569, 22.68853, 
    22.81134, 22.93413, 23.05689, 23.17963, 23.30234, 23.42502, 23.54768, 
    23.67031, 23.79291, 23.91548, 24.03802, 24.16053, 24.28301, 24.40546, 
    24.52787, 24.65026, 24.77261, 24.89492, 25.0172, 25.13945, 25.26166, 
    25.38383, 25.50597, 25.62807, 25.75013, 25.87215, 25.99414, 26.11608, 
    26.23798, 26.35985, 26.48167, 26.60345, 26.72518, 26.84688, 26.96852, 
    27.09013, 27.21169, 27.3332, 27.45467, 27.57609, 27.69747, 27.81879, 
    27.94007, 28.0613, 28.18248, 28.30361, 28.42469, 28.54572, 28.66669, 
    28.78762, 28.90849, 29.02931, 29.15008, 29.27079, 29.39144, 29.51204, 
    29.63259, 29.75308, 29.87351, 29.99388, 30.1142, 30.23446, 30.35466, 
    30.47479, 30.59487, 30.71489, 30.83485, 30.95475, 31.07458, 31.19435, 
    31.31406, 31.43371, 31.55329, 31.67281, 31.79226, 31.91164, 32.03096, 
    32.15022, 32.26941, 32.38853, 32.50758, 32.62656, 32.74548, 32.86432, 
    32.9831, 33.10181, 33.22044, 33.339, 33.4575, 33.57592, 33.69427, 
    33.81254, 33.93074, 34.04887, 34.16693, 34.2849, 34.40281, 34.52064, 
    34.63839, 34.75607, 34.87367, 34.99119, 35.10863, 35.226, 35.34329, 
    35.4605, 35.57763, 35.69468, 35.81165, 35.92854, 36.04535, 36.16208, 
    36.27872, 36.39529, 36.51177, 36.62817, 36.74448, 36.86072, 36.97686, 
    37.09293, 37.20891, 37.3248, 37.44061, 37.55633, 37.67197, 37.78752, 
    37.90298, 38.01836, 38.13365, 38.24885, 38.36396, 38.47898, 38.59392,
  -12.891, -12.78528, -12.67945, -12.57352, -12.46747, -12.36132, -12.25506, 
    -12.14869, -12.04221, -11.93562, -11.82892, -11.72212, -11.61521, 
    -11.50819, -11.40106, -11.29383, -11.18648, -11.07903, -10.97147, 
    -10.86381, -10.75604, -10.64816, -10.54017, -10.43208, -10.32388, 
    -10.21558, -10.10717, -9.998652, -9.89003, -9.781301, -9.672467, 
    -9.563528, -9.454483, -9.345334, -9.236079, -9.12672, -9.017257, 
    -8.907689, -8.798017, -8.688241, -8.578361, -8.468377, -8.358291, 
    -8.2481, -8.137808, -8.027411, -7.916913, -7.806312, -7.695609, 
    -7.584804, -7.473897, -7.362889, -7.251779, -7.140568, -7.029256, 
    -6.917844, -6.806331, -6.694718, -6.583005, -6.471192, -6.35928, 
    -6.247269, -6.135158, -6.022949, -5.910641, -5.798235, -5.685731, 
    -5.573129, -5.46043, -5.347633, -5.23474, -5.12175, -5.008664, -4.895481, 
    -4.782203, -4.668829, -4.555359, -4.441795, -4.328136, -4.214383, 
    -4.100536, -3.986594, -3.87256, -3.758432, -3.644211, -3.529898, 
    -3.415492, -3.300994, -3.186405, -3.071724, -2.956953, -2.84209, 
    -2.727138, -2.612095, -2.496963, -2.381741, -2.26643, -2.151031, 
    -2.035543, -1.919968, -1.804304, -1.688554, -1.572717, -1.456793, 
    -1.340782, -1.224687, -1.108505, -0.9922385, -0.8758873, -0.7594517, 
    -0.6429321, -0.526329, -0.4096427, -0.2928736, -0.176022, -0.05908844, 
    0.05792679, 0.1750232, 0.2922005, 0.4094583, 0.526796, 0.6442134, 
    0.76171, 0.8792855, 0.9969393, 1.114671, 1.23248, 1.350367, 1.46833, 
    1.586369, 1.704485, 1.822675, 1.940941, 2.059281, 2.177696, 2.296183, 
    2.414744, 2.533378, 2.652085, 2.770863, 2.889712, 3.008632, 3.127623, 
    3.246684, 3.365814, 3.485014, 3.604282, 3.723618, 3.843022, 3.962493, 
    4.082031, 4.201634, 4.321304, 4.441039, 4.560839, 4.680703, 4.80063, 
    4.920621, 5.040675, 5.160791, 5.280969, 5.401207, 5.521507, 5.641867, 
    5.762287, 5.882766, 6.003303, 6.123899, 6.244553, 6.365263, 6.48603, 
    6.606853, 6.727732, 6.848666, 6.969654, 7.090696, 7.211792, 7.332941, 
    7.454141, 7.575394, 7.696698, 7.818052, 7.939457, 8.060911, 8.182415, 
    8.303967, 8.425566, 8.547214, 8.668907, 8.790648, 8.912433, 9.034264, 
    9.156139, 9.278059, 9.400022, 9.522028, 9.644075, 9.766165, 9.888296, 
    10.01047, 10.13268, 10.25493, 10.37722, 10.49955, 10.62191, 10.74431, 
    10.86675, 10.98923, 11.11174, 11.23428, 11.35686, 11.47947, 11.60212, 
    11.72479, 11.8475, 11.97024, 12.09301, 12.21581, 12.33864, 12.4615, 
    12.58439, 12.7073, 12.83024, 12.95321, 13.0762, 13.19922, 13.32226, 
    13.44532, 13.56841, 13.69152, 13.81466, 13.93781, 14.06099, 14.18418, 
    14.30739, 14.43063, 14.55388, 14.67715, 14.80044, 14.92374, 15.04706, 
    15.17039, 15.29374, 15.4171, 15.54047, 15.66386, 15.78726, 15.91067, 
    16.03409, 16.15752, 16.28096, 16.40441, 16.52787, 16.65133, 16.77481, 
    16.89828, 17.02177, 17.14526, 17.26875, 17.39225, 17.51575, 17.63925, 
    17.76276, 17.88626, 18.00977, 18.13327, 18.25678, 18.38029, 18.50379, 
    18.62729, 18.75078, 18.87428, 18.99776, 19.12125, 19.24472, 19.3682, 
    19.49166, 19.61512, 19.73856, 19.862, 19.98543, 20.10885, 20.23226, 
    20.35566, 20.47904, 20.60242, 20.72578, 20.84912, 20.97245, 21.09577, 
    21.21907, 21.34235, 21.46562, 21.58887, 21.7121, 21.83531, 21.9585, 
    22.08167, 22.20482, 22.32795, 22.45106, 22.57414, 22.69721, 22.82024, 
    22.94326, 23.06625, 23.18921, 23.31215, 23.43505, 23.55794, 23.68079, 
    23.80361, 23.92641, 24.04918, 24.17191, 24.29461, 24.41729, 24.53993, 
    24.66253, 24.78511, 24.90764, 25.03015, 25.15262, 25.27505, 25.39745, 
    25.51981, 25.64213, 25.76441, 25.88666, 26.00886, 26.13103, 26.25315, 
    26.37523, 26.49727, 26.61927, 26.74123, 26.86314, 26.98501, 27.10683, 
    27.22861, 27.35035, 27.47203, 27.59367, 27.71527, 27.83681, 27.9583, 
    28.07975, 28.20115, 28.32249, 28.44379, 28.56503, 28.68623, 28.80737, 
    28.92845, 29.04949, 29.17047, 29.29139, 29.41226, 29.53308, 29.65384, 
    29.77454, 29.89518, 30.01577, 30.1363, 30.25677, 30.37718, 30.49753, 
    30.61782, 30.73805, 30.85821, 30.97832, 31.09836, 31.21835, 31.33826, 
    31.45812, 31.57791, 31.69763, 31.81729, 31.93688, 32.05641, 32.17587, 
    32.29527, 32.41459, 32.53385, 32.65303, 32.77216, 32.8912, 33.01019, 
    33.12909, 33.24793, 33.3667, 33.48539, 33.60402, 33.72256, 33.84104, 
    33.95944, 34.07777, 34.19603, 34.31421, 34.43231, 34.55033, 34.66829, 
    34.78616, 34.90396, 35.02168, 35.13932, 35.25688, 35.37437, 35.49177, 
    35.6091, 35.72634, 35.84351, 35.96059, 36.07759, 36.19451, 36.31135, 
    36.4281, 36.54478, 36.66137, 36.77787, 36.8943, 37.01064, 37.12689, 
    37.24306, 37.35914, 37.47514, 37.59105, 37.70687, 37.82261, 37.93826, 
    38.05382, 38.16929, 38.28468, 38.39997, 38.51518, 38.6303,
  -12.94244, -12.83658, -12.73062, -12.62454, -12.51836, -12.41206, 
    -12.30566, -12.19915, -12.09252, -11.98579, -11.87895, -11.77201, 
    -11.66495, -11.55779, -11.45051, -11.34313, -11.23564, -11.12804, 
    -11.02034, -10.91253, -10.80461, -10.69658, -10.58844, -10.4802, 
    -10.37185, -10.2634, -10.15484, -10.04617, -9.937392, -9.828511, 
    -9.719524, -9.610431, -9.501232, -9.391928, -9.282518, -9.173004, 
    -9.063384, -8.953659, -8.84383, -8.733896, -8.623858, -8.513717, 
    -8.40347, -8.29312, -8.182668, -8.072111, -7.961452, -7.850689, 
    -7.739824, -7.628857, -7.517787, -7.406615, -7.295341, -7.183966, 
    -7.072489, -6.960911, -6.849233, -6.737453, -6.625573, -6.513593, 
    -6.401513, -6.289333, -6.177054, -6.064675, -5.952198, -5.839622, 
    -5.726947, -5.614174, -5.501303, -5.388335, -5.275269, -5.162106, 
    -5.048845, -4.935489, -4.822036, -4.708487, -4.594842, -4.481102, 
    -4.367267, -4.253337, -4.139312, -4.025193, -3.91098, -3.796673, 
    -3.682273, -3.56778, -3.453194, -3.338516, -3.223746, -3.108884, 
    -2.99393, -2.878885, -2.76375, -2.648524, -2.533207, -2.417802, 
    -2.302306, -2.186722, -2.071048, -1.955287, -1.839437, -1.723499, 
    -1.607474, -1.491362, -1.375164, -1.258879, -1.142509, -1.026052, 
    -0.9095109, -0.7928848, -0.6761743, -0.5593797, -0.4425015, -0.3255401, 
    -0.2084958, -0.09136911, 0.02583969, 0.1431302, 0.2605019, 0.3779545, 
    0.4954875, 0.6131006, 0.7307934, 0.8485653, 0.9664161, 1.084345, 
    1.202352, 1.320437, 1.438599, 1.556837, 1.675152, 1.793542, 1.912008, 
    2.030549, 2.149164, 2.267853, 2.386616, 2.505452, 2.624361, 2.743342, 
    2.862395, 2.981519, 3.100714, 3.219979, 3.339314, 3.458719, 3.578193, 
    3.697735, 3.817345, 3.937023, 4.056767, 4.176579, 4.296456, 4.416399, 
    4.536407, 4.65648, 4.776617, 4.896818, 5.017081, 5.137407, 5.257796, 
    5.378246, 5.498757, 5.619328, 5.73996, 5.860651, 5.981401, 6.10221, 
    6.223076, 6.344, 6.464982, 6.586019, 6.707112, 6.82826, 6.949464, 
    7.070722, 7.192033, 7.313397, 7.434814, 7.556283, 7.677804, 7.799376, 
    7.920998, 8.042669, 8.164391, 8.286161, 8.407979, 8.529845, 8.651758, 
    8.773717, 8.895722, 9.017774, 9.139869, 9.262009, 9.384192, 9.506418, 
    9.628688, 9.750998, 9.873351, 9.995744, 10.11818, 10.24065, 10.36316, 
    10.48571, 10.6083, 10.73092, 10.85359, 10.97628, 11.09902, 11.22179, 
    11.34459, 11.46743, 11.59029, 11.7132, 11.83613, 11.95909, 12.08209, 
    12.20512, 12.32817, 12.45125, 12.57437, 12.6975, 12.82067, 12.94386, 
    13.06708, 13.19033, 13.31359, 13.43689, 13.5602, 13.68354, 13.8069, 
    13.93028, 14.05369, 14.17711, 14.30055, 14.42401, 14.54749, 14.67099, 
    14.7945, 14.91803, 15.04158, 15.16514, 15.28872, 15.41231, 15.53591, 
    15.65952, 15.78315, 15.90679, 16.03044, 16.1541, 16.27777, 16.40145, 
    16.52514, 16.64883, 16.77253, 16.89624, 17.01995, 17.14367, 17.26739, 
    17.39112, 17.51485, 17.63858, 17.76232, 17.88605, 18.00979, 18.13352, 
    18.25726, 18.38099, 18.50472, 18.62845, 18.75218, 18.8759, 18.99962, 
    19.12333, 19.24704, 19.37074, 19.49443, 19.61811, 19.74179, 19.86546, 
    19.98912, 20.11277, 20.2364, 20.36003, 20.48364, 20.60724, 20.73083, 
    20.85441, 20.97797, 21.10151, 21.22504, 21.34855, 21.47204, 21.59552, 
    21.71898, 21.84242, 21.96584, 22.08924, 22.21261, 22.33597, 22.4593, 
    22.58262, 22.70591, 22.82917, 22.95241, 23.07562, 23.19881, 23.32198, 
    23.44511, 23.56822, 23.6913, 23.81435, 23.93737, 24.06036, 24.18332, 
    24.30625, 24.42914, 24.55201, 24.67484, 24.79764, 24.9204, 25.04313, 
    25.16582, 25.28848, 25.41109, 25.53368, 25.65622, 25.77873, 25.90119, 
    26.02362, 26.14601, 26.26835, 26.39066, 26.51292, 26.63514, 26.75731, 
    26.87945, 27.00154, 27.12358, 27.24558, 27.36753, 27.48944, 27.61129, 
    27.7331, 27.85487, 27.97658, 28.09824, 28.21986, 28.34142, 28.46293, 
    28.5844, 28.7058, 28.82716, 28.94846, 29.06971, 29.19091, 29.31205, 
    29.43313, 29.55416, 29.67513, 29.79605, 29.9169, 30.0377, 30.15845, 
    30.27913, 30.39975, 30.52031, 30.64081, 30.76125, 30.88163, 31.00195, 
    31.1222, 31.24239, 31.36252, 31.48258, 31.60258, 31.72251, 31.84238, 
    31.96218, 32.08191, 32.20158, 32.32118, 32.44071, 32.56017, 32.67957, 
    32.79889, 32.91814, 33.03733, 33.15644, 33.27548, 33.39445, 33.51335, 
    33.63218, 33.75093, 33.8696, 33.98821, 34.10674, 34.22519, 34.34357, 
    34.46187, 34.5801, 34.69825, 34.81632, 34.93431, 35.05223, 35.17007, 
    35.28783, 35.40551, 35.52311, 35.64063, 35.75807, 35.87543, 35.99271, 
    36.1099, 36.22702, 36.34405, 36.46099, 36.57786, 36.69464, 36.81134, 
    36.92795, 37.04448, 37.16092, 37.27728, 37.39355, 37.50974, 37.62583, 
    37.74184, 37.85777, 37.9736, 38.08935, 38.20501, 38.32058, 38.43606, 
    38.55146, 38.66676,
  -12.99397, -12.88798, -12.78187, -12.67566, -12.56933, -12.46289, 
    -12.35635, -12.24969, -12.14293, -12.03606, -11.92907, -11.82198, 
    -11.71478, -11.60747, -11.50005, -11.39252, -11.28489, -11.17714, 
    -11.06929, -10.96133, -10.85326, -10.74509, -10.6368, -10.52841, 
    -10.41991, -10.3113, -10.20259, -10.09377, -9.984843, -9.875809, 
    -9.766668, -9.657421, -9.548068, -9.438609, -9.329044, -9.219374, 
    -9.109598, -8.999717, -8.88973, -8.779638, -8.669442, -8.559141, 
    -8.448736, -8.338227, -8.227613, -8.116897, -8.006076, -7.895152, 
    -7.784125, -7.672995, -7.561761, -7.450426, -7.338988, -7.227448, 
    -7.115807, -7.004063, -6.892219, -6.780272, -6.668226, -6.556078, 
    -6.44383, -6.331481, -6.219033, -6.106485, -5.993838, -5.881092, 
    -5.768246, -5.655302, -5.542259, -5.429118, -5.315879, -5.202543, 
    -5.089109, -4.975578, -4.86195, -4.748227, -4.634406, -4.52049, 
    -4.406478, -4.292371, -4.178168, -4.063871, -3.94948, -3.834994, 
    -3.720415, -3.605742, -3.490975, -3.376116, -3.261165, -3.146121, 
    -3.030985, -2.915757, -2.800439, -2.685029, -2.569529, -2.453938, 
    -2.338258, -2.222488, -2.106629, -1.99068, -1.874644, -1.758519, 
    -1.642306, -1.526006, -1.409619, -1.293145, -1.176585, -1.059939, 
    -0.9432073, -0.8263903, -0.7094885, -0.5925022, -0.4754318, -0.3582778, 
    -0.2410405, -0.1237203, -0.006317614, 0.1111672, 0.2287337, 0.3463815, 
    0.4641101, 0.5819193, 0.6998084, 0.8177772, 0.9358253, 1.053952, 
    1.172157, 1.290441, 1.408801, 1.527239, 1.645753, 1.764344, 1.883011, 
    2.001752, 2.120569, 2.23946, 2.358425, 2.477464, 2.596575, 2.71576, 
    2.835016, 2.954344, 3.073744, 3.193214, 3.312754, 3.432365, 3.552044, 
    3.671793, 3.79161, 3.911495, 4.031447, 4.151466, 4.271552, 4.391704, 
    4.51192, 4.632203, 4.752549, 4.87296, 4.993433, 5.11397, 5.23457, 
    5.355231, 5.475954, 5.596737, 5.717581, 5.838485, 5.959448, 6.08047, 
    6.20155, 6.322688, 6.443883, 6.565135, 6.686444, 6.807807, 6.929226, 
    7.0507, 7.172227, 7.293808, 7.415442, 7.537128, 7.658866, 7.780655, 
    7.902495, 8.024385, 8.146325, 8.268313, 8.39035, 8.512436, 8.634568, 
    8.756747, 8.878973, 9.001244, 9.12356, 9.24592, 9.368324, 9.490772, 
    9.613263, 9.735795, 9.85837, 9.980985, 10.10364, 10.22634, 10.34907, 
    10.47184, 10.59466, 10.7175, 10.84039, 10.96331, 11.08627, 11.20926, 
    11.33229, 11.45535, 11.57844, 11.70157, 11.82473, 11.94792, 12.07114, 
    12.19439, 12.31767, 12.44098, 12.56432, 12.68769, 12.81108, 12.9345, 
    13.05795, 13.18142, 13.30491, 13.42843, 13.55197, 13.67554, 13.79913, 
    13.92274, 14.04637, 14.17002, 14.29369, 14.41738, 14.54109, 14.66481, 
    14.78855, 14.91231, 15.03609, 15.15988, 15.28368, 15.4075, 15.53133, 
    15.65518, 15.77904, 15.90291, 16.02678, 16.15067, 16.27457, 16.39848, 
    16.5224, 16.64632, 16.77025, 16.89419, 17.01813, 17.14208, 17.26603, 
    17.38999, 17.51395, 17.63791, 17.76188, 17.88584, 18.00981, 18.13377, 
    18.25773, 18.3817, 18.50566, 18.62962, 18.75357, 18.87753, 19.00147, 
    19.12542, 19.24935, 19.37328, 19.4972, 19.62112, 19.74503, 19.86892, 
    19.99281, 20.11669, 20.24056, 20.36441, 20.48825, 20.61209, 20.7359, 
    20.8597, 20.98349, 21.10727, 21.23102, 21.35476, 21.47849, 21.60219, 
    21.72588, 21.84954, 21.97319, 22.09682, 22.22042, 22.34401, 22.46757, 
    22.59111, 22.71463, 22.83812, 22.96158, 23.08503, 23.20844, 23.33183, 
    23.45519, 23.57853, 23.70183, 23.82511, 23.94835, 24.07157, 24.19476, 
    24.31791, 24.44103, 24.56412, 24.68717, 24.8102, 24.93318, 25.05614, 
    25.17905, 25.30193, 25.42477, 25.54758, 25.67035, 25.79308, 25.91576, 
    26.03841, 26.16102, 26.28359, 26.40612, 26.5286, 26.65104, 26.77344, 
    26.89579, 27.0181, 27.14036, 27.26258, 27.38475, 27.50688, 27.62896, 
    27.75099, 27.87297, 27.9949, 28.11678, 28.23861, 28.3604, 28.48212, 
    28.6038, 28.72543, 28.847, 28.96852, 29.08998, 29.21139, 29.33275, 
    29.45405, 29.57529, 29.69648, 29.81761, 29.93868, 30.05969, 30.18064, 
    30.30154, 30.42237, 30.54315, 30.66386, 30.78451, 30.9051, 31.02563, 
    31.14609, 31.26649, 31.38683, 31.5071, 31.62731, 31.74745, 31.86752, 
    31.98753, 32.10748, 32.22735, 32.34715, 32.46689, 32.58656, 32.70616, 
    32.82569, 32.94515, 33.06454, 33.18385, 33.3031, 33.42227, 33.54137, 
    33.6604, 33.77935, 33.89823, 34.01704, 34.13577, 34.25442, 34.373, 
    34.4915, 34.60993, 34.72828, 34.84655, 34.96474, 35.08286, 35.20089, 
    35.31884, 35.43672, 35.55452, 35.67223, 35.78987, 35.90742, 36.02489, 
    36.14228, 36.25959, 36.37682, 36.49396, 36.61101, 36.72799, 36.84488, 
    36.96168, 37.0784, 37.19503, 37.31158, 37.42804, 37.54441, 37.66069, 
    37.77689, 37.89301, 38.00903, 38.12496, 38.24081, 38.35656, 38.47223, 
    38.58781, 38.70329,
  -13.0456, -12.93946, -12.83322, -12.72686, -12.62039, -12.51382, -12.40713, 
    -12.30033, -12.19342, -12.08641, -11.97928, -11.87204, -11.7647, 
    -11.65724, -11.54968, -11.44201, -11.33422, -11.22633, -11.11833, 
    -11.01022, -10.90201, -10.79368, -10.68525, -10.57671, -10.46806, 
    -10.3593, -10.25043, -10.14146, -10.03238, -9.923195, -9.813901, -9.7045, 
    -9.594993, -9.485378, -9.375658, -9.265832, -9.155899, -9.045861, 
    -8.935718, -8.825468, -8.715114, -8.604653, -8.494089, -8.38342, 
    -8.272647, -8.161769, -8.050787, -7.939701, -7.828511, -7.717218, 
    -7.605822, -7.494323, -7.382721, -7.271016, -7.159209, -7.0473, 
    -6.935289, -6.823176, -6.710962, -6.598647, -6.486231, -6.373714, 
    -6.261097, -6.148379, -6.035562, -5.922645, -5.809628, -5.696512, 
    -5.583297, -5.469984, -5.356572, -5.243062, -5.129455, -5.015749, 
    -4.901947, -4.788047, -4.674051, -4.559958, -4.44577, -4.331485, 
    -4.217105, -4.10263, -3.98806, -3.873395, -3.758636, -3.643782, 
    -3.528836, -3.413795, -3.298662, -3.183436, -3.068118, -2.952708, 
    -2.837205, -2.721612, -2.605927, -2.490152, -2.374286, -2.25833, 
    -2.142285, -2.02615, -1.909926, -1.793614, -1.677213, -1.560725, 
    -1.444149, -1.327486, -1.210736, -1.093899, -0.9769768, -0.8599686, 
    -0.7428752, -0.6256969, -0.5084341, -0.3910871, -0.2736565, -0.1561425, 
    -0.03854556, 0.07913388, 0.1968955, 0.3147388, 0.4326634, 0.5506688, 
    0.6687548, 0.7869208, 0.9051665, 1.023491, 1.141895, 1.260377, 1.378937, 
    1.497575, 1.616289, 1.73508, 1.853948, 1.972891, 2.091909, 2.211002, 
    2.33017, 2.449412, 2.568727, 2.688115, 2.807575, 2.927108, 3.046712, 
    3.166388, 3.286134, 3.40595, 3.525836, 3.645792, 3.765816, 3.885908, 
    4.006068, 4.126296, 4.24659, 4.366951, 4.487377, 4.607869, 4.728425, 
    4.849046, 4.969731, 5.090478, 5.211289, 5.332162, 5.453097, 5.574093, 
    5.69515, 5.816267, 5.937444, 6.058679, 6.179974, 6.301326, 6.422736, 
    6.544203, 6.665727, 6.787306, 6.908941, 7.030631, 7.152375, 7.274172, 
    7.396023, 7.517927, 7.639883, 7.76189, 7.883948, 8.006057, 8.128216, 
    8.250423, 8.37268, 8.494985, 8.617337, 8.739737, 8.862183, 8.984674, 
    9.107211, 9.229794, 9.352419, 9.475088, 9.597801, 9.720556, 9.843352, 
    9.96619, 10.08907, 10.21199, 10.33495, 10.45794, 10.58098, 10.70405, 
    10.82716, 10.95031, 11.07349, 11.19671, 11.31996, 11.44324, 11.56656, 
    11.68992, 11.8133, 11.93672, 12.06016, 12.18364, 12.30715, 12.43069, 
    12.55425, 12.67784, 12.80147, 12.92511, 13.04878, 13.17248, 13.29621, 
    13.41995, 13.54372, 13.66752, 13.79133, 13.91517, 14.03903, 14.16291, 
    14.28681, 14.41073, 14.53466, 14.65862, 14.78259, 14.90658, 15.03058, 
    15.1546, 15.27864, 15.40269, 15.52675, 15.65082, 15.77491, 15.89901, 
    16.02312, 16.14724, 16.27137, 16.39551, 16.51965, 16.64381, 16.76797, 
    16.89213, 17.01631, 17.14049, 17.26467, 17.38885, 17.51304, 17.63724, 
    17.76143, 17.88563, 18.00982, 18.13402, 18.25821, 18.38241, 18.5066, 
    18.63079, 18.75498, 18.87916, 19.00334, 19.12751, 19.25167, 19.37583, 
    19.49999, 19.62413, 19.74827, 19.8724, 19.99652, 20.12062, 20.24472, 
    20.3688, 20.49288, 20.61694, 20.74098, 20.86502, 20.98903, 21.11304, 
    21.23702, 21.36099, 21.48494, 21.60888, 21.73279, 21.85669, 21.98056, 
    22.10442, 22.22825, 22.35207, 22.47585, 22.59962, 22.72337, 22.84709, 
    22.97078, 23.09445, 23.21809, 23.34171, 23.4653, 23.58886, 23.71239, 
    23.83589, 23.95936, 24.08281, 24.20622, 24.3296, 24.45295, 24.57626, 
    24.69954, 24.82279, 24.946, 25.06918, 25.19232, 25.31542, 25.43849, 
    25.56152, 25.68451, 25.80746, 25.93037, 26.05324, 26.17607, 26.29886, 
    26.42161, 26.54432, 26.66698, 26.7896, 26.91217, 27.0347, 27.15719, 
    27.27963, 27.40202, 27.52436, 27.64666, 27.76891, 27.89111, 28.01326, 
    28.13536, 28.25741, 28.37941, 28.50136, 28.62325, 28.7451, 28.86689, 
    28.98862, 29.1103, 29.23193, 29.3535, 29.47502, 29.59647, 29.71787, 
    29.83922, 29.9605, 30.08173, 30.2029, 30.324, 30.44505, 30.56604, 
    30.68696, 30.80783, 30.92863, 31.04936, 31.17004, 31.29065, 31.4112, 
    31.53168, 31.65209, 31.77244, 31.89273, 32.01294, 32.13309, 32.25317, 
    32.37319, 32.49313, 32.61301, 32.73281, 32.85255, 32.97221, 33.0918, 
    33.21133, 33.33078, 33.45015, 33.56945, 33.68869, 33.80784, 33.92692, 
    34.04593, 34.16486, 34.28371, 34.4025, 34.5212, 34.63982, 34.75837, 
    34.87684, 34.99523, 35.11354, 35.23178, 35.34993, 35.468, 35.58599, 
    35.70391, 35.82174, 35.93949, 36.05715, 36.17474, 36.29224, 36.40966, 
    36.52699, 36.64424, 36.7614, 36.87848, 36.99548, 37.11238, 37.22921, 
    37.34595, 37.4626, 37.57916, 37.69563, 37.81202, 37.92832, 38.04453, 
    38.16065, 38.27668, 38.39262, 38.50847, 38.62423, 38.7399,
  -13.09731, -12.99104, -12.88465, -12.77815, -12.67155, -12.56483, -12.458, 
    -12.35106, -12.24401, -12.13685, -12.02958, -11.9222, -11.81471, 
    -11.70711, -11.5994, -11.49158, -11.38365, -11.27561, -11.16746, 
    -11.05921, -10.95084, -10.84237, -10.73378, -10.62509, -10.51629, 
    -10.40738, -10.29837, -10.18924, -10.08001, -9.97067, -9.861222, 
    -9.751667, -9.642005, -9.532236, -9.42236, -9.312378, -9.202289, 
    -9.092093, -8.981792, -8.871386, -8.760872, -8.650253, -8.53953, -8.4287, 
    -8.317766, -8.206728, -8.095584, -7.984336, -7.872984, -7.761528, 
    -7.649969, -7.538306, -7.426539, -7.31467, -7.202698, -7.090623, 
    -6.978446, -6.866166, -6.753785, -6.641302, -6.528717, -6.416031, 
    -6.303245, -6.190357, -6.07737, -5.964282, -5.851094, -5.737806, 
    -5.624419, -5.510933, -5.397348, -5.283665, -5.169883, -5.056003, 
    -4.942025, -4.82795, -4.713778, -4.599509, -4.485143, -4.370681, 
    -4.256123, -4.141469, -4.02672, -3.911875, -3.796937, -3.681903, 
    -3.566775, -3.451554, -3.336239, -3.22083, -3.105329, -2.989736, 
    -2.87405, -2.758272, -2.642403, -2.526443, -2.410391, -2.29425, 
    -2.178018, -2.061696, -1.945285, -1.828785, -1.712196, -1.595518, 
    -1.478753, -1.3619, -1.24496, -1.127933, -1.01082, -0.8936203, 
    -0.7763349, -0.6589643, -0.5415087, -0.4239685, -0.3063442, -0.1886361, 
    -0.07084461, 0.04702981, 0.1649868, 0.2830259, 0.4011468, 0.519349, 
    0.6376321, 0.7559957, 0.8744393, 0.9929626, 1.111565, 1.230246, 1.349006, 
    1.467844, 1.586759, 1.705751, 1.824819, 1.943964, 2.063185, 2.18248, 
    2.301851, 2.421296, 2.540814, 2.660407, 2.780072, 2.899809, 3.019619, 
    3.1395, 3.259452, 3.379475, 3.499568, 3.61973, 3.739962, 3.860262, 
    3.980631, 4.101067, 4.22157, 4.34214, 4.462776, 4.583478, 4.704245, 
    4.825077, 4.945973, 5.066932, 5.187955, 5.30904, 5.430188, 5.551396, 
    5.672667, 5.793997, 5.915388, 6.036838, 6.158346, 6.279914, 6.401539, 
    6.523221, 6.644961, 6.766757, 6.888608, 7.010514, 7.132475, 7.25449, 
    7.376559, 7.498681, 7.620854, 7.74308, 7.865357, 7.987685, 8.110064, 
    8.232491, 8.354967, 8.477492, 8.600065, 8.722686, 8.845352, 8.968065, 
    9.090824, 9.213628, 9.336475, 9.459367, 9.582302, 9.705279, 9.8283, 
    9.951361, 10.07446, 10.19761, 10.32079, 10.44401, 10.56727, 10.69057, 
    10.8139, 10.93727, 11.06068, 11.18412, 11.3076, 11.43111, 11.55466, 
    11.67824, 11.80185, 11.92549, 12.04916, 12.17287, 12.2966, 12.42037, 
    12.54416, 12.66798, 12.79183, 12.9157, 13.0396, 13.16353, 13.28748, 
    13.41146, 13.53545, 13.65948, 13.78352, 13.90759, 14.03168, 14.15579, 
    14.27991, 14.40406, 14.52823, 14.65241, 14.77661, 14.90083, 15.02507, 
    15.14932, 15.27358, 15.39786, 15.52215, 15.64646, 15.77077, 15.8951, 
    16.01944, 16.14379, 16.26815, 16.39252, 16.5169, 16.64128, 16.76568, 
    16.89007, 17.01448, 17.13889, 17.2633, 17.38772, 17.51214, 17.63656, 
    17.76099, 17.88541, 18.00984, 18.13427, 18.25869, 18.38312, 18.50754, 
    18.63196, 18.75638, 18.88079, 19.0052, 19.1296, 19.254, 19.37839, 
    19.50278, 19.62715, 19.75152, 19.87588, 20.00023, 20.12457, 20.24889, 
    20.37321, 20.49751, 20.6218, 20.74608, 20.87034, 20.99459, 21.11882, 
    21.24303, 21.36723, 21.49142, 21.61558, 21.73972, 21.86385, 21.98795, 
    22.11204, 22.2361, 22.36014, 22.48416, 22.60816, 22.73213, 22.85608, 
    22.98, 23.1039, 23.22777, 23.35161, 23.47543, 23.59921, 23.72297, 
    23.8467, 23.9704, 24.09407, 24.21771, 24.34132, 24.46489, 24.58843, 
    24.71194, 24.83541, 24.95885, 25.08225, 25.20561, 25.32894, 25.45223, 
    25.57549, 25.6987, 25.82188, 25.94501, 26.06811, 26.19116, 26.31418, 
    26.43715, 26.56008, 26.68296, 26.8058, 26.9286, 27.05135, 27.17406, 
    27.29671, 27.41933, 27.54189, 27.66441, 27.78688, 27.9093, 28.03167, 
    28.15399, 28.27626, 28.39848, 28.52064, 28.64275, 28.76481, 28.88682, 
    29.00877, 29.13067, 29.25251, 29.3743, 29.49603, 29.6177, 29.73932, 
    29.86088, 29.98238, 30.10382, 30.2252, 30.34652, 30.46778, 30.58898, 
    30.71012, 30.83119, 30.95221, 31.07315, 31.19404, 31.31486, 31.43562, 
    31.55631, 31.67694, 31.7975, 31.91799, 32.03841, 32.15877, 32.27906, 
    32.39928, 32.51943, 32.63951, 32.75953, 32.87947, 32.99934, 33.11914, 
    33.23886, 33.35852, 33.4781, 33.5976, 33.71704, 33.8364, 33.95568, 
    34.07489, 34.19402, 34.31308, 34.43206, 34.55096, 34.66978, 34.78853, 
    34.9072, 35.02579, 35.1443, 35.26273, 35.38108, 35.49936, 35.61754, 
    35.73565, 35.85368, 35.97162, 36.08948, 36.20726, 36.32495, 36.44257, 
    36.56009, 36.67754, 36.7949, 36.91217, 37.02935, 37.14645, 37.26347, 
    37.38039, 37.49723, 37.61398, 37.73064, 37.84722, 37.96371, 38.0801, 
    38.19641, 38.31263, 38.42876, 38.54479, 38.66074, 38.77659,
  -13.14912, -13.0427, -12.93618, -12.82954, -12.72279, -12.61593, -12.50896, 
    -12.40188, -12.29469, -12.18738, -12.07997, -11.97244, -11.86481, 
    -11.75706, -11.64921, -11.54124, -11.43317, -11.32498, -11.21668, 
    -11.10828, -10.99977, -10.89114, -10.78241, -10.67357, -10.56462, 
    -10.45556, -10.34639, -10.23711, -10.12773, -10.01823, -9.908632, 
    -9.798923, -9.689107, -9.579183, -9.469151, -9.359013, -9.248767, 
    -9.138414, -9.027956, -8.917391, -8.806719, -8.695941, -8.585058, 
    -8.474069, -8.362974, -8.251774, -8.14047, -8.029059, -7.917545, 
    -7.805926, -7.694203, -7.582376, -7.470445, -7.35841, -7.246273, 
    -7.134032, -7.021688, -6.909241, -6.796692, -6.684042, -6.571289, 
    -6.458434, -6.345478, -6.23242, -6.119262, -6.006003, -5.892644, 
    -5.779184, -5.665625, -5.551966, -5.438208, -5.32435, -5.210394, 
    -5.09634, -4.982187, -4.867936, -4.753587, -4.639141, -4.524598, 
    -4.409958, -4.295222, -4.180389, -4.065461, -3.950437, -3.835318, 
    -3.720104, -3.604795, -3.489392, -3.373895, -3.258304, -3.14262, 
    -3.026843, -2.910973, -2.795011, -2.678957, -2.562811, -2.446574, 
    -2.330246, -2.213827, -2.097319, -1.98072, -1.864031, -1.747254, 
    -1.630388, -1.513433, -1.39639, -1.27926, -1.162042, -1.044737, 
    -0.9273456, -0.8098681, -0.6923048, -0.5746561, -0.4569224, -0.3391041, 
    -0.2212016, -0.1032152, 0.0148545, 0.1330072, 0.2512425, 0.36956, 
    0.4879592, 0.6064398, 0.7250013, 0.8436432, 0.9623653, 1.081167, 
    1.200048, 1.319008, 1.438046, 1.557161, 1.676355, 1.795625, 1.914972, 
    2.034395, 2.153893, 2.273467, 2.393116, 2.512839, 2.632635, 2.752505, 
    2.872448, 2.992463, 3.11255, 3.232709, 3.352939, 3.473239, 3.593609, 
    3.714049, 3.834557, 3.955134, 4.07578, 4.196493, 4.317272, 4.438118, 
    4.559031, 4.680009, 4.801052, 4.922159, 5.043331, 5.164566, 5.285864, 
    5.407224, 5.528646, 5.65013, 5.771675, 5.89328, 6.014944, 6.136668, 
    6.258451, 6.380291, 6.50219, 6.624146, 6.746158, 6.868226, 6.99035, 
    7.112528, 7.234761, 7.357048, 7.479388, 7.601781, 7.724226, 7.846722, 
    7.96927, 8.091867, 8.214515, 8.337212, 8.459958, 8.582751, 8.705593, 
    8.828482, 8.951416, 9.074397, 9.197423, 9.320493, 9.443607, 9.566766, 
    9.689966, 9.81321, 9.936495, 10.05982, 10.18319, 10.30659, 10.43004, 
    10.55352, 10.67705, 10.80061, 10.9242, 11.04784, 11.1715, 11.29521, 
    11.41895, 11.54272, 11.66652, 11.79036, 11.91423, 12.03813, 12.16206, 
    12.28603, 12.41002, 12.53404, 12.65809, 12.78216, 12.90627, 13.0304, 
    13.15455, 13.27873, 13.40294, 13.52717, 13.65142, 13.77569, 13.89999, 
    14.02431, 14.14864, 14.273, 14.39738, 14.52178, 14.64619, 14.77062, 
    14.89507, 15.01954, 15.14402, 15.26851, 15.39302, 15.51754, 15.64208, 
    15.76663, 15.89119, 16.01576, 16.14034, 16.26493, 16.38953, 16.51414, 
    16.63876, 16.76338, 16.88801, 17.01264, 17.13729, 17.26193, 17.38658, 
    17.51123, 17.63589, 17.76054, 17.8852, 18.00986, 18.13452, 18.25918, 
    18.38383, 18.50849, 18.63314, 18.75779, 18.88243, 19.00707, 19.13171, 
    19.25633, 19.38096, 19.50557, 19.63018, 19.75478, 19.87937, 20.00395, 
    20.12852, 20.25307, 20.37762, 20.50216, 20.62668, 20.75118, 20.87568, 
    21.00015, 21.12462, 21.24906, 21.37349, 21.4979, 21.6223, 21.74667, 
    21.87103, 21.99536, 22.11967, 22.24397, 22.36824, 22.49249, 22.61671, 
    22.74091, 22.86509, 22.98924, 23.11337, 23.23746, 23.36154, 23.48558, 
    23.6096, 23.73358, 23.85754, 23.98147, 24.10536, 24.22923, 24.35306, 
    24.47686, 24.60063, 24.72436, 24.84806, 24.97172, 25.09535, 25.21894, 
    25.34249, 25.46601, 25.58949, 25.71293, 25.83633, 25.95969, 26.08301, 
    26.20629, 26.32952, 26.45272, 26.57587, 26.69898, 26.82204, 26.94506, 
    27.06803, 27.19096, 27.31384, 27.43668, 27.55946, 27.6822, 27.80489, 
    27.92753, 28.05012, 28.17266, 28.29515, 28.41758, 28.53997, 28.6623, 
    28.78458, 28.9068, 29.02897, 29.15109, 29.27315, 29.39515, 29.5171, 
    29.63899, 29.76082, 29.88259, 30.0043, 30.12596, 30.24756, 30.36909, 
    30.49056, 30.61198, 30.73333, 30.85462, 30.97584, 31.097, 31.2181, 
    31.33913, 31.4601, 31.581, 31.70184, 31.82261, 31.94331, 32.06394, 
    32.18451, 32.30501, 32.42544, 32.5458, 32.66608, 32.7863, 32.90645, 
    33.02653, 33.14653, 33.26646, 33.38632, 33.5061, 33.62582, 33.74545, 
    33.86501, 33.9845, 34.10391, 34.22325, 34.34251, 34.46169, 34.58079, 
    34.69981, 34.81876, 34.93763, 35.05642, 35.17513, 35.29376, 35.41231, 
    35.53078, 35.64916, 35.76747, 35.88569, 36.00383, 36.12188, 36.23986, 
    36.35775, 36.47555, 36.59327, 36.71091, 36.82846, 36.94592, 37.0633, 
    37.18059, 37.29779, 37.41491, 37.53194, 37.64888, 37.76573, 37.8825, 
    37.99917, 38.11575, 38.23225, 38.34865, 38.46497, 38.58119, 38.69732, 
    38.81336,
  -13.20101, -13.09446, -12.98779, -12.88101, -12.77412, -12.66712, 
    -12.56001, -12.45279, -12.34545, -12.238, -12.13045, -12.02278, -11.915, 
    -11.80711, -11.69911, -11.59099, -11.48277, -11.37444, -11.266, 
    -11.15744, -11.04878, -10.94001, -10.83112, -10.72213, -10.61303, 
    -10.50382, -10.3945, -10.28507, -10.17553, -10.06589, -9.956132, 
    -9.846269, -9.736298, -9.626218, -9.516031, -9.405736, -9.295334, 
    -9.184825, -9.074208, -8.963485, -8.852654, -8.741717, -8.630674, 
    -8.519525, -8.40827, -8.296908, -8.185442, -8.07387, -7.962193, 
    -7.850411, -7.738524, -7.626533, -7.514437, -7.402237, -7.289934, 
    -7.177527, -7.065017, -6.952403, -6.839686, -6.726867, -6.613945, 
    -6.500922, -6.387796, -6.274569, -6.16124, -6.04781, -5.934279, 
    -5.820647, -5.706915, -5.593083, -5.479152, -5.36512, -5.250989, 
    -5.13676, -5.022431, -4.908004, -4.793479, -4.678856, -4.564136, 
    -4.449318, -4.334403, -4.219392, -4.104284, -3.98908, -3.87378, 
    -3.758385, -3.642895, -3.52731, -3.411631, -3.295857, -3.17999, 
    -3.064029, -2.947975, -2.831829, -2.715589, -2.599258, -2.482835, 
    -2.36632, -2.249715, -2.133018, -2.016232, -1.899355, -1.782388, 
    -1.665333, -1.548188, -1.430955, -1.313634, -1.196225, -1.078729, 
    -0.9611452, -0.8434752, -0.7257189, -0.6078768, -0.4899493, -0.3719366, 
    -0.2538394, -0.1356578, -0.01739248, 0.1009563, 0.2193881, 0.3379025, 
    0.4564992, 0.5751776, 0.6939372, 0.8127779, 0.931699, 1.0507, 1.169781, 
    1.288941, 1.40818, 1.527497, 1.646892, 1.766364, 1.885913, 2.005539, 
    2.125241, 2.245019, 2.364872, 2.484799, 2.6048, 2.724875, 2.845024, 
    2.965245, 3.085539, 3.205904, 3.326341, 3.446849, 3.567427, 3.688075, 
    3.808793, 3.929579, 4.050434, 4.171356, 4.292346, 4.413403, 4.534526, 
    4.655716, 4.77697, 4.89829, 5.019674, 5.141121, 5.262632, 5.384206, 
    5.505843, 5.62754, 5.749299, 5.871119, 5.992999, 6.114938, 6.236937, 
    6.358994, 6.481109, 6.603281, 6.72551, 6.847796, 6.970137, 7.092534, 
    7.214985, 7.337491, 7.46005, 7.582662, 7.705326, 7.828042, 7.950809, 
    8.073627, 8.196496, 8.319414, 8.442381, 8.565396, 8.688459, 8.81157, 
    8.934727, 9.05793, 9.181179, 9.304472, 9.42781, 9.551191, 9.674617, 
    9.798083, 9.921593, 10.04514, 10.16873, 10.29237, 10.41604, 10.53975, 
    10.66349, 10.78728, 10.9111, 11.03496, 11.15886, 11.28279, 11.40675, 
    11.53075, 11.65479, 11.77885, 11.90295, 12.02708, 12.15124, 12.27543, 
    12.39965, 12.5239, 12.64817, 12.77248, 12.89681, 13.02117, 13.14555, 
    13.26996, 13.3944, 13.51886, 13.64334, 13.76784, 13.89237, 14.01692, 
    14.14148, 14.26607, 14.39068, 14.51531, 14.63995, 14.76462, 14.88929, 
    15.01399, 15.1387, 15.26343, 15.38817, 15.51292, 15.63769, 15.76247, 
    15.88726, 16.01206, 16.13688, 16.2617, 16.38653, 16.51137, 16.63622, 
    16.76108, 16.88594, 17.01081, 17.13568, 17.26056, 17.38544, 17.51032, 
    17.63521, 17.7601, 17.88499, 18.00988, 18.13477, 18.25966, 18.38455, 
    18.50943, 18.63432, 18.7592, 18.88408, 19.00895, 19.13381, 19.25867, 
    19.38353, 19.50838, 19.63321, 19.75805, 19.88287, 20.00768, 20.13248, 
    20.25727, 20.38205, 20.50681, 20.63156, 20.7563, 20.88103, 21.00574, 
    21.13043, 21.25511, 21.37977, 21.50441, 21.62903, 21.75364, 21.87822, 
    22.00279, 22.12733, 22.25186, 22.37636, 22.50083, 22.62529, 22.74972, 
    22.87412, 22.9985, 23.12286, 23.24719, 23.37149, 23.49576, 23.62, 
    23.74422, 23.86841, 23.99256, 24.11668, 24.24078, 24.36484, 24.48886, 
    24.61286, 24.73682, 24.86074, 24.98463, 25.10849, 25.2323, 25.35608, 
    25.47983, 25.60353, 25.72719, 25.85082, 25.9744, 26.09795, 26.22145, 
    26.34491, 26.46833, 26.5917, 26.71503, 26.83832, 26.96156, 27.08476, 
    27.20791, 27.33101, 27.45407, 27.57707, 27.70003, 27.82294, 27.9458, 
    28.06861, 28.19137, 28.31408, 28.43674, 28.55934, 28.68189, 28.80439, 
    28.92683, 29.04922, 29.17155, 29.29383, 29.41605, 29.53821, 29.66032, 
    29.78237, 29.90435, 30.02629, 30.14816, 30.26997, 30.39171, 30.5134, 
    30.63503, 30.75659, 30.87809, 30.99953, 31.1209, 31.24221, 31.36346, 
    31.48464, 31.60575, 31.7268, 31.84778, 31.96869, 32.08953, 32.21031, 
    32.33101, 32.45165, 32.57222, 32.69271, 32.81314, 32.93349, 33.05378, 
    33.17399, 33.29412, 33.41419, 33.53418, 33.65409, 33.77393, 33.8937, 
    34.01339, 34.133, 34.25254, 34.372, 34.49138, 34.61069, 34.72991, 
    34.84906, 34.96813, 35.08712, 35.20603, 35.32486, 35.4436, 35.56227, 
    35.68085, 35.79935, 35.91777, 36.03611, 36.15436, 36.27253, 36.39061, 
    36.50861, 36.62652, 36.74435, 36.86209, 36.97975, 37.09732, 37.2148, 
    37.3322, 37.4495, 37.56672, 37.68386, 37.8009, 37.91785, 38.03471, 
    38.15149, 38.26817, 38.38476, 38.50126, 38.61766, 38.73398, 38.85021,
  -13.253, -13.1463, -13.0395, -12.93258, -12.82555, -12.71841, -12.61115, 
    -12.50379, -12.39631, -12.28872, -12.18102, -12.0732, -11.96528, 
    -11.85724, -11.7491, -11.64084, -11.53247, -11.42399, -11.3154, -11.2067, 
    -11.09788, -10.98896, -10.87993, -10.77079, -10.66154, -10.55217, 
    -10.4427, -10.33312, -10.22343, -10.11363, -10.00372, -9.893704, 
    -9.783578, -9.673344, -9.563001, -9.45255, -9.341991, -9.231324, 
    -9.12055, -9.009668, -8.898679, -8.787583, -8.67638, -8.56507, -8.453654, 
    -8.342132, -8.230503, -8.118769, -8.006929, -7.894984, -7.782933, 
    -7.670778, -7.558517, -7.446152, -7.333683, -7.22111, -7.108432, 
    -6.995651, -6.882767, -6.76978, -6.656689, -6.543496, -6.430201, 
    -6.316803, -6.203303, -6.089702, -5.975999, -5.862195, -5.748291, 
    -5.634285, -5.52018, -5.405974, -5.291668, -5.177264, -5.062759, 
    -4.948156, -4.833455, -4.718654, -4.603756, -4.48876, -4.373667, 
    -4.258476, -4.143188, -4.027805, -3.912324, -3.796748, -3.681077, 
    -3.56531, -3.449448, -3.333491, -3.21744, -3.101295, -2.985057, 
    -2.868726, -2.752301, -2.635784, -2.519174, -2.402473, -2.28568, 
    -2.168796, -2.051821, -1.934755, -1.8176, -1.700355, -1.58302, -1.465596, 
    -1.348084, -1.230484, -1.112795, -0.9950196, -0.8771567, -0.7592071, 
    -0.6411713, -0.5230496, -0.4048423, -0.28655, -0.1681729, -0.04971161, 
    0.06883359, 0.1874623, 0.306174, 0.4249683, 0.5438448, 0.6628031, 
    0.7818428, 0.9009634, 1.020164, 1.139446, 1.258806, 1.378246, 1.497765, 
    1.617362, 1.737037, 1.856789, 1.976618, 2.096523, 2.216505, 2.336562, 
    2.456694, 2.576901, 2.697182, 2.817537, 2.937964, 3.058465, 3.179038, 
    3.299682, 3.420398, 3.541184, 3.662041, 3.782968, 3.903964, 4.025028, 
    4.146161, 4.267362, 4.38863, 4.509964, 4.631366, 4.752832, 4.874364, 
    4.995961, 5.117622, 5.239347, 5.361135, 5.482985, 5.604897, 5.726871, 
    5.848906, 5.971001, 6.093157, 6.215372, 6.337645, 6.459977, 6.582366, 
    6.704813, 6.827317, 6.949876, 7.072492, 7.195162, 7.317886, 7.440664, 
    7.563496, 7.68638, 7.809317, 7.932305, 8.055344, 8.178433, 8.301573, 
    8.424762, 8.547998, 8.671285, 8.794618, 8.917997, 9.041423, 9.164895, 
    9.288412, 9.411974, 9.53558, 9.659228, 9.782921, 9.906654, 10.03043, 
    10.15425, 10.2781, 10.402, 10.52594, 10.64991, 10.77392, 10.89797, 
    11.02206, 11.14618, 11.27034, 11.39453, 11.51876, 11.64302, 11.76731, 
    11.89164, 12.01599, 12.14038, 12.2648, 12.38925, 12.51373, 12.63823, 
    12.76277, 12.88733, 13.01192, 13.13653, 13.26117, 13.38584, 13.51052, 
    13.63524, 13.75997, 13.88473, 14.00951, 14.13431, 14.25913, 14.38396, 
    14.50882, 14.6337, 14.75859, 14.8835, 15.00843, 15.13338, 15.25833, 
    15.38331, 15.50829, 15.63329, 15.7583, 15.88333, 16.00836, 16.13341, 
    16.25846, 16.38353, 16.5086, 16.63368, 16.75877, 16.88386, 17.00896, 
    17.13407, 17.25918, 17.38429, 17.50941, 17.63453, 17.75965, 17.88477, 
    18.0099, 18.13502, 18.26014, 18.38526, 18.51038, 18.6355, 18.76061, 
    18.88572, 19.01083, 19.13593, 19.26102, 19.38611, 19.51119, 19.63626, 
    19.76132, 19.88637, 20.01142, 20.13645, 20.26147, 20.38648, 20.51148, 
    20.63646, 20.76143, 20.88639, 21.01133, 21.13626, 21.26116, 21.38605, 
    21.51093, 21.63578, 21.76062, 21.88544, 22.01023, 22.13501, 22.25976, 
    22.38449, 22.5092, 22.63389, 22.75855, 22.88318, 23.00779, 23.13238, 
    23.25693, 23.38146, 23.50597, 23.63044, 23.75488, 23.8793, 24.00368, 
    24.12803, 24.25235, 24.37664, 24.5009, 24.62512, 24.74931, 24.87346, 
    24.99757, 25.12165, 25.2457, 25.3697, 25.49367, 25.6176, 25.74149, 
    25.86534, 25.98915, 26.11292, 26.23665, 26.36033, 26.48398, 26.60757, 
    26.73113, 26.85464, 26.9781, 27.10152, 27.2249, 27.34822, 27.4715, 
    27.59473, 27.71791, 27.84104, 27.96412, 28.08715, 28.21013, 28.33306, 
    28.45594, 28.57876, 28.70153, 28.82425, 28.94691, 29.06952, 29.19206, 
    29.31456, 29.437, 29.55938, 29.6817, 29.80396, 29.92617, 30.04832, 
    30.1704, 30.29243, 30.41439, 30.53629, 30.65813, 30.77991, 30.90163, 
    31.02328, 31.14487, 31.26639, 31.38784, 31.50923, 31.63056, 31.75181, 
    31.873, 31.99413, 32.11518, 32.23616, 32.35708, 32.47793, 32.5987, 
    32.71941, 32.84004, 32.9606, 33.08109, 33.20151, 33.32185, 33.44212, 
    33.56231, 33.68243, 33.80248, 33.92245, 34.04234, 34.16216, 34.2819, 
    34.40156, 34.52114, 34.64065, 34.76008, 34.87943, 34.9987, 35.11789, 
    35.23699, 35.35602, 35.47496, 35.59383, 35.71261, 35.83131, 35.94992, 
    36.06845, 36.1869, 36.30527, 36.42355, 36.54174, 36.65985, 36.77787, 
    36.89581, 37.01366, 37.13142, 37.24909, 37.36668, 37.48418, 37.60159, 
    37.71891, 37.83614, 37.95328, 38.07033, 38.18729, 38.30416, 38.42094, 
    38.53762, 38.65422, 38.77073, 38.88713,
  -13.30508, -13.19824, -13.0913, -12.98424, -12.87707, -12.76978, -12.66239, 
    -12.55488, -12.44726, -12.33953, -12.23168, -12.12372, -12.01565, 
    -11.90747, -11.79918, -11.69077, -11.58226, -11.47363, -11.36489, 
    -11.25604, -11.14708, -11.03801, -10.92883, -10.81953, -10.71013, 
    -10.60062, -10.49099, -10.38126, -10.27142, -10.16146, -10.0514, 
    -9.941231, -9.83095, -9.72056, -9.610061, -9.499454, -9.388738, 
    -9.277914, -9.166982, -9.055942, -8.944794, -8.833538, -8.722175, 
    -8.610705, -8.499128, -8.387444, -8.275654, -8.163757, -8.051754, 
    -7.939645, -7.827431, -7.715111, -7.602685, -7.490155, -7.37752, 
    -7.26478, -7.151936, -7.038988, -6.925935, -6.812779, -6.69952, 
    -6.586157, -6.472692, -6.359124, -6.245453, -6.13168, -6.017806, 
    -5.903829, -5.789752, -5.675573, -5.561293, -5.446913, -5.332433, 
    -5.217852, -5.103172, -4.988392, -4.873514, -4.758536, -4.64346, 
    -4.528286, -4.413013, -4.297643, -4.182176, -4.066612, -3.950951, 
    -3.835193, -3.71934, -3.60339, -3.487345, -3.371206, -3.254971, 
    -3.138642, -3.022219, -2.905702, -2.789092, -2.672389, -2.555592, 
    -2.438704, -2.321723, -2.204651, -2.087488, -1.970233, -1.852888, 
    -1.735453, -1.617928, -1.500314, -1.38261, -1.264818, -1.146937, 
    -1.028969, -0.9109131, -0.7927699, -0.67454, -0.5562238, -0.4378216, 
    -0.3193339, -0.200761, -0.08210333, 0.0366386, 0.1554644, 0.2743738, 
    0.3933662, 0.5124412, 0.6315985, 0.7508375, 0.8701579, 0.9895592, 
    1.109041, 1.228603, 1.348244, 1.467965, 1.587764, 1.707642, 1.827597, 
    1.94763, 2.067739, 2.187925, 2.308187, 2.428525, 2.548937, 2.669424, 
    2.789985, 2.91062, 3.031327, 3.152108, 3.27296, 3.393885, 3.51488, 
    3.635946, 3.757082, 3.878288, 3.999563, 4.120907, 4.242319, 4.363798, 
    4.485345, 4.606958, 4.728637, 4.850382, 4.972192, 5.094067, 5.216005, 
    5.338007, 5.460073, 5.5822, 5.704389, 5.82664, 5.948951, 6.071323, 
    6.193755, 6.316245, 6.438795, 6.561402, 6.684067, 6.806788, 6.929567, 
    7.052401, 7.17529, 7.298234, 7.421233, 7.544284, 7.667389, 7.790546, 
    7.913755, 8.037016, 8.160327, 8.283689, 8.4071, 8.53056, 8.654067, 
    8.777623, 8.901226, 9.024877, 9.148572, 9.272313, 9.396099, 9.519929, 
    9.643804, 9.76772, 9.891679, 10.01568, 10.13972, 10.26381, 10.38793, 
    10.51209, 10.63629, 10.76053, 10.88481, 11.00912, 11.13347, 11.25786, 
    11.38228, 11.50673, 11.63122, 11.75574, 11.8803, 12.00488, 12.1295, 
    12.25415, 12.37883, 12.50353, 12.62827, 12.75303, 12.87782, 13.00264, 
    13.12749, 13.25236, 13.37725, 13.50217, 13.62712, 13.75208, 13.87707, 
    14.00208, 14.12711, 14.25216, 14.37723, 14.50232, 14.62743, 14.75256, 
    14.8777, 15.00286, 15.12803, 15.25323, 15.37843, 15.50365, 15.62888, 
    15.75413, 15.87938, 16.00465, 16.12993, 16.25522, 16.38051, 16.50582, 
    16.63113, 16.75645, 16.88178, 17.00711, 17.13245, 17.2578, 17.38314, 
    17.50849, 17.63385, 17.7592, 17.88456, 18.00991, 18.13527, 18.26063, 
    18.38598, 18.51134, 18.63668, 18.76203, 18.88737, 19.01271, 19.13804, 
    19.26337, 19.38869, 19.514, 19.63931, 19.7646, 19.88989, 20.01517, 
    20.14043, 20.26569, 20.39093, 20.51616, 20.64138, 20.76658, 20.89177, 
    21.01694, 21.1421, 21.26724, 21.39236, 21.51747, 21.64255, 21.76762, 
    21.89267, 22.0177, 22.1427, 22.26769, 22.39265, 22.51759, 22.64251, 
    22.7674, 22.89226, 23.0171, 23.14192, 23.2667, 23.39146, 23.5162, 
    23.6409, 23.76557, 23.89021, 24.01483, 24.13941, 24.26396, 24.38848, 
    24.51296, 24.63741, 24.76182, 24.8862, 25.01055, 25.13485, 25.25912, 
    25.38336, 25.50755, 25.63171, 25.75583, 25.8799, 26.00394, 26.12793, 
    26.25188, 26.3758, 26.49966, 26.62349, 26.74726, 26.871, 26.99469, 
    27.11833, 27.24192, 27.36547, 27.48897, 27.61242, 27.73583, 27.85918, 
    27.98248, 28.10574, 28.22894, 28.35209, 28.47518, 28.59823, 28.72122, 
    28.84415, 28.96703, 29.08986, 29.21263, 29.33534, 29.458, 29.5806, 
    29.70313, 29.82562, 29.94804, 30.0704, 30.1927, 30.31494, 30.43712, 
    30.55924, 30.6813, 30.80329, 30.92522, 31.04708, 31.16888, 31.29062, 
    31.41228, 31.53389, 31.65542, 31.77689, 31.89829, 32.01963, 32.14089, 
    32.26208, 32.38321, 32.50426, 32.62525, 32.74616, 32.867, 32.98777, 
    33.10847, 33.22909, 33.34964, 33.47012, 33.59052, 33.71084, 33.83109, 
    33.95126, 34.07136, 34.19138, 34.31133, 34.43119, 34.55098, 34.67068, 
    34.79031, 34.90987, 35.02934, 35.14872, 35.26803, 35.38726, 35.5064, 
    35.62546, 35.74444, 35.86334, 35.98215, 36.10088, 36.21952, 36.33808, 
    36.45656, 36.57494, 36.69325, 36.81146, 36.92959, 37.04763, 37.16559, 
    37.28346, 37.40123, 37.51892, 37.63652, 37.75404, 37.87146, 37.98879, 
    38.10603, 38.22318, 38.34023, 38.4572, 38.57407, 38.69086, 38.80754, 
    38.92414,
  -13.35725, -13.25028, -13.14319, -13.03599, -12.92868, -12.82125, 
    -12.71372, -12.60606, -12.4983, -12.39042, -12.28244, -12.17433, 
    -12.06612, -11.95779, -11.84935, -11.7408, -11.63214, -11.52336, 
    -11.41448, -11.30548, -11.19637, -11.08715, -10.97782, -10.86837, 
    -10.75882, -10.64915, -10.53938, -10.42949, -10.3195, -10.20939, 
    -10.09917, -9.988849, -9.878412, -9.767867, -9.657212, -9.546449, 
    -9.435575, -9.324594, -9.213504, -9.102305, -8.990998, -8.879583, 
    -8.76806, -8.656429, -8.544692, -8.432846, -8.320894, -8.208835, 
    -8.096668, -7.984396, -7.872018, -7.759533, -7.646943, -7.534246, 
    -7.421445, -7.308539, -7.195528, -7.082411, -6.969191, -6.855866, 
    -6.742438, -6.628906, -6.51527, -6.401531, -6.287689, -6.173745, 
    -6.059698, -5.945549, -5.831298, -5.716946, -5.602492, -5.487937, 
    -5.373281, -5.258525, -5.143669, -5.028713, -4.913657, -4.798502, 
    -4.683248, -4.567894, -4.452443, -4.336894, -4.221246, -4.105501, 
    -3.989659, -3.87372, -3.757684, -3.641553, -3.525325, -3.409002, 
    -3.292583, -3.176069, -3.059461, -2.942759, -2.825963, -2.709073, 
    -2.59209, -2.475014, -2.357846, -2.240585, -2.123233, -2.00579, 
    -1.888255, -1.770629, -1.652914, -1.535108, -1.417213, -1.299229, 
    -1.181156, -1.062994, -0.9447448, -0.8264077, -0.7079835, -0.5894724, 
    -0.4708749, -0.3521914, -0.2334224, -0.1145681, 0.004370888, 0.1233943, 
    0.2425016, 0.3616924, 0.4809662, 0.6003228, 0.7197616, 0.8392821, 
    0.958884, 1.078567, 1.19833, 1.318174, 1.438096, 1.558098, 1.678179, 
    1.798338, 1.918575, 2.038889, 2.15928, 2.279747, 2.40029, 2.520908, 
    2.641602, 2.76237, 2.883212, 3.004127, 3.125115, 3.246176, 3.36731, 
    3.488514, 3.60979, 3.731136, 3.852552, 3.974038, 4.095593, 4.217216, 
    4.338908, 4.460666, 4.582492, 4.704385, 4.826343, 4.948367, 5.070456, 
    5.192608, 5.314825, 5.437105, 5.559448, 5.681853, 5.80432, 5.926848, 
    6.049437, 6.172086, 6.294794, 6.417561, 6.540387, 6.66327, 6.786211, 
    6.909208, 7.032261, 7.155371, 7.278535, 7.401753, 7.525026, 7.648352, 
    7.77173, 7.895161, 8.018643, 8.142177, 8.26576, 8.389394, 8.513077, 
    8.636808, 8.760588, 8.884415, 9.008288, 9.132209, 9.256174, 9.380185, 
    9.504241, 9.62834, 9.752482, 9.876667, 10.00089, 10.12516, 10.24947, 
    10.37382, 10.49821, 10.62264, 10.74711, 10.87161, 10.99615, 11.12073, 
    11.24534, 11.36999, 11.49468, 11.61939, 11.74414, 11.86893, 11.99374, 
    12.11859, 12.24347, 12.36838, 12.49331, 12.61828, 12.74327, 12.8683, 
    12.99335, 13.11842, 13.24352, 13.36865, 13.4938, 13.61897, 13.74417, 
    13.86939, 13.99463, 14.1199, 14.24518, 14.37048, 14.4958, 14.62115, 
    14.7465, 14.87188, 14.99727, 15.12268, 15.24811, 15.37354, 15.49899, 
    15.62446, 15.74994, 15.87543, 16.00093, 16.12644, 16.25196, 16.37749, 
    16.50303, 16.62858, 16.75413, 16.87969, 17.00526, 17.13083, 17.25641, 
    17.38199, 17.50758, 17.63316, 17.75875, 17.88434, 18.00993, 18.13552, 
    18.26111, 18.3867, 18.51229, 18.63787, 18.76345, 18.88903, 19.0146, 
    19.14017, 19.26573, 19.39128, 19.51683, 19.64236, 19.76789, 19.89342, 
    20.01892, 20.14442, 20.26991, 20.39539, 20.52085, 20.6463, 20.77174, 
    20.89716, 21.02256, 21.14795, 21.27333, 21.39868, 21.52402, 21.64934, 
    21.77464, 21.89992, 22.02518, 22.15042, 22.27563, 22.40083, 22.526, 
    22.65115, 22.77627, 22.90137, 23.02644, 23.15148, 23.2765, 23.40149, 
    23.52645, 23.65138, 23.77629, 23.90116, 24.026, 24.15081, 24.27559, 
    24.40034, 24.52505, 24.64973, 24.77437, 24.89898, 25.02355, 25.14809, 
    25.27258, 25.39705, 25.52147, 25.64585, 25.7702, 25.8945, 26.01876, 
    26.14298, 26.26716, 26.39129, 26.51539, 26.63943, 26.76344, 26.8874, 
    27.01131, 27.13518, 27.259, 27.38277, 27.50649, 27.63017, 27.75379, 
    27.87737, 28.00089, 28.12437, 28.24779, 28.37116, 28.49448, 28.61774, 
    28.74095, 28.86411, 28.98721, 29.11025, 29.23324, 29.35617, 29.47905, 
    29.60186, 29.72462, 29.84732, 29.96996, 30.09254, 30.21506, 30.33751, 
    30.45991, 30.58224, 30.70451, 30.82672, 30.94886, 31.07094, 31.19295, 
    31.3149, 31.43678, 31.5586, 31.68035, 31.80203, 31.92364, 32.04519, 
    32.16666, 32.28806, 32.4094, 32.53066, 32.65186, 32.77298, 32.89403, 
    33.015, 33.13591, 33.25674, 33.37749, 33.49818, 33.61878, 33.73932, 
    33.85977, 33.98015, 34.10045, 34.22067, 34.34082, 34.46089, 34.58088, 
    34.70079, 34.82062, 34.94037, 35.06004, 35.17963, 35.29914, 35.41856, 
    35.53791, 35.65717, 35.77634, 35.89544, 36.01445, 36.13337, 36.25222, 
    36.37097, 36.48964, 36.60822, 36.72672, 36.84513, 36.96346, 37.08169, 
    37.19984, 37.3179, 37.43587, 37.55375, 37.67154, 37.78924, 37.90685, 
    38.02437, 38.1418, 38.25914, 38.37638, 38.49354, 38.6106, 38.72757, 
    38.84444, 38.96123,
  -13.40951, -13.3024, -13.19518, -13.08784, -12.98038, -12.87282, -12.76514, 
    -12.65734, -12.54944, -12.44142, -12.33328, -12.22504, -12.11668, 
    -12.00821, -11.89962, -11.79092, -11.68211, -11.57319, -11.46416, 
    -11.35501, -11.24575, -11.13638, -11.0269, -10.9173, -10.8076, -10.69778, 
    -10.58786, -10.47782, -10.36767, -10.25741, -10.14704, -10.03656, 
    -9.925966, -9.815266, -9.704455, -9.593534, -9.482505, -9.371366, 
    -9.260117, -9.14876, -9.037293, -8.925719, -8.814036, -8.702245, 
    -8.590345, -8.478338, -8.366224, -8.254002, -8.141673, -8.029237, 
    -7.916694, -7.804045, -7.691289, -7.578427, -7.465459, -7.352386, 
    -7.239208, -7.125924, -7.012535, -6.899042, -6.785444, -6.671742, 
    -6.557936, -6.444026, -6.330013, -6.215897, -6.101678, -5.987356, 
    -5.872932, -5.758405, -5.643777, -5.529047, -5.414217, -5.299284, 
    -5.184252, -5.069119, -4.953886, -4.838552, -4.72312, -4.607588, 
    -4.491957, -4.376228, -4.2604, -4.144475, -4.028451, -3.91233, -3.796112, 
    -3.679797, -3.563386, -3.446879, -3.330276, -3.213578, -3.096785, 
    -2.979897, -2.862914, -2.745838, -2.628668, -2.511404, -2.394048, 
    -2.276599, -2.159057, -2.041424, -1.923699, -1.805884, -1.687977, 
    -1.56998, -1.451893, -1.333716, -1.21545, -1.097096, -0.9786524, 
    -0.8601211, -0.7415021, -0.6227959, -0.5040028, -0.3851233, -0.2661577, 
    -0.1471065, -0.02797002, 0.09125121, 0.2105568, 0.3299464, 0.4494195, 
    0.5689757, 0.6886145, 0.8083356, 0.9281384, 1.048023, 1.167988, 1.288033, 
    1.408159, 1.528364, 1.648648, 1.769011, 1.889452, 2.009971, 2.130567, 
    2.25124, 2.371989, 2.492814, 2.613714, 2.734689, 2.855739, 2.976863, 
    3.09806, 3.219329, 3.340672, 3.462086, 3.583572, 3.705128, 3.826755, 
    3.948452, 4.070219, 4.192054, 4.313958, 4.435929, 4.557969, 4.680074, 
    4.802247, 4.924484, 5.046788, 5.169156, 5.291587, 5.414083, 5.536642, 
    5.659264, 5.781947, 5.904692, 6.027498, 6.150364, 6.273291, 6.396276, 
    6.51932, 6.642423, 6.765583, 6.8888, 7.012074, 7.135403, 7.258788, 
    7.382227, 7.505721, 7.629268, 7.752868, 7.876521, 8.000226, 8.123981, 
    8.247788, 8.371645, 8.495551, 8.619507, 8.74351, 8.867561, 8.99166, 
    9.115805, 9.239996, 9.364232, 9.488513, 9.612838, 9.737206, 9.861618, 
    9.986072, 10.11057, 10.2351, 10.35968, 10.4843, 10.60895, 10.73365, 
    10.85838, 10.98315, 11.10796, 11.2328, 11.35768, 11.48259, 11.60754, 
    11.73252, 11.85753, 11.98258, 12.10765, 12.23276, 12.3579, 12.48307, 
    12.60827, 12.73349, 12.85875, 12.98403, 13.10933, 13.23467, 13.36002, 
    13.48541, 13.61081, 13.73624, 13.8617, 13.98717, 14.11266, 14.23818, 
    14.36372, 14.48927, 14.61485, 14.74044, 14.86605, 14.99167, 15.11731, 
    15.24297, 15.36864, 15.49433, 15.62003, 15.74574, 15.87146, 15.9972, 
    16.12294, 16.2487, 16.37446, 16.50024, 16.62602, 16.75181, 16.8776, 
    17.0034, 17.12921, 17.25502, 17.38084, 17.50666, 17.63248, 17.7583, 
    17.88413, 18.00995, 18.13578, 18.2616, 18.38742, 18.51324, 18.63906, 
    18.76488, 18.89069, 19.01649, 19.1423, 19.26809, 19.39388, 19.51966, 
    19.64543, 19.77119, 19.89695, 20.02269, 20.14843, 20.27415, 20.39986, 
    20.52555, 20.65124, 20.77691, 20.90256, 21.0282, 21.15382, 21.27943, 
    21.40502, 21.53059, 21.65614, 21.78168, 21.90719, 22.03268, 22.15815, 
    22.2836, 22.40903, 22.53443, 22.65981, 22.78516, 22.91049, 23.03579, 
    23.16107, 23.28632, 23.41154, 23.53673, 23.6619, 23.78703, 23.91213, 
    24.03721, 24.16225, 24.28725, 24.41223, 24.53717, 24.66208, 24.78695, 
    24.91179, 25.03659, 25.16135, 25.28608, 25.41077, 25.53542, 25.66003, 
    25.7846, 25.90913, 26.03362, 26.15806, 26.28247, 26.40683, 26.53115, 
    26.65542, 26.77965, 26.90384, 27.02797, 27.15207, 27.27611, 27.4001, 
    27.52405, 27.64795, 27.7718, 27.8956, 28.01935, 28.14304, 28.26669, 
    28.39028, 28.51382, 28.6373, 28.76073, 28.88411, 29.00743, 29.1307, 
    29.2539, 29.37705, 29.50015, 29.62318, 29.74616, 29.86908, 29.99193, 
    30.11473, 30.23746, 30.36014, 30.48275, 30.6053, 30.72778, 30.85021, 
    30.97256, 31.09486, 31.21708, 31.33924, 31.46134, 31.58337, 31.70533, 
    31.82722, 31.94905, 32.0708, 32.19249, 32.31411, 32.43565, 32.55713, 
    32.67853, 32.79986, 32.92112, 33.0423, 33.16341, 33.28445, 33.40541, 
    33.5263, 33.64712, 33.76785, 33.88852, 34.0091, 34.1296, 34.25003, 
    34.37038, 34.49065, 34.61085, 34.73096, 34.85099, 34.97095, 35.09082, 
    35.21061, 35.33031, 35.44994, 35.56948, 35.68895, 35.80832, 35.92761, 
    36.04682, 36.16594, 36.28498, 36.40393, 36.5228, 36.64158, 36.76027, 
    36.87888, 36.99739, 37.11582, 37.23417, 37.35242, 37.47058, 37.58865, 
    37.70663, 37.82453, 37.94233, 38.06004, 38.17766, 38.29519, 38.41262, 
    38.52996, 38.64721, 38.76436, 38.88142, 38.99839,
  -13.46187, -13.35462, -13.24725, -13.13978, -13.03218, -12.92447, 
    -12.81665, -12.70872, -12.60067, -12.4925, -12.38422, -12.27583, 
    -12.16733, -12.05871, -11.94998, -11.84114, -11.73218, -11.62311, 
    -11.51393, -11.40463, -11.29523, -11.18571, -11.07607, -10.96633, 
    -10.85647, -10.7465, -10.63643, -10.52623, -10.41593, -10.30552, 
    -10.19499, -10.08436, -9.973613, -9.862757, -9.75179, -9.640713, 
    -9.529526, -9.418228, -9.306822, -9.195306, -9.08368, -8.971946, 
    -8.860103, -8.748151, -8.63609, -8.523922, -8.411645, -8.29926, 
    -8.186768, -8.074167, -7.96146, -7.848646, -7.735725, -7.622697, 
    -7.509563, -7.396323, -7.282977, -7.169525, -7.055968, -6.942306, 
    -6.828538, -6.714666, -6.60069, -6.486609, -6.372425, -6.258136, 
    -6.143745, -6.02925, -5.914652, -5.799952, -5.685149, -5.570244, 
    -5.455238, -5.34013, -5.224921, -5.109611, -4.9942, -4.878688, -4.763077, 
    -4.647366, -4.531556, -4.415647, -4.299638, -4.183531, -4.067326, 
    -3.951023, -3.834623, -3.718125, -3.601531, -3.484839, -3.368052, 
    -3.251169, -3.13419, -3.017116, -2.899947, -2.782684, -2.665326, 
    -2.547874, -2.43033, -2.312692, -2.194961, -2.077138, -1.959223, 
    -1.841216, -1.723118, -1.60493, -1.48665, -1.368281, -1.249822, 
    -1.131274, -1.012636, -0.8939103, -0.7750964, -0.6561947, -0.5372057, 
    -0.4181297, -0.2989673, -0.1797188, -0.06038459, 0.05903485, 0.1785391, 
    0.2981278, 0.4178004, 0.5375566, 0.6573959, 0.7773179, 0.8973221, 
    1.017408, 1.137575, 1.257824, 1.378152, 1.498561, 1.619049, 1.739616, 
    1.860262, 1.980986, 2.101788, 2.222667, 2.343622, 2.464654, 2.585762, 
    2.706944, 2.828202, 2.949534, 3.07094, 3.192419, 3.313971, 3.435595, 
    3.557292, 3.679059, 3.800897, 3.922806, 4.044785, 4.166832, 4.288949, 
    4.411133, 4.533386, 4.655705, 4.778092, 4.900545, 5.023063, 5.145646, 
    5.268294, 5.391006, 5.513781, 5.63662, 5.75952, 5.882483, 6.005507, 
    6.128591, 6.251736, 6.37494, 6.498203, 6.621525, 6.744905, 6.868342, 
    6.991836, 7.115386, 7.238992, 7.362653, 7.486368, 7.610137, 7.73396, 
    7.857835, 7.981763, 8.105742, 8.229773, 8.353853, 8.477983, 8.602162, 
    8.726391, 8.850667, 8.974991, 9.09936, 9.223778, 9.34824, 9.472747, 
    9.597299, 9.721893, 9.846532, 9.971212, 10.09594, 10.2207, 10.3455, 
    10.47035, 10.59523, 10.72016, 10.84512, 10.97012, 11.09515, 11.22022, 
    11.34533, 11.47047, 11.59565, 11.72086, 11.84611, 11.97138, 12.09669, 
    12.22203, 12.3474, 12.4728, 12.59823, 12.72368, 12.84917, 12.97468, 
    13.10022, 13.22579, 13.35138, 13.47699, 13.60263, 13.72829, 13.85398, 
    13.97969, 14.10541, 14.23116, 14.35693, 14.48272, 14.60853, 14.73435, 
    14.8602, 14.98606, 15.11193, 15.23782, 15.36373, 15.48965, 15.61558, 
    15.74153, 15.86749, 15.99346, 16.11944, 16.24543, 16.37143, 16.49744, 
    16.62345, 16.74948, 16.87551, 17.00154, 17.12758, 17.25363, 17.37968, 
    17.50574, 17.63179, 17.75785, 17.88391, 18.00997, 18.13603, 18.26209, 
    18.38815, 18.5142, 18.64026, 18.76631, 18.89235, 19.01839, 19.14443, 
    19.27046, 19.39648, 19.5225, 19.6485, 19.7745, 19.90049, 20.02647, 
    20.15244, 20.27839, 20.40434, 20.53027, 20.65619, 20.78209, 20.90798, 
    21.03385, 21.15971, 21.28555, 21.41137, 21.53718, 21.66296, 21.78873, 
    21.91447, 22.0402, 22.1659, 22.29159, 22.41724, 22.54288, 22.66849, 
    22.79408, 22.91964, 23.04517, 23.17068, 23.29616, 23.42162, 23.54704, 
    23.67244, 23.7978, 23.92313, 24.04844, 24.17371, 24.29895, 24.42415, 
    24.54932, 24.67446, 24.79956, 24.92463, 25.04966, 25.17465, 25.29961, 
    25.42452, 25.5494, 25.67424, 25.79904, 25.9238, 26.04851, 26.17319, 
    26.29782, 26.42241, 26.54695, 26.67145, 26.79591, 26.92031, 27.04468, 
    27.16899, 27.29326, 27.41748, 27.54166, 27.66578, 27.78985, 27.91387, 
    28.03784, 28.16176, 28.28563, 28.40944, 28.53321, 28.65691, 28.78057, 
    28.90416, 29.0277, 29.15119, 29.27462, 29.39799, 29.5213, 29.64455, 
    29.76775, 29.89088, 30.01396, 30.13697, 30.25993, 30.38282, 30.50564, 
    30.62841, 30.75111, 30.87375, 30.99632, 31.11883, 31.24127, 31.36365, 
    31.48596, 31.6082, 31.73037, 31.85248, 31.97452, 32.09648, 32.21838, 
    32.34021, 32.46196, 32.58365, 32.70526, 32.8268, 32.94827, 33.06966, 
    33.19098, 33.31223, 33.4334, 33.5545, 33.67552, 33.79646, 33.91733, 
    34.03812, 34.15883, 34.27946, 34.40002, 34.52049, 34.64089, 34.7612, 
    34.88144, 35.00159, 35.12167, 35.24166, 35.36156, 35.48139, 35.60114, 
    35.72079, 35.84037, 35.95986, 36.07927, 36.19859, 36.31782, 36.43697, 
    36.55603, 36.67501, 36.7939, 36.9127, 37.03141, 37.15003, 37.26857, 
    37.38701, 37.50537, 37.62363, 37.74181, 37.85989, 37.97788, 38.09578, 
    38.21359, 38.33131, 38.44893, 38.56646, 38.6839, 38.80124, 38.91849, 
    39.03564,
  -13.51432, -13.40693, -13.29943, -13.19181, -13.08407, -12.97622, 
    -12.86826, -12.76018, -12.65199, -12.54368, -12.43526, -12.32673, 
    -12.21808, -12.10931, -12.00044, -11.89145, -11.78234, -11.67312, 
    -11.56379, -11.45435, -11.34479, -11.23512, -11.12534, -11.01545, 
    -10.90544, -10.79532, -10.68509, -10.57475, -10.46429, -10.35372, 
    -10.24304, -10.13225, -10.02135, -9.91034, -9.799217, -9.687983, 
    -9.576638, -9.465184, -9.353619, -9.241944, -9.130159, -9.018265, 
    -8.906261, -8.794148, -8.681927, -8.569596, -8.457156, -8.344609, 
    -8.231953, -8.119189, -8.006317, -7.893338, -7.780252, -7.667058, 
    -7.553757, -7.44035, -7.326836, -7.213216, -7.099491, -6.985659, 
    -6.871722, -6.75768, -6.643533, -6.529281, -6.414925, -6.300464, -6.1859, 
    -6.071232, -5.95646, -5.841586, -5.726608, -5.611528, -5.496346, 
    -5.381062, -5.265676, -5.150188, -5.034599, -4.91891, -4.80312, -4.68723, 
    -4.571239, -4.45515, -4.338961, -4.222672, -4.106286, -3.9898, -3.873217, 
    -3.756536, -3.639758, -3.522882, -3.40591, -3.288842, -3.171677, 
    -3.054417, -2.937061, -2.81961, -2.702065, -2.584425, -2.466692, 
    -2.348865, -2.230944, -2.112931, -1.994826, -1.876628, -1.758338, 
    -1.639958, -1.521486, -1.402923, -1.284271, -1.165529, -1.046697, 
    -0.9277761, -0.8087668, -0.6896693, -0.570484, -0.4512114, -0.3318518, 
    -0.2124056, -0.0928733, 0.0267447, 0.146448, 0.2662361, 0.3861087, 
    0.5060652, 0.6261053, 0.7462285, 0.8664344, 0.9867225, 1.107092, 
    1.227544, 1.348076, 1.468688, 1.589381, 1.710153, 1.831004, 1.951933, 
    2.072941, 2.194026, 2.315188, 2.436428, 2.557743, 2.679134, 2.8006, 
    2.922141, 3.043756, 3.165445, 3.287207, 3.409042, 3.530949, 3.652928, 
    3.774978, 3.897098, 4.019289, 4.14155, 4.263879, 4.386278, 4.508744, 
    4.631279, 4.75388, 4.876547, 4.999281, 5.12208, 5.244944, 5.367872, 
    5.490865, 5.61392, 5.737039, 5.860219, 5.983461, 6.106764, 6.230128, 
    6.353551, 6.477034, 6.600576, 6.724176, 6.847834, 6.971549, 7.09532, 
    7.219148, 7.34303, 7.466968, 7.59096, 7.715005, 7.839104, 7.963254, 
    8.087458, 8.211712, 8.336017, 8.460371, 8.584776, 8.709229, 8.833731, 
    8.95828, 9.082876, 9.207519, 9.332207, 9.456941, 9.581719, 9.706542, 
    9.831408, 9.956316, 10.08127, 10.20626, 10.33129, 10.45637, 10.58148, 
    10.70663, 10.83182, 10.95705, 11.08232, 11.20762, 11.33296, 11.45833, 
    11.58374, 11.70918, 11.83465, 11.96016, 12.0857, 12.21127, 12.33687, 
    12.4625, 12.58816, 12.71385, 12.83957, 12.96531, 13.09109, 13.21688, 
    13.34271, 13.46856, 13.59443, 13.72032, 13.84624, 13.97218, 14.09815, 
    14.22413, 14.35013, 14.47616, 14.6022, 14.72826, 14.85433, 14.98043, 
    15.10654, 15.23267, 15.35881, 15.48496, 15.61113, 15.73731, 15.8635, 
    15.98971, 16.11592, 16.24215, 16.36838, 16.49463, 16.62088, 16.74714, 
    16.87341, 16.99968, 17.12595, 17.25224, 17.37852, 17.50481, 17.6311, 
    17.7574, 17.88369, 18.00999, 18.13629, 18.26258, 18.38887, 18.51517, 
    18.64145, 18.76774, 18.89402, 19.0203, 19.14657, 19.27283, 19.39909, 
    19.52534, 19.65158, 19.77782, 19.90404, 20.03026, 20.15646, 20.28265, 
    20.40883, 20.535, 20.66115, 20.78729, 20.91341, 21.03952, 21.16561, 
    21.29169, 21.41774, 21.54378, 21.6698, 21.7958, 21.92178, 22.04774, 
    22.17368, 22.29959, 22.42548, 22.55135, 22.6772, 22.80302, 22.92881, 
    23.05458, 23.18032, 23.30603, 23.43172, 23.55737, 23.683, 23.8086, 
    23.93416, 24.0597, 24.1852, 24.31067, 24.4361, 24.56151, 24.68687, 
    24.81221, 24.9375, 25.06276, 25.18798, 25.31317, 25.43831, 25.56342, 
    25.68849, 25.81351, 25.9385, 26.06344, 26.18835, 26.31321, 26.43802, 
    26.56279, 26.68752, 26.8122, 26.93684, 27.06143, 27.18597, 27.31046, 
    27.43491, 27.5593, 27.68365, 27.80795, 27.93219, 28.05639, 28.18053, 
    28.30462, 28.42866, 28.55264, 28.67657, 28.80044, 28.92426, 29.04803, 
    29.17173, 29.29538, 29.41897, 29.5425, 29.66598, 29.78939, 29.91274, 
    30.03604, 30.15927, 30.28244, 30.40555, 30.52859, 30.65158, 30.7745, 
    30.89735, 31.02014, 31.14286, 31.26552, 31.38811, 31.51063, 31.63309, 
    31.75548, 31.87779, 32.00005, 32.12222, 32.24434, 32.36637, 32.48834, 
    32.61024, 32.73206, 32.85381, 32.97549, 33.09709, 33.21862, 33.34007, 
    33.46145, 33.58276, 33.70398, 33.82513, 33.94621, 34.0672, 34.18812, 
    34.30896, 34.42972, 34.5504, 34.671, 34.79152, 34.91195, 35.03231, 
    35.15258, 35.27278, 35.39289, 35.51292, 35.63286, 35.75272, 35.87249, 
    35.99218, 36.11179, 36.2313, 36.35074, 36.47009, 36.58934, 36.70852, 
    36.8276, 36.94659, 37.0655, 37.18432, 37.30305, 37.42168, 37.54023, 
    37.65869, 37.77706, 37.89533, 38.01352, 38.13161, 38.2496, 38.36751, 
    38.48532, 38.60304, 38.72066, 38.8382, 38.95563, 39.07297,
  -13.56687, -13.45934, -13.3517, -13.24394, -13.13606, -13.02807, -12.91996, 
    -12.81174, -12.70341, -12.59496, -12.48639, -12.37771, -12.26892, 
    -12.16001, -12.05099, -11.94185, -11.8326, -11.72323, -11.61375, 
    -11.50416, -11.39446, -11.28464, -11.1747, -11.06466, -10.9545, 
    -10.84423, -10.73385, -10.62335, -10.51274, -10.40202, -10.29119, 
    -10.18024, -10.06919, -9.958016, -9.846737, -9.735347, -9.623845, 
    -9.512232, -9.400509, -9.288675, -9.176731, -9.064676, -8.952513, 
    -8.840239, -8.727855, -8.615362, -8.50276, -8.39005, -8.27723, -8.164302, 
    -8.051266, -7.938121, -7.824869, -7.711509, -7.598042, -7.484467, 
    -7.370786, -7.256998, -7.143103, -7.029102, -6.914995, -6.800783, 
    -6.686465, -6.572042, -6.457513, -6.342881, -6.228143, -6.113302, 
    -5.998356, -5.883307, -5.768155, -5.6529, -5.537541, -5.422081, 
    -5.306518, -5.190853, -5.075086, -4.959218, -4.843249, -4.727179, 
    -4.611009, -4.494739, -4.378368, -4.261899, -4.145329, -4.028662, 
    -3.911896, -3.795031, -3.678069, -3.561009, -3.443851, -3.326597, 
    -3.209247, -3.0918, -2.974257, -2.856619, -2.738886, -2.621058, 
    -2.503135, -2.385118, -2.267008, -2.148805, -2.030508, -1.912119, 
    -1.793638, -1.675064, -1.5564, -1.437644, -1.318798, -1.199861, 
    -1.080835, -0.9617189, -0.8425139, -0.7232202, -0.6038383, -0.4843686, 
    -0.3648115, -0.2451673, -0.1254366, -0.005619704, 0.1142829, 0.2342709, 
    0.3543437, 0.474501, 0.5947422, 0.715067, 0.835475, 0.9559656, 1.076538, 
    1.197193, 1.317929, 1.438746, 1.559643, 1.68062, 1.801676, 1.922812, 
    2.044026, 2.165318, 2.286688, 2.408134, 2.529658, 2.651257, 2.772932, 
    2.894682, 3.016507, 3.138406, 3.260379, 3.382425, 3.504543, 3.626734, 
    3.748996, 3.871329, 3.993733, 4.116207, 4.23875, 4.361362, 4.484044, 
    4.606792, 4.729609, 4.852492, 4.975441, 5.098457, 5.221538, 5.344683, 
    5.467893, 5.591166, 5.714502, 5.837901, 5.961362, 6.084884, 6.208467, 
    6.33211, 6.455813, 6.579576, 6.703397, 6.827276, 6.951212, 7.075205, 
    7.199255, 7.323359, 7.44752, 7.571735, 7.696003, 7.820325, 7.9447, 
    8.069127, 8.193606, 8.318135, 8.442716, 8.567346, 8.692024, 8.816751, 
    8.941527, 9.06635, 9.191219, 9.316134, 9.441096, 9.566102, 9.691152, 
    9.816246, 9.941382, 10.06656, 10.19178, 10.31705, 10.44235, 10.56769, 
    10.69307, 10.81849, 10.94395, 11.06945, 11.19498, 11.32055, 11.44615, 
    11.57179, 11.69746, 11.82317, 11.94891, 12.07468, 12.20048, 12.32631, 
    12.45218, 12.57807, 12.70399, 12.82994, 12.95592, 13.08193, 13.20796, 
    13.33402, 13.4601, 13.5862, 13.71233, 13.83849, 13.96466, 14.09086, 
    14.21708, 14.34332, 14.46957, 14.59585, 14.72214, 14.84846, 14.97478, 
    15.10113, 15.22749, 15.35387, 15.48026, 15.60666, 15.73308, 15.85951, 
    15.98595, 16.1124, 16.23886, 16.36533, 16.49181, 16.6183, 16.74479, 
    16.8713, 16.9978, 17.12432, 17.25084, 17.37736, 17.50389, 17.63041, 
    17.75694, 17.88348, 18.01001, 18.13654, 18.26307, 18.3896, 18.51613, 
    18.64265, 18.76918, 18.89569, 19.02221, 19.14871, 19.27522, 19.40171, 
    19.5282, 19.65467, 19.78114, 19.9076, 20.03405, 20.16049, 20.28692, 
    20.41333, 20.53974, 20.66612, 20.7925, 20.91886, 21.0452, 21.17153, 
    21.29784, 21.42413, 21.5504, 21.67665, 21.80289, 21.9291, 22.0553, 
    22.18147, 22.30762, 22.43374, 22.55985, 22.68592, 22.81198, 22.93801, 
    23.06401, 23.18998, 23.31593, 23.44184, 23.56773, 23.69359, 23.81942, 
    23.94522, 24.07098, 24.19672, 24.32242, 24.44809, 24.57372, 24.69932, 
    24.82488, 24.95041, 25.0759, 25.20135, 25.32676, 25.45214, 25.57748, 
    25.70277, 25.82803, 25.95324, 26.07841, 26.20354, 26.32863, 26.45367, 
    26.57867, 26.70363, 26.82854, 26.9534, 27.07821, 27.20298, 27.3277, 
    27.45237, 27.57699, 27.70157, 27.82609, 27.95056, 28.07498, 28.19934, 
    28.32366, 28.44792, 28.57212, 28.69628, 28.82037, 28.94441, 29.0684, 
    29.19232, 29.31619, 29.44001, 29.56376, 29.68745, 29.81109, 29.93466, 
    30.05817, 30.18162, 30.30501, 30.42834, 30.5516, 30.6748, 30.79794, 
    30.92101, 31.04401, 31.16695, 31.28982, 31.41263, 31.53537, 31.65804, 
    31.78064, 31.90317, 32.02563, 32.14803, 32.27035, 32.3926, 32.51478, 
    32.63689, 32.75892, 32.88088, 33.00277, 33.12458, 33.24632, 33.36798, 
    33.48957, 33.61108, 33.73252, 33.85387, 33.97515, 34.09636, 34.21748, 
    34.33852, 34.45949, 34.58037, 34.70118, 34.8219, 34.94254, 35.0631, 
    35.18358, 35.30397, 35.42428, 35.54451, 35.66465, 35.78471, 35.90469, 
    36.02458, 36.14438, 36.2641, 36.38373, 36.50327, 36.62273, 36.7421, 
    36.86138, 36.98057, 37.09967, 37.21868, 37.3376, 37.45644, 37.57518, 
    37.69383, 37.81239, 37.93085, 38.04923, 38.16751, 38.2857, 38.40379, 
    38.52179, 38.6397, 38.75751, 38.87523, 38.99286, 39.11039,
  -13.61951, -13.51184, -13.40406, -13.29616, -13.18814, -13.08001, 
    -12.97176, -12.8634, -12.75492, -12.64633, -12.53762, -12.42879, 
    -12.31985, -12.2108, -12.10163, -11.99235, -11.88295, -11.77344, 
    -11.66381, -11.55407, -11.44421, -11.33424, -11.22416, -11.11397, 
    -11.00366, -10.89323, -10.7827, -10.67205, -10.56129, -10.45041, 
    -10.33942, -10.22832, -10.11711, -10.00579, -9.894351, -9.782804, 
    -9.671144, -9.559374, -9.447492, -9.335499, -9.223395, -9.111181, 
    -8.998857, -8.886421, -8.773876, -8.661221, -8.548456, -8.435582, 
    -8.322599, -8.209507, -8.096306, -7.982996, -7.869578, -7.756052, 
    -7.642417, -7.528676, -7.414826, -7.300869, -7.186806, -7.072636, 
    -6.958359, -6.843976, -6.729487, -6.614892, -6.500192, -6.385386, 
    -6.270476, -6.155461, -6.040341, -5.925118, -5.80979, -5.694359, 
    -5.578825, -5.463187, -5.347447, -5.231604, -5.115659, -4.999612, 
    -4.883464, -4.767215, -4.650864, -4.534413, -4.417861, -4.30121, 
    -4.184459, -4.067608, -3.950659, -3.833611, -3.716464, -3.599219, 
    -3.481876, -3.364436, -3.2469, -3.129266, -3.011536, -2.89371, -2.775788, 
    -2.657772, -2.53966, -2.421453, -2.303153, -2.184758, -2.066271, 
    -1.94769, -1.829016, -1.71025, -1.591393, -1.472443, -1.353403, 
    -1.234272, -1.11505, -0.995739, -0.8763381, -0.7568479, -0.6372691, 
    -0.517602, -0.397847, -0.2780045, -0.158075, -0.03805884, 0.0820435, 
    0.2022316, 0.3225051, 0.4428634, 0.5633062, 0.6838329, 0.8044433, 
    0.9251368, 1.045913, 1.166771, 1.287711, 1.408733, 1.529835, 1.651018, 
    1.77228, 1.893622, 2.015043, 2.136542, 2.258119, 2.379774, 2.501506, 
    2.623314, 2.745199, 2.867159, 2.989194, 3.111303, 3.233487, 3.355744, 
    3.478074, 3.600477, 3.722951, 3.845498, 3.968115, 4.090803, 4.21356, 
    4.336387, 4.459283, 4.582247, 4.705279, 4.828378, 4.951544, 5.074776, 
    5.198074, 5.321437, 5.444864, 5.568356, 5.691911, 5.815528, 5.939209, 
    6.06295, 6.186753, 6.310617, 6.434541, 6.558524, 6.682566, 6.806666, 
    6.930825, 7.05504, 7.179312, 7.30364, 7.428024, 7.552462, 7.676955, 
    7.801501, 7.9261, 8.050752, 8.175455, 8.30021, 8.425015, 8.549871, 
    8.674777, 8.79973, 8.924732, 9.049782, 9.174879, 9.300022, 9.425211, 
    9.550445, 9.675723, 9.801045, 9.926412, 10.05182, 10.17727, 10.30276, 
    10.42829, 10.55387, 10.67948, 10.80513, 10.93082, 11.05655, 11.18231, 
    11.30811, 11.43394, 11.55981, 11.68572, 11.81166, 11.93763, 12.06363, 
    12.18967, 12.31573, 12.44183, 12.56796, 12.69411, 12.8203, 12.94651, 
    13.07275, 13.19901, 13.3253, 13.45162, 13.57796, 13.70432, 13.83071, 
    13.95712, 14.08355, 14.21001, 14.33648, 14.46297, 14.58948, 14.71601, 
    14.84256, 14.96913, 15.09571, 15.22231, 15.34892, 15.47554, 15.60218, 
    15.72884, 15.8555, 15.98218, 16.10887, 16.23557, 16.36227, 16.48899, 
    16.61571, 16.74244, 16.86918, 16.99593, 17.12268, 17.24944, 17.37619, 
    17.50296, 17.62972, 17.75649, 17.88326, 18.01003, 18.1368, 18.26356, 
    18.39033, 18.5171, 18.64386, 18.77062, 18.89737, 19.02412, 19.15086, 
    19.2776, 19.40433, 19.53106, 19.65777, 19.78448, 19.91117, 20.03786, 
    20.16454, 20.2912, 20.41785, 20.54449, 20.67111, 20.79772, 20.92432, 
    21.05089, 21.17746, 21.304, 21.43053, 21.55704, 21.68353, 21.81, 
    21.93645, 22.06288, 22.18928, 22.31567, 22.44203, 22.56836, 22.69468, 
    22.82096, 22.94722, 23.07346, 23.19967, 23.32585, 23.452, 23.57812, 
    23.70421, 23.83027, 23.9563, 24.0823, 24.20827, 24.3342, 24.4601, 
    24.58596, 24.71179, 24.83759, 24.96335, 25.08907, 25.21475, 25.34039, 
    25.466, 25.59157, 25.71709, 25.84258, 25.96802, 26.09342, 26.21878, 
    26.3441, 26.46937, 26.59459, 26.71978, 26.84491, 26.97, 27.09504, 
    27.22004, 27.34498, 27.46988, 27.59473, 27.71953, 27.84427, 27.96897, 
    28.09361, 28.2182, 28.34274, 28.46723, 28.59166, 28.71603, 28.84035, 
    28.96461, 29.08882, 29.21297, 29.33706, 29.46109, 29.58507, 29.70898, 
    29.83283, 29.95663, 30.08036, 30.20403, 30.32764, 30.45118, 30.57467, 
    30.69808, 30.82143, 30.94472, 31.06794, 31.1911, 31.31419, 31.43721, 
    31.56016, 31.68305, 31.80586, 31.92861, 32.05128, 32.17389, 32.29643, 
    32.41889, 32.54128, 32.6636, 32.78585, 32.90802, 33.03012, 33.15214, 
    33.27409, 33.39596, 33.51775, 33.63948, 33.76112, 33.88268, 34.00417, 
    34.12558, 34.24691, 34.36816, 34.48933, 34.61042, 34.73143, 34.85235, 
    34.9732, 35.09396, 35.21464, 35.33524, 35.45575, 35.57618, 35.69653, 
    35.81679, 35.93696, 36.05705, 36.17705, 36.29697, 36.4168, 36.53654, 
    36.65619, 36.77576, 36.89523, 37.01462, 37.13391, 37.25312, 37.37224, 
    37.49126, 37.6102, 37.72904, 37.84779, 37.96645, 38.08502, 38.20349, 
    38.32187, 38.44016, 38.55835, 38.67645, 38.79445, 38.91235, 39.03017, 
    39.14788,
  -13.67225, -13.56444, -13.45652, -13.34848, -13.24032, -13.13205, 
    -13.02366, -12.91515, -12.80653, -12.69779, -12.58894, -12.47997, 
    -12.37088, -12.26168, -12.15237, -12.04294, -11.93339, -11.82373, 
    -11.71396, -11.60407, -11.49407, -11.38395, -11.27371, -11.16337, 
    -11.05291, -10.94233, -10.83164, -10.72084, -10.60993, -10.4989, 
    -10.38775, -10.2765, -10.16513, -10.05365, -9.94206, -9.830355, 
    -9.718538, -9.606609, -9.494569, -9.382417, -9.270153, -9.157779, 
    -9.045293, -8.932697, -8.81999, -8.707172, -8.594245, -8.481208, 
    -8.368061, -8.254804, -8.141438, -8.027963, -7.914379, -7.800686, 
    -7.686884, -7.572975, -7.458958, -7.344832, -7.2306, -7.11626, -7.001813, 
    -6.887259, -6.772599, -6.657833, -6.54296, -6.427982, -6.312898, 
    -6.19771, -6.082416, -5.967017, -5.851514, -5.735907, -5.620196, 
    -5.504382, -5.388464, -5.272444, -5.15632, -5.040094, -4.923767, 
    -4.807337, -4.690806, -4.574174, -4.457441, -4.340608, -4.223674, 
    -4.10664, -3.989507, -3.872275, -3.754943, -3.637514, -3.519985, 
    -3.402359, -3.284636, -3.166815, -3.048898, -2.930884, -2.812774, 
    -2.694568, -2.576266, -2.45787, -2.339379, -2.220793, -2.102114, 
    -1.983341, -1.864475, -1.745517, -1.626465, -1.507322, -1.388087, 
    -1.268761, -1.149344, -1.029837, -0.9102398, -0.7905529, -0.6707768, 
    -0.550912, -0.4309588, -0.3109176, -0.190789, -0.0705732, 0.04972921, 
    0.1701178, 0.2905923, 0.411152, 0.5317967, 0.6525258, 0.773339, 
    0.8942357, 1.015216, 1.136278, 1.257423, 1.378649, 1.499957, 1.621345, 
    1.742814, 1.864363, 1.985991, 2.107698, 2.229483, 2.351346, 2.473287, 
    2.595305, 2.717399, 2.839569, 2.961815, 3.084135, 3.20653, 3.328999, 
    3.451541, 3.574157, 3.696844, 3.819604, 3.942435, 4.065337, 4.188309, 
    4.311351, 4.434462, 4.557642, 4.68089, 4.804205, 4.927588, 5.051038, 
    5.174553, 5.298134, 5.42178, 5.54549, 5.669263, 5.793101, 5.917, 
    6.040962, 6.164986, 6.28907, 6.413215, 6.53742, 6.661684, 6.786006, 
    6.910387, 7.034825, 7.15932, 7.283872, 7.408479, 7.533141, 7.657858, 
    7.782629, 7.907454, 8.032331, 8.15726, 8.28224, 8.407272, 8.532354, 
    8.657486, 8.782666, 8.907896, 9.033174, 9.158498, 9.283869, 9.409286, 
    9.534748, 9.660255, 9.785808, 9.911403, 10.03704, 10.16272, 10.28844, 
    10.4142, 10.54001, 10.66585, 10.79173, 10.91765, 11.04361, 11.16961, 
    11.29564, 11.4217, 11.54781, 11.67394, 11.80011, 11.92632, 12.05256, 
    12.17882, 12.30512, 12.43145, 12.55781, 12.6842, 12.81062, 12.93707, 
    13.06354, 13.19004, 13.31657, 13.44312, 13.56969, 13.69629, 13.82292, 
    13.94956, 14.07623, 14.20292, 14.32963, 14.45636, 14.5831, 14.70987, 
    14.83665, 14.96346, 15.09027, 15.21711, 15.34396, 15.47082, 15.5977, 
    15.72458, 15.85149, 15.9784, 16.10533, 16.23226, 16.35921, 16.48616, 
    16.61312, 16.74009, 16.86707, 16.99405, 17.12104, 17.24803, 17.37502, 
    17.50203, 17.62903, 17.75603, 17.88304, 18.01005, 18.13705, 18.26406, 
    18.39106, 18.51806, 18.64506, 18.77206, 18.89905, 19.02604, 19.15302, 
    19.27999, 19.40696, 19.53392, 19.66088, 19.78782, 19.91475, 20.04168, 
    20.16859, 20.29549, 20.42238, 20.54925, 20.67611, 20.80296, 20.92979, 
    21.0566, 21.1834, 21.31018, 21.43695, 21.56369, 21.69042, 21.81712, 
    21.94381, 22.07047, 22.19711, 22.32373, 22.45033, 22.5769, 22.70345, 
    22.82997, 22.95647, 23.08294, 23.20938, 23.33579, 23.46218, 23.58853, 
    23.71486, 23.84115, 23.96741, 24.09365, 24.21984, 24.34601, 24.47214, 
    24.59824, 24.7243, 24.85033, 24.97632, 25.10227, 25.22818, 25.35406, 
    25.47989, 25.60569, 25.73145, 25.85716, 25.98284, 26.10847, 26.23406, 
    26.3596, 26.4851, 26.61056, 26.73597, 26.86133, 26.98665, 27.11192, 
    27.23714, 27.36231, 27.48744, 27.61251, 27.73753, 27.8625, 27.98743, 
    28.1123, 28.23711, 28.36187, 28.48658, 28.61124, 28.73583, 28.86038, 
    28.98486, 29.10929, 29.23366, 29.35798, 29.48223, 29.60643, 29.73056, 
    29.85464, 29.97865, 30.1026, 30.22649, 30.35032, 30.47408, 30.59778, 
    30.72142, 30.84499, 30.96849, 31.09193, 31.21531, 31.33861, 31.46185, 
    31.58502, 31.70812, 31.83115, 31.95411, 32.077, 32.19982, 32.32257, 
    32.44524, 32.56785, 32.69038, 32.81284, 32.93522, 33.05753, 33.17976, 
    33.30192, 33.424, 33.54601, 33.66793, 33.78979, 33.91156, 34.03325, 
    34.15487, 34.27641, 34.39786, 34.51924, 34.64053, 34.76175, 34.88288, 
    35.00393, 35.12489, 35.24578, 35.36658, 35.48729, 35.60793, 35.72847, 
    35.84893, 35.96931, 36.0896, 36.2098, 36.32991, 36.44994, 36.56988, 
    36.68973, 36.80949, 36.92916, 37.04875, 37.16824, 37.28764, 37.40696, 
    37.52618, 37.6453, 37.76434, 37.88329, 38.00214, 38.1209, 38.23956, 
    38.35813, 38.4766, 38.59499, 38.71327, 38.83146, 38.94956, 39.06756, 
    39.18546,
  -13.72509, -13.61714, -13.50908, -13.40089, -13.2926, -13.18418, -13.07565, 
    -12.967, -12.85823, -12.74935, -12.64036, -12.53124, -12.42201, 
    -12.31267, -12.20321, -12.09363, -11.98394, -11.87413, -11.7642, 
    -11.65417, -11.54401, -11.43375, -11.32336, -11.21286, -11.10225, 
    -10.99152, -10.88068, -10.76973, -10.65866, -10.54748, -10.43618, 
    -10.32477, -10.21325, -10.10161, -9.989862, -9.878, -9.766026, -9.653939, 
    -9.54174, -9.429429, -9.317005, -9.204471, -9.091825, -8.979067, 
    -8.866198, -8.753218, -8.640127, -8.526927, -8.413615, -8.300194, 
    -8.186663, -8.073022, -7.959272, -7.845413, -7.731444, -7.617367, 
    -7.503181, -7.388887, -7.274486, -7.159976, -7.045359, -6.930634, 
    -6.815803, -6.700864, -6.585819, -6.470668, -6.355411, -6.240048, 
    -6.124579, -6.009006, -5.893328, -5.777544, -5.661657, -5.545665, 
    -5.42957, -5.313371, -5.197069, -5.080665, -4.964157, -4.847547, 
    -4.730835, -4.614022, -4.497108, -4.380092, -4.262975, -4.145758, 
    -4.028441, -3.911025, -3.793508, -3.675893, -3.558179, -3.440367, 
    -3.322457, -3.204449, -3.086343, -2.968141, -2.849842, -2.731447, 
    -2.612955, -2.494369, -2.375687, -2.25691, -2.138039, -2.019074, 
    -1.900015, -1.780863, -1.661618, -1.542281, -1.422851, -1.30333, 
    -1.183717, -1.064014, -0.9442197, -0.8243357, -0.704362, -0.584299, 
    -0.4641473, -0.3439071, -0.2235789, -0.1031632, 0.01733959, 0.1379291, 
    0.2586049, 0.3793665, 0.5002134, 0.6211452, 0.7421616, 0.8632619, 
    0.9844458, 1.105713, 1.227062, 1.348494, 1.470008, 1.591603, 1.713278, 
    1.835034, 1.95687, 2.078785, 2.200778, 2.322851, 2.445001, 2.567228, 
    2.689532, 2.811913, 2.93437, 3.056901, 3.179508, 3.302189, 3.424944, 
    3.547773, 3.670674, 3.793647, 3.916692, 4.039809, 4.162996, 4.286253, 
    4.40958, 4.532976, 4.656441, 4.779974, 4.903574, 5.027241, 5.150974, 
    5.274774, 5.398638, 5.522567, 5.646561, 5.770617, 5.894738, 6.01892, 
    6.143165, 6.26747, 6.391837, 6.516263, 6.640749, 6.765295, 6.889898, 
    7.01456, 7.139278, 7.264054, 7.388885, 7.513772, 7.638714, 7.76371, 
    7.88876, 8.013863, 8.139018, 8.264225, 8.389483, 8.514792, 8.640151, 
    8.765559, 8.891017, 9.016522, 9.142075, 9.267674, 9.393321, 9.519012, 
    9.644749, 9.770531, 9.896355, 10.02222, 10.14813, 10.27409, 10.40008, 
    10.52611, 10.65219, 10.7783, 10.90445, 11.03064, 11.15687, 11.28313, 
    11.40943, 11.53577, 11.66214, 11.78854, 11.91498, 12.04145, 12.16795, 
    12.29449, 12.42105, 12.54765, 12.67427, 12.80092, 12.92761, 13.05431, 
    13.18105, 13.30781, 13.4346, 13.56141, 13.68824, 13.8151, 13.94198, 
    14.06889, 14.19581, 14.32276, 14.44972, 14.57671, 14.70371, 14.83073, 
    14.95777, 15.08482, 15.21189, 15.33898, 15.46608, 15.59319, 15.72032, 
    15.84746, 15.97461, 16.10177, 16.22895, 16.35613, 16.48332, 16.61052, 
    16.73773, 16.86494, 16.99216, 17.11939, 17.24662, 17.37385, 17.50109, 
    17.62833, 17.75558, 17.88282, 18.01006, 18.13731, 18.26455, 18.3918, 
    18.51904, 18.64627, 18.77351, 18.90074, 19.02796, 19.15518, 19.28239, 
    19.4096, 19.5368, 19.66399, 19.79117, 19.91834, 20.0455, 20.17265, 
    20.29979, 20.42691, 20.55403, 20.68112, 20.80821, 20.93528, 21.06233, 
    21.18936, 21.31638, 21.44338, 21.57036, 21.69733, 21.82427, 21.95119, 
    22.07809, 22.20497, 22.33182, 22.45865, 22.58546, 22.71224, 22.839, 
    22.96573, 23.09244, 23.21911, 23.34576, 23.47238, 23.59897, 23.72553, 
    23.85206, 23.97856, 24.10502, 24.23145, 24.35785, 24.48422, 24.61055, 
    24.73684, 24.8631, 24.98932, 25.11551, 25.24165, 25.36776, 25.49383, 
    25.61985, 25.74584, 25.87179, 25.99769, 26.12355, 26.24937, 26.37514, 
    26.50087, 26.62656, 26.7522, 26.87779, 27.00333, 27.12883, 27.25428, 
    27.37968, 27.50503, 27.63033, 27.75558, 27.88078, 28.00593, 28.13103, 
    28.25607, 28.38105, 28.50599, 28.63087, 28.75569, 28.88045, 29.00516, 
    29.12982, 29.25441, 29.37895, 29.50342, 29.62784, 29.7522, 29.87649, 
    30.00073, 30.1249, 30.24901, 30.37306, 30.49704, 30.62096, 30.74481, 
    30.8686, 30.99233, 31.11598, 31.23957, 31.36309, 31.48655, 31.60993, 
    31.73325, 31.85649, 31.97967, 32.10278, 32.22581, 32.34877, 32.47166, 
    32.59448, 32.71722, 32.83989, 32.96249, 33.08501, 33.20745, 33.32982, 
    33.45211, 33.57433, 33.69646, 33.81852, 33.94051, 34.06241, 34.18423, 
    34.30597, 34.42764, 34.54922, 34.67072, 34.79214, 34.91348, 35.03473, 
    35.1559, 35.27699, 35.39799, 35.51891, 35.63974, 35.76049, 35.88115, 
    36.00173, 36.12222, 36.24262, 36.36293, 36.48316, 36.6033, 36.72335, 
    36.8433, 36.96318, 37.08295, 37.20264, 37.32224, 37.44175, 37.56116, 
    37.68049, 37.79972, 37.91885, 38.0379, 38.15685, 38.2757, 38.39447, 
    38.51313, 38.63171, 38.75018, 38.86856, 38.98685, 39.10503, 39.22312,
  -13.77802, -13.66993, -13.56173, -13.45341, -13.34497, -13.23641, 
    -13.12774, -13.01895, -12.91004, -12.80101, -12.69187, -12.58261, 
    -12.47324, -12.36375, -12.25414, -12.14441, -12.03458, -11.92462, 
    -11.81455, -11.70436, -11.59406, -11.48364, -11.37311, -11.26246, 
    -11.15169, -11.04082, -10.92982, -10.81871, -10.70749, -10.59615, 
    -10.4847, -10.37314, -10.26146, -10.14967, -10.03776, -9.925742, 
    -9.81361, -9.701365, -9.589006, -9.476536, -9.363953, -9.251257, 
    -9.13845, -9.025531, -8.912499, -8.799357, -8.686104, -8.57274, 
    -8.459264, -8.345678, -8.231981, -8.118176, -8.004259, -7.890233, 
    -7.776097, -7.661852, -7.547498, -7.433035, -7.318463, -7.203784, 
    -7.088996, -6.974101, -6.859097, -6.743987, -6.628769, -6.513445, 
    -6.398014, -6.282477, -6.166834, -6.051085, -5.935231, -5.819272, 
    -5.703207, -5.587039, -5.470765, -5.354388, -5.237907, -5.121323, 
    -5.004635, -4.887845, -4.770953, -4.653958, -4.536861, -4.419662, 
    -4.302363, -4.184963, -4.067461, -3.94986, -3.832159, -3.714358, 
    -3.596458, -3.478459, -3.360362, -3.242166, -3.123873, -3.005482, 
    -2.886994, -2.768409, -2.649728, -2.53095, -2.412077, -2.293109, 
    -2.174046, -2.054888, -1.935636, -1.81629, -1.696851, -1.577319, 
    -1.457695, -1.337978, -1.218169, -1.098269, -0.9782782, -0.8581967, 
    -0.7380251, -0.6177637, -0.497413, -0.3769735, -0.2564455, -0.1358295, 
    -0.01512585, 0.1056649, 0.2265424, 0.3475061, 0.4685557, 0.5896906, 
    0.7109105, 0.8322149, 0.9536032, 1.075075, 1.19663, 1.318268, 1.439988, 
    1.561789, 1.683672, 1.805635, 1.927679, 2.049802, 2.172005, 2.294286, 
    2.416646, 2.539084, 2.661599, 2.78419, 2.906858, 3.029602, 3.152421, 
    3.275315, 3.398283, 3.521325, 3.64444, 3.767627, 3.890887, 4.014219, 
    4.137621, 4.261095, 4.384638, 4.50825, 4.631932, 4.755682, 4.8795, 
    5.003385, 5.127337, 5.251355, 5.375439, 5.499588, 5.623802, 5.748079, 
    5.87242, 5.996823, 6.121289, 6.245816, 6.370405, 6.495054, 6.619763, 
    6.744532, 6.869359, 6.994244, 7.119186, 7.244186, 7.369243, 7.494355, 
    7.619522, 7.744743, 7.870019, 7.995348, 8.12073, 8.246164, 8.37165, 
    8.497186, 8.622773, 8.748409, 8.874095, 8.999828, 9.12561, 9.251439, 
    9.377315, 9.503236, 9.629203, 9.755215, 9.881269, 10.00737, 10.13351, 
    10.25969, 10.38592, 10.51218, 10.63849, 10.76484, 10.89122, 11.01764, 
    11.1441, 11.2706, 11.39713, 11.5237, 11.65031, 11.77694, 11.90361, 
    12.03032, 12.15706, 12.28382, 12.41062, 12.53745, 12.66431, 12.7912, 
    12.91812, 13.04506, 13.17203, 13.29903, 13.42605, 13.5531, 13.68017, 
    13.80727, 13.93438, 14.06152, 14.18869, 14.31587, 14.44307, 14.57029, 
    14.69753, 14.82479, 14.95207, 15.07936, 15.20667, 15.33399, 15.46133, 
    15.58868, 15.71605, 15.84342, 15.97081, 16.09822, 16.22563, 16.35305, 
    16.48048, 16.60791, 16.73536, 16.86281, 16.99027, 17.11773, 17.2452, 
    17.37268, 17.50015, 17.62763, 17.75512, 17.8826, 18.01008, 18.13757, 
    18.26505, 18.39253, 18.52001, 18.64749, 18.77496, 18.90243, 19.02989, 
    19.15735, 19.2848, 19.41224, 19.53968, 19.66711, 19.79453, 19.92194, 
    20.04934, 20.17673, 20.3041, 20.43147, 20.55882, 20.68615, 20.81347, 
    20.94078, 21.06807, 21.19534, 21.3226, 21.44983, 21.57705, 21.70425, 
    21.83143, 21.95859, 22.08573, 22.21284, 22.33993, 22.467, 22.59404, 
    22.72106, 22.84805, 22.97502, 23.10196, 23.22887, 23.35576, 23.48261, 
    23.60944, 23.73623, 23.86299, 23.98973, 24.11642, 24.24309, 24.36972, 
    24.49632, 24.62288, 24.74941, 24.8759, 25.00236, 25.12877, 25.25515, 
    25.38149, 25.50779, 25.63405, 25.76027, 25.88645, 26.01258, 26.13867, 
    26.26472, 26.39073, 26.51669, 26.6426, 26.76847, 26.89429, 27.02006, 
    27.14579, 27.27147, 27.3971, 27.52267, 27.6482, 27.77368, 27.89911, 
    28.02448, 28.1498, 28.27507, 28.40028, 28.52544, 28.65054, 28.77559, 
    28.90058, 29.02551, 29.15039, 29.27521, 29.39997, 29.52467, 29.64931, 
    29.77389, 29.8984, 30.02286, 30.14725, 30.27158, 30.39585, 30.52005, 
    30.64419, 30.76827, 30.89227, 31.01622, 31.14009, 31.2639, 31.38764, 
    31.51131, 31.63491, 31.75844, 31.8819, 32.00529, 32.12862, 32.25187, 
    32.37504, 32.49814, 32.62117, 32.74413, 32.86701, 32.98982, 33.11255, 
    33.23521, 33.35779, 33.48029, 33.60271, 33.72506, 33.84733, 33.96952, 
    34.09163, 34.21366, 34.33561, 34.45749, 34.57927, 34.70098, 34.82261, 
    34.94415, 35.06561, 35.18698, 35.30827, 35.42948, 35.5506, 35.67163, 
    35.79258, 35.91345, 36.03423, 36.15491, 36.27552, 36.39603, 36.51646, 
    36.6368, 36.75704, 36.8772, 36.99726, 37.11724, 37.23713, 37.35692, 
    37.47662, 37.59623, 37.71575, 37.83517, 37.95451, 38.07374, 38.19289, 
    38.31194, 38.43089, 38.54974, 38.66851, 38.78717, 38.90574, 39.02422, 
    39.14259, 39.26087,
  -13.83105, -13.72283, -13.61448, -13.50602, -13.39744, -13.28874, 
    -13.17992, -13.07099, -12.96194, -12.85277, -12.74348, -12.63408, 
    -12.52456, -12.41492, -12.30517, -12.1953, -12.08531, -11.97521, 
    -11.86499, -11.75465, -11.6442, -11.53363, -11.42295, -11.31215, 
    -11.20123, -11.0902, -10.97906, -10.86779, -10.75642, -10.64493, 
    -10.53332, -10.4216, -10.30977, -10.19782, -10.08576, -9.973579, 
    -9.861289, -9.748885, -9.636368, -9.523738, -9.410995, -9.298139, 
    -9.18517, -9.072089, -8.958897, -8.845592, -8.732175, -8.618647, 
    -8.505007, -8.391256, -8.277394, -8.163422, -8.049339, -7.935146, 
    -7.820843, -7.706429, -7.591907, -7.477275, -7.362534, -7.247684, 
    -7.132726, -7.017659, -6.902484, -6.787201, -6.671811, -6.556314, 
    -6.440709, -6.324997, -6.209179, -6.093255, -5.977225, -5.861089, 
    -5.744848, -5.628501, -5.51205, -5.395494, -5.278834, -5.16207, 
    -5.045203, -4.928232, -4.811158, -4.693981, -4.576702, -4.459321, 
    -4.341838, -4.224254, -4.106569, -3.988783, -3.870896, -3.752909, 
    -3.634823, -3.516637, -3.398353, -3.279969, -3.161487, -3.042907, 
    -2.92423, -2.805455, -2.686583, -2.567615, -2.44855, -2.32939, -2.210135, 
    -2.090784, -1.971338, -1.851799, -1.732165, -1.612438, -1.492618, 
    -1.372706, -1.252701, -1.132604, -1.012416, -0.8921365, -0.7717665, 
    -0.6513064, -0.5307565, -0.4101172, -0.289389, -0.1685724, -0.0476676, 
    0.07332477, 0.1944043, 0.3155706, 0.4368232, 0.5581616, 0.6795854, 
    0.8010941, 0.9226874, 1.044365, 1.166125, 1.287969, 1.409896, 1.531904, 
    1.653994, 1.776166, 1.898418, 2.02075, 2.143162, 2.265653, 2.388223, 
    2.510871, 2.633597, 2.7564, 2.87928, 3.002236, 3.125268, 3.248375, 
    3.371556, 3.494812, 3.618141, 3.741544, 3.865019, 3.988566, 4.112185, 
    4.235874, 4.359634, 4.483464, 4.607363, 4.731331, 4.855367, 4.979471, 
    5.103642, 5.22788, 5.352183, 5.476552, 5.600986, 5.725484, 5.850046, 
    5.974671, 6.099359, 6.224109, 6.34892, 6.473792, 6.598724, 6.723716, 
    6.848767, 6.973876, 7.099044, 7.224269, 7.34955, 7.474888, 7.600281, 
    7.725729, 7.851231, 7.976787, 8.102396, 8.228058, 8.353771, 8.479535, 
    8.60535, 8.731215, 8.85713, 8.983093, 9.109104, 9.235163, 9.361268, 
    9.48742, 9.613617, 9.73986, 9.866145, 9.992476, 10.11885, 10.24526, 
    10.37172, 10.49822, 10.62476, 10.75134, 10.87795, 11.00461, 11.1313, 
    11.25803, 11.3848, 11.5116, 11.63844, 11.76531, 11.89222, 12.01916, 
    12.14613, 12.27313, 12.40017, 12.52723, 12.65433, 12.78145, 12.9086, 
    13.03578, 13.16299, 13.29023, 13.41748, 13.54477, 13.67208, 13.79941, 
    13.92676, 14.05414, 14.18154, 14.30896, 14.4364, 14.56386, 14.69134, 
    14.81884, 14.94635, 15.07388, 15.20143, 15.32899, 15.45657, 15.58416, 
    15.71176, 15.83938, 15.96701, 16.09464, 16.2223, 16.34995, 16.47762, 
    16.6053, 16.73299, 16.86068, 16.98838, 17.11608, 17.24379, 17.3715, 
    17.49922, 17.62694, 17.75466, 17.88238, 18.0101, 18.13783, 18.26555, 
    18.39327, 18.52099, 18.6487, 18.77641, 18.90412, 19.03182, 19.15952, 
    19.28721, 19.4149, 19.54257, 19.67024, 19.7979, 19.92555, 20.05318, 
    20.18081, 20.30843, 20.43603, 20.56362, 20.69119, 20.81875, 20.94629, 
    21.07382, 21.20133, 21.32883, 21.4563, 21.58376, 21.7112, 21.83861, 
    21.96601, 22.09338, 22.22073, 22.34806, 22.47537, 22.60265, 22.7299, 
    22.85713, 22.98433, 23.11151, 23.23866, 23.36578, 23.49287, 23.61993, 
    23.74696, 23.87396, 24.00092, 24.12786, 24.25476, 24.38163, 24.50846, 
    24.63526, 24.76202, 24.88874, 25.01543, 25.14208, 25.26869, 25.39526, 
    25.52179, 25.64828, 25.77474, 25.90114, 26.02751, 26.15383, 26.28011, 
    26.40635, 26.53254, 26.65868, 26.78478, 26.91083, 27.03684, 27.16279, 
    27.2887, 27.41455, 27.54036, 27.66612, 27.79182, 27.91748, 28.04308, 
    28.16862, 28.29412, 28.41956, 28.54494, 28.67027, 28.79554, 28.92076, 
    29.04592, 29.17102, 29.29606, 29.42104, 29.54597, 29.67083, 29.79563, 
    29.92037, 30.04505, 30.16966, 30.29421, 30.4187, 30.54313, 30.66748, 
    30.79178, 30.916, 31.04016, 31.16426, 31.28828, 31.41224, 31.53613, 
    31.65995, 31.7837, 31.90738, 32.03098, 32.15452, 32.27798, 32.40137, 
    32.52469, 32.64793, 32.7711, 32.8942, 33.01722, 33.14016, 33.26303, 
    33.38582, 33.50853, 33.63117, 33.75373, 33.87621, 33.99861, 34.12093, 
    34.24316, 34.36532, 34.4874, 34.6094, 34.73131, 34.85314, 34.97489, 
    35.09655, 35.21813, 35.33963, 35.46104, 35.58236, 35.7036, 35.82475, 
    35.94582, 36.0668, 36.18769, 36.30849, 36.42921, 36.54983, 36.67037, 
    36.79081, 36.91117, 37.03143, 37.15161, 37.27169, 37.39168, 37.51158, 
    37.63138, 37.75109, 37.87072, 37.99024, 38.10967, 38.229, 38.34825, 
    38.46739, 38.58644, 38.70539, 38.82425, 38.94301, 39.06167, 39.18024, 
    39.2987,
  -13.88418, -13.77582, -13.66733, -13.55873, -13.45, -13.34116, -13.23221, 
    -13.12313, -13.01394, -12.90462, -12.79519, -12.68565, -12.57598, 
    -12.4662, -12.3563, -12.24628, -12.13615, -12.0259, -11.91553, -11.80504, 
    -11.69444, -11.58372, -11.47289, -11.36194, -11.25087, -11.13969, 
    -11.02839, -10.91697, -10.80544, -10.6938, -10.58204, -10.47016, 
    -10.35817, -10.24607, -10.13385, -10.02151, -9.909064, -9.796502, 
    -9.683826, -9.571036, -9.458133, -9.345117, -9.231987, -9.118744, 
    -9.005389, -8.891921, -8.778341, -8.664649, -8.550845, -8.436929, 
    -8.322902, -8.208763, -8.094514, -7.980154, -7.865683, -7.751101, 
    -7.63641, -7.521609, -7.406698, -7.291678, -7.176548, -7.06131, 
    -6.945964, -6.830508, -6.714945, -6.599274, -6.483495, -6.367609, 
    -6.251616, -6.135516, -6.01931, -5.902997, -5.786579, -5.670054, 
    -5.553425, -5.43669, -5.319851, -5.202907, -5.085859, -4.968708, 
    -4.851452, -4.734094, -4.616632, -4.499068, -4.381402, -4.263633, 
    -4.145763, -4.027792, -3.90972, -3.791547, -3.673274, -3.554901, 
    -3.436429, -3.317857, -3.199187, -3.080417, -2.96155, -2.842585, 
    -2.723523, -2.604363, -2.485107, -2.365755, -2.246306, -2.126762, 
    -2.007123, -1.887389, -1.767561, -1.647639, -1.527623, -1.407515, 
    -1.287313, -1.167019, -1.046633, -0.9261555, -0.8055869, -0.6849277, 
    -0.5641782, -0.4433389, -0.3224101, -0.2013924, -0.08028615, 0.0409082, 
    0.1621902, 0.2835594, 0.4050153, 0.5265576, 0.6481857, 0.7698992, 
    0.8916976, 1.013581, 1.135547, 1.257598, 1.379731, 1.501947, 1.624246, 
    1.746625, 1.869086, 1.991628, 2.114249, 2.236951, 2.359731, 2.48259, 
    2.605528, 2.728543, 2.851635, 2.974803, 3.098048, 3.221369, 3.344764, 
    3.468235, 3.591779, 3.715396, 3.839087, 3.96285, 4.086685, 4.210591, 
    4.334568, 4.458616, 4.582733, 4.706919, 4.831174, 4.955497, 5.079887, 
    5.204345, 5.328868, 5.453458, 5.578113, 5.702833, 5.827616, 5.952464, 
    6.077374, 6.202346, 6.327381, 6.452476, 6.577632, 6.702848, 6.828124, 
    6.953458, 7.078851, 7.204301, 7.329808, 7.455372, 7.580991, 7.706666, 
    7.832396, 7.958179, 8.084016, 8.209905, 8.335847, 8.46184, 8.587884, 
    8.713978, 8.840121, 8.966314, 9.092555, 9.218844, 9.345181, 9.471563, 
    9.597991, 9.724464, 9.850983, 9.977545, 10.10415, 10.2308, 10.35749, 
    10.48422, 10.61099, 10.7378, 10.86465, 10.99154, 11.11847, 11.24543, 
    11.37243, 11.49947, 11.62654, 11.75365, 11.88079, 12.00797, 12.13518, 
    12.26241, 12.38969, 12.51699, 12.64432, 12.77168, 12.89907, 13.02648, 
    13.15393, 13.2814, 13.4089, 13.53642, 13.66396, 13.79153, 13.91913, 
    14.04674, 14.17438, 14.30204, 14.42972, 14.55741, 14.68513, 14.81287, 
    14.94062, 15.06839, 15.19617, 15.32397, 15.45179, 15.57962, 15.70746, 
    15.83532, 15.96319, 16.09107, 16.21896, 16.34686, 16.47476, 16.60268, 
    16.73061, 16.85854, 16.98647, 17.11442, 17.24237, 17.37032, 17.49828, 
    17.62623, 17.7542, 17.88216, 18.01012, 18.13808, 18.26605, 18.39401, 
    18.52197, 18.64992, 18.77787, 18.90582, 19.03376, 19.1617, 19.28963, 
    19.41755, 19.54547, 19.67338, 19.80128, 19.92916, 20.05704, 20.18491, 
    20.31276, 20.4406, 20.56843, 20.69624, 20.82404, 20.95182, 21.07959, 
    21.20734, 21.33507, 21.46279, 21.59048, 21.71816, 21.84581, 21.97345, 
    22.10106, 22.22865, 22.35621, 22.48376, 22.61127, 22.73877, 22.86623, 
    22.99367, 23.12109, 23.24847, 23.37583, 23.50315, 23.63045, 23.75772, 
    23.88495, 24.01215, 24.13932, 24.26646, 24.39356, 24.52063, 24.64766, 
    24.77465, 24.90161, 25.02853, 25.15542, 25.28226, 25.40907, 25.53583, 
    25.66256, 25.78924, 25.91588, 26.04248, 26.16903, 26.29554, 26.42201, 
    26.54843, 26.67481, 26.80114, 26.92742, 27.05365, 27.17984, 27.30597, 
    27.43206, 27.55809, 27.68408, 27.81001, 27.93589, 28.06172, 28.1875, 
    28.31322, 28.43888, 28.56449, 28.69005, 28.81555, 28.94099, 29.06637, 
    29.1917, 29.31696, 29.44217, 29.56732, 29.6924, 29.81743, 29.94239, 
    30.06729, 30.19213, 30.3169, 30.44161, 30.56625, 30.69083, 30.81535, 
    30.93979, 31.06417, 31.18849, 31.31273, 31.4369, 31.56101, 31.68505, 
    31.80901, 31.93291, 32.05673, 32.18048, 32.30416, 32.42777, 32.5513, 
    32.67476, 32.79815, 32.92145, 33.04469, 33.16784, 33.29092, 33.41393, 
    33.53685, 33.65969, 33.78246, 33.90515, 34.02776, 34.15029, 34.27274, 
    34.39511, 34.51739, 34.6396, 34.76171, 34.88375, 35.00571, 35.12757, 
    35.24936, 35.37106, 35.49268, 35.6142, 35.73565, 35.857, 35.97827, 
    36.09945, 36.22054, 36.34155, 36.46246, 36.58329, 36.70402, 36.82467, 
    36.94522, 37.06568, 37.18605, 37.30633, 37.42652, 37.54662, 37.66661, 
    37.78652, 37.90633, 38.02605, 38.14568, 38.26521, 38.38464, 38.50398, 
    38.62322, 38.74236, 38.86141, 38.98036, 39.09921, 39.21796, 39.33662,
  -13.93741, -13.8289, -13.72028, -13.61153, -13.50267, -13.39369, -13.28459, 
    -13.17537, -13.06603, -12.95658, -12.847, -12.73731, -12.6275, -12.51757, 
    -12.40753, -12.29736, -12.18708, -12.07668, -11.96616, -11.85553, 
    -11.74478, -11.63391, -11.52292, -11.41182, -11.3006, -11.18927, 
    -11.07782, -10.96625, -10.85457, -10.74277, -10.63085, -10.51882, 
    -10.40667, -10.29441, -10.18203, -10.06954, -9.956937, -9.844216, 
    -9.73138, -9.618431, -9.505367, -9.39219, -9.278899, -9.165495, 
    -9.051977, -8.938346, -8.824603, -8.710747, -8.596778, -8.482697, 
    -8.368505, -8.254199, -8.139783, -8.025256, -7.910617, -7.795867, 
    -7.681007, -7.566037, -7.450956, -7.335765, -7.220465, -7.105055, 
    -6.989536, -6.873909, -6.758172, -6.642327, -6.526374, -6.410313, 
    -6.294145, -6.177869, -6.061486, -5.944997, -5.828401, -5.711699, 
    -5.594891, -5.477977, -5.360958, -5.243834, -5.126606, -5.009273, 
    -4.891836, -4.774295, -4.656651, -4.538903, -4.421053, -4.303101, 
    -4.185046, -4.066889, -3.948631, -3.830272, -3.711812, -3.593252, 
    -3.474591, -3.355831, -3.236972, -3.118013, -2.998956, -2.8798, 
    -2.760547, -2.641196, -2.521748, -2.402203, -2.282561, -2.162824, 
    -2.042991, -1.923062, -1.803039, -1.682922, -1.56271, -1.442404, 
    -1.322006, -1.201514, -1.08093, -0.9602543, -0.8394868, -0.718628, 
    -0.5976786, -0.4766389, -0.3555092, -0.2342901, -0.112982, 0.008414708, 
    0.1298995, 0.251472, 0.3731317, 0.4948782, 0.616711, 0.7386296, 
    0.8606337, 0.9827226, 1.104896, 1.227154, 1.349494, 1.471918, 1.594425, 
    1.717013, 1.839684, 1.962435, 2.085267, 2.208179, 2.33117, 2.454241, 
    2.57739, 2.700617, 2.823922, 2.947304, 3.070762, 3.194297, 3.317907, 
    3.441592, 3.565351, 3.689184, 3.813091, 3.93707, 4.061122, 4.185246, 
    4.30944, 4.433706, 4.558042, 4.682446, 4.806921, 4.931463, 5.056074, 
    5.180751, 5.305496, 5.430307, 5.555183, 5.680124, 5.80513, 5.9302, 
    6.055333, 6.180529, 6.305787, 6.431107, 6.556487, 6.681928, 6.807428, 
    6.932988, 7.058606, 7.184282, 7.310016, 7.435806, 7.561653, 7.687555, 
    7.813512, 7.939523, 8.065588, 8.191706, 8.317876, 8.444098, 8.570372, 
    8.696695, 8.82307, 8.949492, 9.075964, 9.202484, 9.329051, 9.455666, 
    9.582325, 9.70903, 9.83578, 9.962575, 10.08941, 10.21629, 10.34322, 
    10.47018, 10.59719, 10.72423, 10.85132, 10.97844, 11.1056, 11.2328, 
    11.36004, 11.48731, 11.61462, 11.74196, 11.86934, 11.99675, 12.12419, 
    12.25167, 12.37918, 12.50671, 12.63428, 12.76188, 12.88951, 13.01716, 
    13.14484, 13.27255, 13.40028, 13.52804, 13.65583, 13.78364, 13.91147, 
    14.03932, 14.1672, 14.29509, 14.42301, 14.55095, 14.6789, 14.80688, 
    14.93487, 15.06288, 15.19091, 15.31895, 15.447, 15.57507, 15.70316, 
    15.83125, 15.95936, 16.08748, 16.21561, 16.34375, 16.4719, 16.60005, 
    16.72822, 16.85639, 16.98457, 17.11275, 17.24094, 17.36913, 17.49733, 
    17.62553, 17.75373, 17.88194, 18.01014, 18.13834, 18.26655, 18.39475, 
    18.52295, 18.65114, 18.77934, 18.90752, 19.03571, 19.16389, 19.29206, 
    19.42022, 19.54838, 19.67652, 19.80466, 19.93279, 20.06091, 20.18901, 
    20.31711, 20.44519, 20.57326, 20.70131, 20.82935, 20.95737, 21.08538, 
    21.21337, 21.34134, 21.46929, 21.59723, 21.72514, 21.85303, 21.9809, 
    22.10876, 22.23658, 22.36439, 22.49217, 22.61992, 22.74765, 22.87536, 
    23.00303, 23.13069, 23.25831, 23.3859, 23.51346, 23.641, 23.7685, 
    23.89597, 24.02341, 24.15081, 24.27818, 24.40552, 24.53283, 24.66009, 
    24.78732, 24.91452, 25.04167, 25.16879, 25.29587, 25.42291, 25.54991, 
    25.67686, 25.80378, 25.93065, 26.05749, 26.18427, 26.31102, 26.43771, 
    26.56437, 26.69097, 26.81753, 26.94404, 27.07051, 27.19692, 27.32329, 
    27.44961, 27.57587, 27.70209, 27.82825, 27.95436, 28.08041, 28.20642, 
    28.33237, 28.45826, 28.5841, 28.70988, 28.8356, 28.96127, 29.08688, 
    29.21243, 29.33792, 29.46335, 29.58872, 29.71403, 29.83928, 29.96447, 
    30.08959, 30.21465, 30.33964, 30.46457, 30.58944, 30.71424, 30.83898, 
    30.96364, 31.08824, 31.21277, 31.33724, 31.46163, 31.58596, 31.71021, 
    31.83439, 31.95851, 32.08255, 32.20651, 32.33041, 32.45423, 32.57798, 
    32.70165, 32.82525, 32.94877, 33.07222, 33.19559, 33.31888, 33.4421, 
    33.56523, 33.68829, 33.81127, 33.93417, 34.05699, 34.17973, 34.30238, 
    34.42496, 34.54745, 34.66986, 34.79219, 34.91444, 35.03659, 35.15867, 
    35.28066, 35.40257, 35.52439, 35.64612, 35.76777, 35.88932, 36.0108, 
    36.13218, 36.25347, 36.37468, 36.49579, 36.61682, 36.73775, 36.8586, 
    36.97935, 37.10001, 37.22058, 37.34106, 37.46144, 37.58173, 37.70193, 
    37.82203, 37.94204, 38.06195, 38.18177, 38.30149, 38.42112, 38.54065, 
    38.66008, 38.77942, 38.89865, 39.0178, 39.13684, 39.25578, 39.37462,
  -13.99074, -13.88209, -13.77333, -13.66444, -13.55544, -13.44631, 
    -13.33707, -13.22771, -13.11823, -13.00863, -12.89891, -12.78907, 
    -12.67912, -12.56904, -12.45885, -12.34854, -12.23811, -12.12756, 
    -12.0169, -11.90611, -11.79521, -11.6842, -11.57306, -11.46181, 
    -11.35044, -11.23895, -11.12734, -11.01562, -10.90379, -10.79183, 
    -10.67976, -10.56758, -10.45527, -10.34285, -10.23032, -10.11767, 
    -10.00491, -9.892027, -9.779033, -9.665923, -9.552699, -9.439362, 
    -9.325909, -9.212342, -9.098662, -8.984868, -8.870961, -8.756941, 
    -8.642807, -8.528561, -8.414203, -8.299731, -8.185148, -8.070454, 
    -7.955647, -7.840729, -7.725699, -7.610559, -7.495308, -7.379947, 
    -7.264475, -7.148894, -7.033203, -6.917402, -6.801492, -6.685473, 
    -6.569346, -6.45311, -6.336766, -6.220315, -6.103755, -5.987089, 
    -5.870315, -5.753435, -5.636448, -5.519355, -5.402156, -5.284852, 
    -5.167442, -5.049928, -4.932309, -4.814586, -4.696759, -4.578828, 
    -4.460793, -4.342657, -4.224417, -4.106074, -3.98763, -3.869085, 
    -3.750437, -3.63169, -3.512841, -3.393892, -3.274843, -3.155695, 
    -3.036447, -2.917101, -2.797656, -2.678113, -2.558473, -2.438735, 
    -2.3189, -2.198969, -2.078942, -1.958818, -1.8386, -1.718286, -1.597878, 
    -1.477376, -1.35678, -1.23609, -1.115308, -0.9944334, -0.8734666, 
    -0.752408, -0.6312582, -0.5100177, -0.3886868, -0.2672659, -0.1457556, 
    -0.02415619, 0.0975318, 0.2193079, 0.3411718, 0.4631229, 0.5851607, 
    0.7072849, 0.829495, 0.9517905, 1.074171, 1.196636, 1.319184, 1.441817, 
    1.564532, 1.68733, 1.810209, 1.933171, 2.056213, 2.179336, 2.302539, 
    2.425821, 2.549183, 2.672623, 2.796141, 2.919736, 3.043409, 3.167158, 
    3.290982, 3.414883, 3.538858, 3.662907, 3.78703, 3.911227, 4.035496, 
    4.159837, 4.28425, 4.408734, 4.533288, 4.657913, 4.782607, 4.907369, 
    5.0322, 5.157099, 5.282064, 5.407097, 5.532195, 5.657359, 5.782588, 
    5.90788, 6.033237, 6.158657, 6.284139, 6.409683, 6.535288, 6.660954, 
    6.78668, 6.912466, 7.03831, 7.164213, 7.290174, 7.416191, 7.542265, 
    7.668395, 7.79458, 7.92082, 8.047113, 8.17346, 8.29986, 8.426311, 
    8.552815, 8.679369, 8.805974, 8.932628, 9.059331, 9.186082, 9.312881, 
    9.439726, 9.566618, 9.693556, 9.820539, 9.947566, 10.07464, 10.20175, 
    10.32891, 10.45611, 10.58335, 10.71063, 10.83794, 10.9653, 11.0927, 
    11.22014, 11.34761, 11.47512, 11.60266, 11.73024, 11.85785, 11.9855, 
    12.11318, 12.24089, 12.36864, 12.49641, 12.62422, 12.75205, 12.87992, 
    13.00781, 13.13573, 13.26368, 13.39165, 13.51965, 13.64767, 13.77572, 
    13.90379, 14.03188, 14.16, 14.28813, 14.41629, 14.54447, 14.67266, 
    14.80088, 14.92911, 15.05736, 15.18562, 15.31391, 15.4422, 15.57051, 
    15.69884, 15.82717, 15.95552, 16.08388, 16.21225, 16.34063, 16.46902, 
    16.59742, 16.72583, 16.85424, 16.98266, 17.11108, 17.23951, 17.36795, 
    17.49639, 17.62483, 17.75327, 17.88171, 18.01016, 18.1386, 18.26705, 
    18.39549, 18.52393, 18.65237, 18.7808, 18.90923, 19.03765, 19.16607, 
    19.29449, 19.42289, 19.55129, 19.67968, 19.80806, 19.93642, 20.06478, 
    20.19313, 20.32146, 20.44979, 20.57809, 20.70639, 20.83467, 20.96293, 
    21.09118, 21.21941, 21.34762, 21.47581, 21.60398, 21.73214, 21.86027, 
    21.98838, 22.11647, 22.24454, 22.37258, 22.5006, 22.6286, 22.75656, 
    22.88451, 23.01242, 23.14031, 23.26817, 23.396, 23.5238, 23.65157, 
    23.77931, 23.90702, 24.03469, 24.16234, 24.28994, 24.41752, 24.54506, 
    24.67256, 24.80003, 24.92745, 25.05485, 25.1822, 25.30951, 25.43678, 
    25.56402, 25.69121, 25.81836, 25.94547, 26.07253, 26.19955, 26.32653, 
    26.45346, 26.58034, 26.70718, 26.83397, 26.96071, 27.08741, 27.21406, 
    27.34065, 27.4672, 27.59369, 27.72014, 27.84653, 27.97287, 28.09915, 
    28.22538, 28.35156, 28.47768, 28.60375, 28.72976, 28.85571, 28.9816, 
    29.10744, 29.23321, 29.35893, 29.48458, 29.61018, 29.73571, 29.86119, 
    29.9866, 30.11194, 30.23723, 30.36244, 30.4876, 30.61269, 30.73771, 
    30.86266, 30.98755, 31.11237, 31.23712, 31.3618, 31.48642, 31.61096, 
    31.73544, 31.85984, 31.98417, 32.10843, 32.23261, 32.35672, 32.48076, 
    32.60472, 32.72861, 32.85242, 32.97616, 33.09982, 33.2234, 33.34691, 
    33.47034, 33.59369, 33.71696, 33.84015, 33.96326, 34.08628, 34.20923, 
    34.3321, 34.45488, 34.57759, 34.70021, 34.82274, 34.94519, 35.06756, 
    35.18984, 35.31204, 35.43415, 35.55618, 35.67811, 35.79996, 35.92172, 
    36.0434, 36.16498, 36.28648, 36.40789, 36.5292, 36.65043, 36.77156, 
    36.89261, 37.01356, 37.13442, 37.25519, 37.37586, 37.49644, 37.61693, 
    37.73732, 37.85762, 37.97783, 38.09793, 38.21795, 38.33786, 38.45768, 
    38.5774, 38.69703, 38.81656, 38.93599, 39.05532, 39.17455, 39.29368, 
    39.41272,
  -14.04416, -13.93538, -13.82647, -13.71745, -13.6083, -13.49904, -13.38965, 
    -13.28015, -13.17053, -13.06078, -12.95092, -12.84094, -12.73084, 
    -12.62062, -12.51028, -12.39982, -12.28924, -12.17855, -12.06773, 
    -11.9568, -11.84575, -11.73458, -11.62329, -11.51189, -11.40037, 
    -11.28873, -11.17697, -11.0651, -10.9531, -10.841, -10.72877, -10.61643, 
    -10.50397, -10.3914, -10.2787, -10.1659, -10.05297, -9.939937, -9.826782, 
    -9.713513, -9.600129, -9.486629, -9.373015, -9.259287, -9.145444, 
    -9.031487, -8.917416, -8.803231, -8.688933, -8.574521, -8.459997, 
    -8.34536, -8.230609, -8.115746, -8.000772, -7.885685, -7.770487, 
    -7.655177, -7.539756, -7.424223, -7.308581, -7.192827, -7.076963, 
    -6.96099, -6.844906, -6.728714, -6.612411, -6.496, -6.379481, -6.262853, 
    -6.146117, -6.029273, -5.912321, -5.795262, -5.678097, -5.560824, 
    -5.443446, -5.325961, -5.20837, -5.090674, -4.972873, -4.854967, 
    -4.736957, -4.618842, -4.500624, -4.382302, -4.263876, -4.145349, 
    -4.026718, -3.907985, -3.789151, -3.670215, -3.551178, -3.43204, 
    -3.312801, -3.193463, -3.074025, -2.954488, -2.834851, -2.715116, 
    -2.595283, -2.475352, -2.355324, -2.235198, -2.114976, -1.994658, 
    -1.874243, -1.753734, -1.633129, -1.512429, -1.391636, -1.270748, 
    -1.149767, -1.028693, -0.9075267, -0.7862681, -0.6649176, -0.543476, 
    -0.4219434, -0.3003204, -0.1786075, -0.05680501, 0.06508655, 0.1870667, 
    0.3091351, 0.4312912, 0.5535345, 0.6758646, 0.7982811, 0.9207833, 
    1.043371, 1.166044, 1.288801, 1.411642, 1.534566, 1.657573, 1.780663, 
    1.903835, 2.027088, 2.150423, 2.273838, 2.397332, 2.520906, 2.64456, 
    2.768291, 2.892101, 3.015988, 3.139951, 3.263992, 3.388108, 3.512299, 
    3.636564, 3.760905, 3.885319, 4.009805, 4.134365, 4.258996, 4.383699, 
    4.508473, 4.633317, 4.758232, 4.883215, 5.008266, 5.133387, 5.258574, 
    5.383829, 5.50915, 5.634536, 5.759988, 5.885504, 6.011085, 6.136729, 
    6.262435, 6.388205, 6.514035, 6.639927, 6.765879, 6.891891, 7.017962, 
    7.144092, 7.27028, 7.396525, 7.522827, 7.649185, 7.775599, 7.902068, 
    8.028591, 8.155168, 8.281797, 8.40848, 8.535213, 8.661998, 8.788834, 
    8.915719, 9.042654, 9.169637, 9.296668, 9.423746, 9.550871, 9.678041, 
    9.805258, 9.932519, 10.05982, 10.18717, 10.31456, 10.442, 10.56947, 
    10.69698, 10.82454, 10.95213, 11.07977, 11.20744, 11.33515, 11.46289, 
    11.59067, 11.71849, 11.84634, 11.97422, 12.10214, 12.23009, 12.35807, 
    12.48609, 12.61413, 12.7422, 12.87031, 12.99844, 13.1266, 13.25478, 
    13.38299, 13.51123, 13.63949, 13.76778, 13.89609, 14.02442, 14.15278, 
    14.28115, 14.40955, 14.53797, 14.6664, 14.79486, 14.92333, 15.05182, 
    15.18033, 15.30885, 15.43739, 15.56594, 15.6945, 15.82308, 15.95167, 
    16.08027, 16.20889, 16.33751, 16.46614, 16.59478, 16.72343, 16.85208, 
    16.98074, 17.10941, 17.23808, 17.36676, 17.49544, 17.62412, 17.75281, 
    17.88149, 18.01018, 18.13886, 18.26755, 18.39623, 18.52492, 18.6536, 
    18.78227, 18.91094, 19.03961, 19.16827, 19.29692, 19.42557, 19.55421, 
    19.68284, 19.81146, 19.94007, 20.06867, 20.19726, 20.32583, 20.4544, 
    20.58294, 20.71148, 20.84, 20.9685, 21.09699, 21.22546, 21.35391, 
    21.48235, 21.61076, 21.73915, 21.86753, 21.99588, 22.12421, 22.25252, 
    22.3808, 22.50906, 22.63729, 22.7655, 22.89368, 23.02183, 23.14996, 
    23.27806, 23.40613, 23.53417, 23.66217, 23.79015, 23.9181, 24.04601, 
    24.17389, 24.30173, 24.42954, 24.55732, 24.68506, 24.81276, 24.94043, 
    25.06805, 25.19564, 25.32319, 25.4507, 25.57817, 25.70559, 25.83298, 
    25.96032, 26.08761, 26.21487, 26.34208, 26.46924, 26.59636, 26.72343, 
    26.85045, 26.97743, 27.10435, 27.23123, 27.35806, 27.48484, 27.61156, 
    27.73824, 27.86486, 27.99143, 28.11794, 28.2444, 28.37081, 28.49716, 
    28.62345, 28.74969, 28.87586, 29.00198, 29.12805, 29.25405, 29.37999, 
    29.50587, 29.63169, 29.75745, 29.88315, 30.00879, 30.13436, 30.25986, 
    30.3853, 30.51068, 30.63599, 30.76123, 30.88641, 31.01152, 31.13656, 
    31.26153, 31.38644, 31.51127, 31.63603, 31.76072, 31.88534, 32.00989, 
    32.13437, 32.25877, 32.3831, 32.50735, 32.63153, 32.75563, 32.87966, 
    33.00362, 33.12749, 33.25129, 33.375, 33.49865, 33.62221, 33.74569, 
    33.86909, 33.99241, 34.11565, 34.23881, 34.36189, 34.48489, 34.6078, 
    34.73062, 34.85337, 34.97602, 35.0986, 35.22109, 35.34349, 35.46581, 
    35.58804, 35.71018, 35.83223, 35.9542, 36.07608, 36.19787, 36.31956, 
    36.44117, 36.56269, 36.68412, 36.80545, 36.9267, 37.04785, 37.16891, 
    37.28988, 37.41075, 37.53153, 37.65221, 37.7728, 37.8933, 38.01369, 
    38.134, 38.25421, 38.37432, 38.49433, 38.61425, 38.73406, 38.85378, 
    38.9734, 39.09293, 39.21235, 39.33167, 39.45089,
  -14.09769, -13.98877, -13.87972, -13.77056, -13.66127, -13.55186, 
    -13.44234, -13.33269, -13.22292, -13.11304, -13.00303, -12.8929, 
    -12.78265, -12.67229, -12.5618, -12.4512, -12.34047, -12.22963, 
    -12.11867, -12.00759, -11.89639, -11.78507, -11.67363, -11.56207, 
    -11.4504, -11.33861, -11.2267, -11.11467, -11.00252, -10.89026, 
    -10.77788, -10.66538, -10.55277, -10.44004, -10.32719, -10.21422, 
    -10.10114, -9.987945, -9.874631, -9.761201, -9.647656, -9.533996, 
    -9.42022, -9.30633, -9.192324, -9.078203, -8.963968, -8.849619, 
    -8.735156, -8.620579, -8.505888, -8.391084, -8.276167, -8.161137, 
    -8.045994, -7.930738, -7.81537, -7.699891, -7.584299, -7.468596, 
    -7.352781, -7.236856, -7.120819, -7.004673, -6.888415, -6.772048, 
    -6.655571, -6.538985, -6.422289, -6.305485, -6.188571, -6.07155, 
    -5.954421, -5.837183, -5.719838, -5.602386, -5.484827, -5.367161, 
    -5.24939, -5.131512, -5.013528, -4.895439, -4.777246, -4.658947, 
    -4.540544, -4.422037, -4.303426, -4.184712, -4.065895, -3.946975, 
    -3.827953, -3.708828, -3.589602, -3.470275, -3.350847, -3.231318, 
    -3.111689, -2.991961, -2.872132, -2.752205, -2.632179, -2.512054, 
    -2.391832, -2.271512, -2.151095, -2.030581, -1.909971, -1.789265, 
    -1.668463, -1.547566, -1.426574, -1.305488, -1.184308, -1.063035, 
    -0.9416679, -0.8202087, -0.6986573, -0.5770141, -0.4552795, -0.3334541, 
    -0.2115382, -0.08953223, 0.03256327, 0.1547479, 0.2770211, 0.3993826, 
    0.5218318, 0.6443682, 0.7669914, 0.889701, 1.012496, 1.135377, 1.258343, 
    1.381393, 1.504527, 1.627744, 1.751045, 1.874427, 1.997892, 2.121438, 
    2.245065, 2.368773, 2.49256, 2.616427, 2.740373, 2.864397, 2.988498, 
    3.112678, 3.236933, 3.361266, 3.485673, 3.610156, 3.734714, 3.859346, 
    3.984051, 4.108829, 4.23368, 4.358602, 4.483596, 4.60866, 4.733795, 
    4.858999, 4.984272, 5.109614, 5.235024, 5.360501, 5.486045, 5.611655, 
    5.73733, 5.863071, 5.988876, 6.114745, 6.240677, 6.366671, 6.492728, 
    6.618845, 6.745024, 6.871264, 6.997562, 7.123919, 7.250335, 7.376809, 
    7.503339, 7.629927, 7.756569, 7.883268, 8.01002, 8.136827, 8.263688, 
    8.3906, 8.517566, 8.644582, 8.771649, 8.898767, 9.025933, 9.153149, 
    9.280413, 9.407724, 9.535083, 9.662487, 9.789937, 9.917432, 10.04497, 
    10.17255, 10.30018, 10.42785, 10.55556, 10.68331, 10.8111, 10.93893, 
    11.0668, 11.19471, 11.32265, 11.45063, 11.57865, 11.7067, 11.83479, 
    11.96291, 12.09107, 12.21926, 12.34748, 12.47573, 12.60401, 12.73233, 
    12.86067, 12.98904, 13.11744, 13.24586, 13.37431, 13.50279, 13.63129, 
    13.75982, 13.88837, 14.01694, 14.14554, 14.27416, 14.40279, 14.53145, 
    14.66013, 14.78883, 14.91754, 15.04627, 15.17502, 15.30378, 15.43256, 
    15.56135, 15.69016, 15.81898, 15.94781, 16.07666, 16.20551, 16.33438, 
    16.46325, 16.59213, 16.72102, 16.84992, 16.97882, 17.10773, 17.23665, 
    17.36556, 17.49449, 17.62341, 17.75234, 17.88127, 18.0102, 18.13913, 
    18.26805, 18.39698, 18.52591, 18.65483, 18.78375, 18.91266, 19.04157, 
    19.17047, 19.29937, 19.42826, 19.55714, 19.68601, 19.81487, 19.94373, 
    20.07257, 20.2014, 20.33022, 20.45902, 20.58781, 20.71659, 20.84535, 
    20.97409, 21.10282, 21.23153, 21.36023, 21.4889, 21.61756, 21.74619, 
    21.8748, 22.0034, 22.13197, 22.26051, 22.38904, 22.51753, 22.64601, 
    22.77446, 22.90288, 23.03127, 23.15964, 23.28797, 23.41628, 23.54456, 
    23.67281, 23.80102, 23.9292, 24.05736, 24.18547, 24.31355, 24.4416, 
    24.56961, 24.69759, 24.82553, 24.95343, 25.0813, 25.20912, 25.3369, 
    25.46465, 25.59235, 25.72001, 25.84763, 25.97521, 26.10274, 26.23023, 
    26.35767, 26.48507, 26.61242, 26.73972, 26.86698, 26.99419, 27.12135, 
    27.24846, 27.37551, 27.50252, 27.62948, 27.75638, 27.88323, 28.01003, 
    28.13678, 28.26347, 28.3901, 28.51668, 28.6432, 28.76967, 28.89607, 
    29.02242, 29.14871, 29.27494, 29.40111, 29.52722, 29.65326, 29.77925, 
    29.90517, 30.03103, 30.15682, 30.28255, 30.40822, 30.53382, 30.65935, 
    30.78482, 30.91022, 31.03555, 31.16081, 31.286, 31.41113, 31.53618, 
    31.66116, 31.78608, 31.91091, 32.03568, 32.16037, 32.28499, 32.40954, 
    32.53401, 32.65841, 32.78273, 32.90697, 33.03114, 33.15523, 33.27924, 
    33.40317, 33.52703, 33.6508, 33.77449, 33.89811, 34.02164, 34.1451, 
    34.26847, 34.39175, 34.51496, 34.63808, 34.76111, 34.88407, 35.00694, 
    35.12971, 35.25241, 35.37502, 35.49754, 35.61998, 35.74232, 35.86459, 
    35.98676, 36.10884, 36.23083, 36.35273, 36.47454, 36.59626, 36.71789, 
    36.83943, 36.96087, 37.08223, 37.20348, 37.32465, 37.44572, 37.5667, 
    37.68758, 37.80836, 37.92905, 38.04965, 38.17015, 38.29055, 38.41085, 
    38.53106, 38.65117, 38.77118, 38.89109, 39.01091, 39.13062, 39.25023, 
    39.36975, 39.48916,
  -14.15132, -14.04226, -13.93307, -13.82376, -13.71434, -13.60479, 
    -13.49512, -13.38533, -13.27542, -13.16539, -13.05524, -12.94497, 
    -12.83457, -12.72406, -12.61343, -12.50268, -12.39181, -12.28081, 
    -12.1697, -12.05847, -11.94712, -11.83565, -11.72406, -11.61236, 
    -11.50053, -11.38859, -11.27652, -11.16434, -11.05204, -10.93962, 
    -10.82709, -10.71444, -10.60166, -10.48878, -10.37577, -10.26265, 
    -10.14941, -10.03605, -9.922578, -9.808989, -9.695283, -9.581461, 
    -9.467524, -9.35347, -9.239302, -9.125018, -9.010619, -8.896105, 
    -8.781477, -8.666734, -8.551877, -8.436906, -8.321821, -8.206623, 
    -8.091312, -7.975888, -7.86035, -7.7447, -7.628938, -7.513064, -7.397078, 
    -7.28098, -7.164771, -7.04845, -6.932019, -6.815477, -6.698825, 
    -6.582064, -6.465192, -6.348211, -6.23112, -6.113921, -5.996613, 
    -5.879197, -5.761672, -5.644041, -5.526301, -5.408454, -5.290501, 
    -5.172441, -5.054275, -4.936003, -4.817626, -4.699142, -4.580554, 
    -4.461862, -4.343066, -4.224165, -4.105161, -3.986054, -3.866843, 
    -3.747531, -3.628116, -3.508599, -3.388981, -3.269261, -3.149441, 
    -3.029521, -2.9095, -2.78938, -2.669161, -2.548842, -2.428426, -2.307911, 
    -2.187299, -2.066589, -1.945782, -1.824879, -1.70388, -1.582785, 
    -1.461595, -1.34031, -1.218931, -1.097458, -0.9758906, -0.8542305, 
    -0.7324777, -0.6106326, -0.4886957, -0.3666674, -0.2445481, -0.1223384, 
    -3.855618e-05, 0.1223508, 0.2448294, 0.3673966, 0.490052, 0.6127952, 
    0.7356256, 0.8585429, 0.9815464, 1.104636, 1.227811, 1.35107, 1.474414, 
    1.597842, 1.721353, 1.844947, 1.968624, 2.092382, 2.216222, 2.340143, 
    2.464144, 2.588225, 2.712385, 2.836624, 2.960941, 3.085336, 3.209808, 
    3.334357, 3.458982, 3.583682, 3.708457, 3.833308, 3.958231, 4.083229, 
    4.208299, 4.333441, 4.458655, 4.583941, 4.709297, 4.834723, 4.960218, 
    5.085782, 5.211414, 5.337114, 5.462882, 5.588716, 5.714615, 5.84058, 
    5.96661, 6.092705, 6.218862, 6.345083, 6.471366, 6.597711, 6.724116, 
    6.850583, 6.977109, 7.103694, 7.230339, 7.357041, 7.483801, 7.610618, 
    7.737491, 7.864419, 7.991402, 8.11844, 8.245531, 8.372675, 8.499872, 
    8.62712, 8.754419, 8.881769, 9.00917, 9.136618, 9.264115, 9.391661, 
    9.519253, 9.646892, 9.774576, 9.902306, 10.03008, 10.1579, 10.28576, 
    10.41366, 10.54161, 10.6696, 10.79762, 10.92569, 11.0538, 11.18194, 
    11.31012, 11.43834, 11.5666, 11.69489, 11.82322, 11.95158, 12.07997, 
    12.2084, 12.33686, 12.46535, 12.59387, 12.72242, 12.851, 12.97961, 
    13.10825, 13.23692, 13.36561, 13.49433, 13.62307, 13.75184, 13.88063, 
    14.00944, 14.13828, 14.26714, 14.39602, 14.52492, 14.65384, 14.78278, 
    14.91173, 15.04071, 15.1697, 15.2987, 15.42772, 15.55676, 15.68581, 
    15.81487, 15.94394, 16.07303, 16.20213, 16.33123, 16.46035, 16.58948, 
    16.71861, 16.84775, 16.9769, 17.10605, 17.23521, 17.36437, 17.49353, 
    17.6227, 17.75187, 17.88104, 18.01022, 18.13939, 18.26856, 18.39773, 
    18.5269, 18.65606, 18.78522, 18.91438, 19.04353, 19.17268, 19.30182, 
    19.43095, 19.56007, 19.68919, 19.81829, 19.94739, 20.07648, 20.20555, 
    20.33461, 20.46365, 20.59269, 20.72171, 20.85071, 20.9797, 21.10867, 
    21.23762, 21.36656, 21.49547, 21.62437, 21.75324, 21.8821, 22.01093, 
    22.13974, 22.26853, 22.39729, 22.52604, 22.65475, 22.78344, 22.9121, 
    23.04073, 23.16934, 23.29791, 23.42646, 23.55498, 23.68346, 23.81192, 
    23.94034, 24.06873, 24.19709, 24.32541, 24.45369, 24.58194, 24.71016, 
    24.83833, 24.96647, 25.09457, 25.22263, 25.35065, 25.47863, 25.60657, 
    25.73447, 25.86232, 25.99014, 26.1179, 26.24562, 26.3733, 26.50093, 
    26.62852, 26.75606, 26.88354, 27.01099, 27.13838, 27.26572, 27.39301, 
    27.52025, 27.64744, 27.77458, 27.90166, 28.02869, 28.15566, 28.28258, 
    28.40945, 28.53625, 28.663, 28.7897, 28.91633, 29.04291, 29.16943, 
    29.29588, 29.42228, 29.54861, 29.67489, 29.8011, 29.92725, 30.05333, 
    30.17935, 30.3053, 30.43119, 30.55702, 30.68277, 30.80846, 30.93409, 
    31.05964, 31.18512, 31.31054, 31.43588, 31.56116, 31.68636, 31.81149, 
    31.93655, 32.06153, 32.18645, 32.31129, 32.43605, 32.56074, 32.68535, 
    32.80989, 32.93435, 33.05873, 33.18303, 33.30726, 33.43141, 33.55548, 
    33.67947, 33.80337, 33.9272, 34.05095, 34.17461, 34.29819, 34.42169, 
    34.5451, 34.66843, 34.79168, 34.91484, 35.03792, 35.16091, 35.28381, 
    35.40663, 35.52936, 35.652, 35.77455, 35.89701, 36.01939, 36.14168, 
    36.26387, 36.38597, 36.50799, 36.62991, 36.75174, 36.87348, 36.99513, 
    37.11668, 37.23814, 37.3595, 37.48077, 37.60195, 37.72303, 37.84401, 
    37.9649, 38.08569, 38.20638, 38.32698, 38.44748, 38.56788, 38.68818, 
    38.80839, 38.92849, 39.0485, 39.1684, 39.2882, 39.40791, 39.52751,
  -14.20505, -14.09585, -13.98652, -13.87708, -13.76751, -13.65782, 
    -13.54801, -13.43807, -13.32802, -13.21784, -13.10755, -12.99713, 
    -12.88659, -12.77594, -12.66516, -12.55426, -12.44324, -12.3321, 
    -12.22084, -12.10946, -11.99796, -11.88634, -11.7746, -11.66274, 
    -11.55076, -11.43867, -11.32645, -11.21412, -11.10166, -10.98909, 
    -10.8764, -10.76359, -10.65066, -10.53762, -10.42445, -10.31117, 
    -10.19777, -10.08426, -9.970625, -9.856875, -9.743009, -9.629025, 
    -9.514926, -9.40071, -9.286379, -9.171931, -9.057368, -8.94269, 
    -8.827896, -8.712988, -8.597964, -8.482826, -8.367575, -8.252208, 
    -8.136728, -8.021134, -7.905427, -7.789607, -7.673674, -7.557628, 
    -7.44147, -7.3252, -7.208818, -7.092324, -6.975719, -6.859003, -6.742175, 
    -6.625237, -6.50819, -6.391031, -6.273764, -6.156386, -6.0389, -5.921305, 
    -5.803601, -5.685789, -5.567868, -5.449841, -5.331705, -5.213463, 
    -5.095114, -4.976658, -4.858097, -4.739429, -4.620656, -4.501779, 
    -4.382796, -4.263709, -4.144517, -4.025222, -3.905824, -3.786322, 
    -3.666718, -3.547011, -3.427203, -3.307292, -3.187281, -3.067168, 
    -2.946955, -2.826642, -2.706229, -2.585717, -2.465106, -2.344396, 
    -2.223588, -2.102682, -1.981679, -1.860578, -1.739382, -1.618088, 
    -1.4967, -1.375216, -1.253636, -1.131963, -1.010195, -0.8883339, 
    -0.7663794, -0.6443321, -0.5221924, -0.3999608, -0.2776379, -0.1552239, 
    -0.03271941, 0.08987517, 0.2125594, 0.3353328, 0.4581948, 0.581145, 
    0.7041831, 0.8273084, 0.9505205, 1.073819, 1.197203, 1.320673, 1.444227, 
    1.567866, 1.691588, 1.815394, 1.939283, 2.063254, 2.187307, 2.311441, 
    2.435657, 2.559952, 2.684327, 2.808781, 2.933314, 3.057925, 3.182614, 
    3.30738, 3.432222, 3.557141, 3.682135, 3.807204, 3.932347, 4.057564, 
    4.182854, 4.308217, 4.433652, 4.559158, 4.684736, 4.810384, 4.936101, 
    5.061889, 5.187744, 5.313668, 5.439659, 5.565718, 5.691842, 5.818032, 
    5.944288, 6.070608, 6.196991, 6.323439, 6.449949, 6.576521, 6.703154, 
    6.829849, 6.956604, 7.083417, 7.210291, 7.337223, 7.464212, 7.591259, 
    7.718362, 7.845521, 7.972735, 8.100004, 8.227327, 8.354703, 8.482132, 
    8.609613, 8.737145, 8.864728, 8.992361, 9.120044, 9.247775, 9.375554, 
    9.503381, 9.631255, 9.759174, 9.887139, 10.01515, 10.1432, 10.2713, 
    10.39944, 10.52762, 10.65585, 10.78411, 10.91242, 11.04076, 11.16914, 
    11.29756, 11.42602, 11.55451, 11.68304, 11.81161, 11.94021, 12.06884, 
    12.19751, 12.32621, 12.45494, 12.5837, 12.71249, 12.84131, 12.97017, 
    13.09904, 13.22795, 13.35688, 13.48584, 13.61483, 13.74384, 13.87287, 
    14.00193, 14.131, 14.26011, 14.38923, 14.51837, 14.64753, 14.77671, 
    14.90591, 15.03512, 15.16436, 15.29361, 15.42287, 15.55215, 15.68144, 
    15.81075, 15.94006, 16.06939, 16.19873, 16.32808, 16.45745, 16.58681, 
    16.71619, 16.84557, 16.97496, 17.10436, 17.23376, 17.36317, 17.49258, 
    17.62199, 17.7514, 17.88082, 18.01024, 18.13965, 18.26907, 18.39848, 
    18.52789, 18.6573, 18.78671, 18.91611, 19.0455, 19.17489, 19.30428, 
    19.43365, 19.56302, 19.69238, 19.82173, 19.95107, 20.08039, 20.20971, 
    20.33901, 20.4683, 20.59758, 20.72684, 20.85609, 20.98532, 21.11453, 
    21.24372, 21.3729, 21.50206, 21.6312, 21.76032, 21.88942, 22.01849, 
    22.14754, 22.27657, 22.40558, 22.53456, 22.66351, 22.79244, 22.92134, 
    23.05022, 23.17907, 23.30788, 23.43667, 23.56543, 23.69415, 23.82285, 
    23.95151, 24.08014, 24.20873, 24.33729, 24.46581, 24.5943, 24.72276, 
    24.85117, 24.97955, 25.10788, 25.23618, 25.36444, 25.49266, 25.62083, 
    25.74896, 25.87706, 26.0051, 26.13311, 26.26106, 26.38898, 26.51684, 
    26.64466, 26.77243, 26.90016, 27.02783, 27.15546, 27.28303, 27.41056, 
    27.53803, 27.66545, 27.79282, 27.92013, 28.04739, 28.1746, 28.30175, 
    28.42884, 28.55588, 28.68286, 28.80978, 28.93665, 29.06345, 29.1902, 
    29.31688, 29.4435, 29.57007, 29.69657, 29.823, 29.94938, 30.07569, 
    30.20193, 30.32811, 30.45423, 30.58027, 30.70625, 30.83217, 30.95801, 
    31.08379, 31.2095, 31.33513, 31.4607, 31.58619, 31.71162, 31.83697, 
    31.96225, 32.08746, 32.21259, 32.33764, 32.46262, 32.58753, 32.71236, 
    32.83712, 32.96179, 33.08639, 33.21091, 33.33535, 33.45972, 33.584, 
    33.7082, 33.83232, 33.95636, 34.08032, 34.2042, 34.32799, 34.4517, 
    34.57532, 34.69886, 34.82232, 34.94569, 35.06898, 35.19217, 35.31528, 
    35.43831, 35.56124, 35.68409, 35.80685, 35.92952, 36.0521, 36.17459, 
    36.29699, 36.4193, 36.54152, 36.66364, 36.78568, 36.90762, 37.02946, 
    37.15121, 37.27287, 37.39444, 37.51591, 37.63728, 37.75856, 37.87974, 
    38.00083, 38.12181, 38.2427, 38.3635, 38.48419, 38.60479, 38.72528, 
    38.84568, 38.96598, 39.08617, 39.20627, 39.32627, 39.44616, 39.56595,
  -14.25888, -14.14954, -14.04008, -13.93049, -13.82078, -13.71095, 
    -13.60099, -13.49092, -13.38072, -13.2704, -13.15996, -13.0494, 
    -12.93872, -12.82791, -12.71699, -12.60594, -12.49477, -12.38349, 
    -12.27208, -12.16055, -12.0489, -11.93713, -11.82524, -11.71323, 
    -11.6011, -11.48885, -11.37648, -11.26399, -11.15138, -11.03866, 
    -10.92581, -10.81284, -10.69976, -10.58656, -10.47324, -10.3598, 
    -10.24624, -10.13256, -10.01877, -9.904862, -9.790834, -9.67669, 
    -9.562428, -9.44805, -9.333555, -9.218944, -9.104217, -8.989373, 
    -8.874414, -8.759339, -8.64415, -8.528845, -8.413425, -8.297891, 
    -8.182242, -8.066479, -7.950602, -7.834611, -7.718508, -7.60229, 
    -7.48596, -7.369517, -7.252962, -7.136294, -7.019515, -6.902624, 
    -6.785621, -6.668507, -6.551282, -6.433948, -6.316502, -6.198946, 
    -6.081281, -5.963507, -5.845623, -5.727631, -5.609529, -5.49132, 
    -5.373003, -5.254578, -5.136045, -5.017406, -4.898661, -4.779809, 
    -4.660851, -4.541787, -4.422617, -4.303343, -4.183965, -4.064481, 
    -3.944894, -3.825204, -3.70541, -3.585513, -3.465514, -3.345412, 
    -3.225209, -3.104904, -2.984498, -2.863992, -2.743385, -2.622679, 
    -2.501872, -2.380967, -2.259963, -2.138861, -2.01766, -1.896363, 
    -1.774968, -1.653476, -1.531888, -1.410204, -1.288425, -1.166551, 
    -1.044582, -0.9225194, -0.8003628, -0.6781129, -0.5557702, -0.433335, 
    -0.3108079, -0.1881894, -0.06547982, 0.05732033, 0.1802106, 0.3031905, 
    0.4262596, 0.5494174, 0.6726634, 0.7959971, 0.9194182, 1.042926, 1.16652, 
    1.2902, 1.413965, 1.537815, 1.66175, 1.785768, 1.909869, 2.034054, 
    2.15832, 2.282668, 2.407098, 2.531608, 2.656199, 2.780869, 2.905618, 
    3.030446, 3.155352, 3.280335, 3.405396, 3.530533, 3.655746, 3.781034, 
    3.906396, 4.031834, 4.157344, 4.282928, 4.408585, 4.534313, 4.660112, 
    4.785983, 4.911923, 5.037934, 5.164013, 5.290162, 5.416377, 5.54266, 
    5.66901, 5.795426, 5.921907, 6.048454, 6.175065, 6.301739, 6.428476, 
    6.555276, 6.682138, 6.809061, 6.936044, 7.063088, 7.190191, 7.317352, 
    7.444572, 7.571849, 7.699183, 7.826574, 7.95402, 8.08152, 8.209076, 
    8.336684, 8.464346, 8.59206, 8.719826, 8.847642, 8.97551, 9.103426, 
    9.231392, 9.359406, 9.487468, 9.615577, 9.743732, 9.871933, 10.00018, 
    10.12847, 10.2568, 10.38518, 10.5136, 10.64206, 10.77056, 10.89911, 
    11.02769, 11.15631, 11.28497, 11.41366, 11.5424, 11.67117, 11.79997, 
    11.92881, 12.05768, 12.18659, 12.31553, 12.4445, 12.5735, 12.70254, 
    12.8316, 12.96069, 13.08981, 13.21896, 13.34813, 13.47733, 13.60656, 
    13.73581, 13.86509, 13.99439, 14.12371, 14.25305, 14.38241, 14.5118, 
    14.6412, 14.77063, 14.90007, 15.02953, 15.15901, 15.2885, 15.418, 
    15.54753, 15.67706, 15.80661, 15.93617, 16.06575, 16.19533, 16.32493, 
    16.45453, 16.58414, 16.71376, 16.84339, 16.97303, 17.10267, 17.23232, 
    17.36197, 17.49162, 17.62127, 17.75093, 17.88059, 18.01026, 18.13992, 
    18.26958, 18.39923, 18.52889, 18.65854, 18.78819, 18.91784, 19.04748, 
    19.17711, 19.30674, 19.43636, 19.56597, 19.69557, 19.82517, 19.95475, 
    20.08432, 20.21388, 20.34343, 20.47296, 20.60248, 20.73199, 20.86148, 
    20.99095, 21.12041, 21.24985, 21.37927, 21.50867, 21.63805, 21.76741, 
    21.89675, 22.02607, 22.15536, 22.28464, 22.41388, 22.5431, 22.6723, 
    22.80147, 22.93062, 23.05973, 23.18882, 23.31788, 23.44691, 23.5759, 
    23.70487, 23.8338, 23.9627, 24.09157, 24.22041, 24.34921, 24.47797, 
    24.6067, 24.73539, 24.86404, 24.99265, 25.12123, 25.24977, 25.37826, 
    25.50672, 25.63513, 25.7635, 25.89183, 26.02011, 26.14835, 26.27654, 
    26.40469, 26.53279, 26.66085, 26.78885, 26.91681, 27.04472, 27.17258, 
    27.30039, 27.42815, 27.55585, 27.68351, 27.81111, 27.93865, 28.06614, 
    28.19358, 28.32096, 28.44829, 28.57556, 28.70277, 28.82992, 28.95701, 
    29.08405, 29.21102, 29.33793, 29.46479, 29.59158, 29.7183, 29.84497, 
    29.97157, 30.0981, 30.22458, 30.35098, 30.47732, 30.60359, 30.7298, 
    30.85593, 30.982, 31.108, 31.23393, 31.35979, 31.48558, 31.6113, 
    31.73694, 31.86251, 31.98801, 32.11344, 32.23879, 32.36407, 32.48927, 
    32.61439, 32.73944, 32.86441, 32.9893, 33.11412, 33.23886, 33.36351, 
    33.48809, 33.61259, 33.73701, 33.86134, 33.9856, 34.10977, 34.23386, 
    34.35786, 34.48178, 34.60562, 34.72937, 34.85303, 34.97662, 35.10011, 
    35.22352, 35.34684, 35.47007, 35.59321, 35.71627, 35.83923, 35.96211, 
    36.0849, 36.20759, 36.3302, 36.45271, 36.57513, 36.69746, 36.81969, 
    36.94183, 37.06388, 37.18584, 37.30769, 37.42946, 37.55113, 37.6727, 
    37.79418, 37.91556, 38.03684, 38.15802, 38.27911, 38.4001, 38.52099, 
    38.64178, 38.76247, 38.88306, 39.00355, 39.12394, 39.24423, 39.36442, 
    39.4845, 39.60448,
  -14.31282, -14.20334, -14.09373, -13.984, -13.87415, -13.76418, -13.65408, 
    -13.54387, -13.43353, -13.32306, -13.21248, -13.10177, -12.99094, 
    -12.87999, -12.76892, -12.65773, -12.54641, -12.43498, -12.32342, 
    -12.21174, -12.09994, -11.98802, -11.87598, -11.76382, -11.65154, 
    -11.53913, -11.42661, -11.31397, -11.20121, -11.08832, -10.97532, 
    -10.8622, -10.74896, -10.6356, -10.52212, -10.40852, -10.29481, 
    -10.18097, -10.06702, -9.95295, -9.838761, -9.724455, -9.610031, 
    -9.49549, -9.380832, -9.266057, -9.151165, -9.036157, -8.921032, 
    -8.805792, -8.690435, -8.574963, -8.459375, -8.343673, -8.227855, 
    -8.111922, -7.995875, -7.879714, -7.763439, -7.64705, -7.530548, 
    -7.413932, -7.297203, -7.180361, -7.063407, -6.946341, -6.829163, 
    -6.711873, -6.594472, -6.476959, -6.359336, -6.241602, -6.123758, 
    -6.005804, -5.88774, -5.769567, -5.651285, -5.532894, -5.414394, 
    -5.295786, -5.177071, -5.058248, -4.939317, -4.82028, -4.701137, 
    -4.581887, -4.462531, -4.34307, -4.223503, -4.103832, -3.984056, 
    -3.864176, -3.744192, -3.624104, -3.503914, -3.383621, -3.263226, 
    -3.142729, -3.02213, -2.901429, -2.780629, -2.659727, -2.538726, 
    -2.417625, -2.296424, -2.175125, -2.053728, -1.932232, -1.810639, 
    -1.688948, -1.567161, -1.445277, -1.323298, -1.201223, -1.079053, 
    -0.9567876, -0.8344285, -0.7119757, -0.5894295, -0.4667904, -0.3440588, 
    -0.2212353, -0.09832029, 0.02468582, 0.1477825, 0.2709694, 0.3942459, 
    0.5176116, 0.641066, 0.7646086, 0.888239, 1.011957, 1.135761, 1.259652, 
    1.383628, 1.50769, 1.631837, 1.756068, 1.880382, 2.00478, 2.129261, 
    2.253823, 2.378468, 2.503193, 2.628, 2.752886, 2.877852, 3.002897, 
    3.128021, 3.253222, 3.378501, 3.503857, 3.629289, 3.754797, 3.88038, 
    4.006038, 4.13177, 4.257575, 4.383453, 4.509403, 4.635426, 4.761519, 
    4.887683, 5.013918, 5.140222, 5.266594, 5.393035, 5.519544, 5.646119, 
    5.772761, 5.899469, 6.026242, 6.15308, 6.279983, 6.406948, 6.533976, 
    6.661067, 6.788218, 6.915431, 7.042705, 7.170038, 7.29743, 7.424881, 
    7.552389, 7.679955, 7.807577, 7.935255, 8.062988, 8.190776, 8.318618, 
    8.446512, 8.57446, 8.70246, 8.830511, 8.958612, 9.086764, 9.214965, 
    9.343215, 9.471513, 9.599857, 9.728249, 9.856687, 9.985169, 10.1137, 
    10.24227, 10.37088, 10.49954, 10.62824, 10.75698, 10.88576, 11.01458, 
    11.14344, 11.27234, 11.40127, 11.53025, 11.65926, 11.7883, 11.91738, 
    12.0465, 12.17564, 12.30482, 12.43404, 12.56328, 12.69255, 12.82186, 
    12.95119, 13.08055, 13.20994, 13.33936, 13.4688, 13.59827, 13.72777, 
    13.85729, 13.98683, 14.11639, 14.24598, 14.37559, 14.50521, 14.63486, 
    14.76453, 14.89421, 15.02392, 15.15364, 15.28337, 15.41313, 15.54289, 
    15.67267, 15.80247, 15.93227, 16.06209, 16.19192, 16.32176, 16.45161, 
    16.58147, 16.71133, 16.84121, 16.97109, 17.10097, 17.23086, 17.36076, 
    17.49066, 17.62056, 17.75046, 17.88037, 18.01027, 18.14018, 18.27009, 
    18.39999, 18.52989, 18.65979, 18.78968, 18.91957, 19.04946, 19.17934, 
    19.30921, 19.43908, 19.56893, 19.69878, 19.82862, 19.95844, 20.08826, 
    20.21807, 20.34786, 20.47763, 20.6074, 20.73715, 20.86688, 20.9966, 
    21.1263, 21.25598, 21.38565, 21.51529, 21.64492, 21.77452, 21.90411, 
    22.03367, 22.1632, 22.29272, 22.42221, 22.55167, 22.68111, 22.81053, 
    22.93991, 23.06927, 23.1986, 23.3279, 23.45717, 23.58641, 23.71561, 
    23.84479, 23.97393, 24.10304, 24.23211, 24.36115, 24.49016, 24.61912, 
    24.74805, 24.87695, 25.0058, 25.13461, 25.26339, 25.39212, 25.52081, 
    25.64947, 25.77807, 25.90664, 26.03516, 26.16363, 26.29206, 26.42045, 
    26.54879, 26.67708, 26.80532, 26.93351, 27.06166, 27.18975, 27.31779, 
    27.44578, 27.57372, 27.70161, 27.82944, 27.95722, 28.08495, 28.21261, 
    28.34023, 28.46778, 28.59528, 28.72272, 28.85011, 28.97743, 29.1047, 
    29.2319, 29.35904, 29.48612, 29.61314, 29.7401, 29.86699, 29.99382, 
    30.12058, 30.24728, 30.37391, 30.50047, 30.62697, 30.7534, 30.87976, 
    31.00606, 31.13228, 31.25843, 31.38451, 31.51052, 31.63646, 31.76233, 
    31.88812, 32.01384, 32.13949, 32.26506, 32.39056, 32.51598, 32.64132, 
    32.76659, 32.89178, 33.01689, 33.14192, 33.26687, 33.39175, 33.51654, 
    33.64125, 33.76588, 33.89043, 34.0149, 34.13929, 34.26359, 34.38781, 
    34.51194, 34.63599, 34.75995, 34.88383, 35.00762, 35.13132, 35.25494, 
    35.37847, 35.50191, 35.62526, 35.74852, 35.8717, 35.99478, 36.11777, 
    36.24067, 36.36348, 36.48619, 36.60882, 36.73135, 36.85379, 36.97614, 
    37.09838, 37.22054, 37.3426, 37.46457, 37.58643, 37.70821, 37.82988, 
    37.95146, 38.07294, 38.19432, 38.3156, 38.43679, 38.55787, 38.67886, 
    38.79974, 38.92053, 39.04121, 39.1618, 39.28228, 39.40266, 39.52293, 
    39.64311,
  -14.36686, -14.25724, -14.14749, -14.03762, -13.92763, -13.81752, 
    -13.70728, -13.59692, -13.48643, -13.37583, -13.2651, -13.15425, 
    -13.04327, -12.93218, -12.82096, -12.70962, -12.59815, -12.48657, 
    -12.37486, -12.26303, -12.15108, -12.03901, -11.92682, -11.81451, 
    -11.70207, -11.58952, -11.47684, -11.36405, -11.25113, -11.13809, 
    -11.02493, -10.91166, -10.79826, -10.68474, -10.57111, -10.45735, 
    -10.34348, -10.22948, -10.11537, -10.00114, -9.886788, -9.772321, 
    -9.657735, -9.543031, -9.428209, -9.31327, -9.198214, -9.08304, -8.96775, 
    -8.852344, -8.73682, -8.621181, -8.505424, -8.389554, -8.273567, 
    -8.157465, -8.041247, -7.924916, -7.808469, -7.691908, -7.575233, 
    -7.458445, -7.341542, -7.224526, -7.107398, -6.990156, -6.872802, 
    -6.755336, -6.637758, -6.520068, -6.402267, -6.284354, -6.16633, 
    -6.048197, -5.929953, -5.811599, -5.693135, -5.574562, -5.45588, 
    -5.337089, -5.21819, -5.099183, -4.980068, -4.860845, -4.741516, 
    -4.622079, -4.502537, -4.382888, -4.263133, -4.143273, -4.023308, 
    -3.903239, -3.783065, -3.662787, -3.542405, -3.42192, -3.301332, 
    -3.180642, -3.05985, -2.938956, -2.817961, -2.696864, -2.575667, 
    -2.45437, -2.332973, -2.211477, -2.089881, -1.968188, -1.846396, 
    -1.724506, -1.602519, -1.480435, -1.358255, -1.235978, -1.113606, 
    -0.9911391, -0.8685772, -0.745921, -0.6231709, -0.5003275, -0.3773911, 
    -0.2543622, -0.1312413, -0.008028875, 0.1152747, 0.2386689, 0.3621532, 
    0.4857272, 0.6093904, 0.7331424, 0.8569825, 0.9809104, 1.104926, 
    1.229028, 1.353216, 1.47749, 1.601849, 1.726293, 1.850821, 1.975433, 
    2.100128, 2.224905, 2.349765, 2.474707, 2.59973, 2.724833, 2.850016, 
    2.975279, 3.10062, 3.22604, 3.351538, 3.477113, 3.602765, 3.728493, 
    3.854297, 3.980176, 4.106129, 4.232156, 4.358257, 4.48443, 4.610676, 
    4.736993, 4.863381, 4.98984, 5.116368, 5.242966, 5.369632, 5.496367, 
    5.623169, 5.750038, 5.876973, 6.003973, 6.131039, 6.258169, 6.385363, 
    6.51262, 6.63994, 6.767322, 6.894765, 7.022269, 7.149832, 7.277456, 
    7.405138, 7.532877, 7.660675, 7.78853, 7.91644, 8.044407, 8.172428, 
    8.300503, 8.428632, 8.556814, 8.685048, 8.813334, 8.941671, 9.070058, 
    9.198495, 9.326981, 9.455514, 9.584096, 9.712725, 9.841399, 9.970119, 
    10.09888, 10.22769, 10.35655, 10.48544, 10.61438, 10.74336, 10.87238, 
    11.00144, 11.13054, 11.25968, 11.38885, 11.51807, 11.64732, 11.7766, 
    11.90592, 12.03528, 12.16467, 12.29409, 12.42354, 12.55303, 12.68254, 
    12.81209, 12.94167, 13.07127, 13.2009, 13.33056, 13.46025, 13.58996, 
    13.7197, 13.84946, 13.97925, 14.10905, 14.23888, 14.36874, 14.49861, 
    14.6285, 14.75841, 14.88834, 15.01829, 15.14826, 15.27824, 15.40823, 
    15.53825, 15.66827, 15.79831, 15.92836, 16.05843, 16.1885, 16.31859, 
    16.44868, 16.57878, 16.70889, 16.83901, 16.96914, 17.09927, 17.22941, 
    17.35955, 17.48969, 17.61984, 17.74999, 17.88014, 18.01029, 18.14045, 
    18.2706, 18.40075, 18.53089, 18.66104, 18.79118, 18.92131, 19.05145, 
    19.18157, 19.31169, 19.4418, 19.5719, 19.70199, 19.83208, 19.96215, 
    20.09221, 20.22226, 20.3523, 20.48232, 20.61233, 20.74232, 20.8723, 
    21.00227, 21.13221, 21.26214, 21.39205, 21.52194, 21.6518, 21.78165, 
    21.91148, 22.04128, 22.17107, 22.30083, 22.43056, 22.56027, 22.68995, 
    22.8196, 22.94923, 23.07883, 23.2084, 23.33795, 23.46746, 23.59694, 
    23.72639, 23.8558, 23.98519, 24.11454, 24.24385, 24.37313, 24.50238, 
    24.63158, 24.76075, 24.88988, 25.01898, 25.14803, 25.27705, 25.40602, 
    25.53495, 25.66384, 25.79268, 25.92149, 26.05025, 26.17896, 26.30763, 
    26.43625, 26.56482, 26.69335, 26.82183, 26.95025, 27.07863, 27.20696, 
    27.33524, 27.46347, 27.59164, 27.71976, 27.84783, 27.97584, 28.1038, 
    28.2317, 28.35954, 28.48733, 28.61506, 28.74274, 28.87035, 28.9979, 
    29.1254, 29.25283, 29.3802, 29.50751, 29.63476, 29.76195, 29.88906, 
    30.01612, 30.14311, 30.27003, 30.39689, 30.52369, 30.65041, 30.77707, 
    30.90365, 31.03017, 31.15662, 31.28299, 31.4093, 31.53553, 31.6617, 
    31.78778, 31.9138, 32.03974, 32.16561, 32.2914, 32.41711, 32.54276, 
    32.66832, 32.7938, 32.91921, 33.04454, 33.16979, 33.29496, 33.42005, 
    33.54506, 33.66999, 33.79484, 33.9196, 34.04428, 34.16888, 34.2934, 
    34.41783, 34.54218, 34.66644, 34.79061, 34.9147, 35.0387, 35.16261, 
    35.28644, 35.41018, 35.53382, 35.65739, 35.78086, 35.90424, 36.02753, 
    36.15072, 36.27383, 36.39684, 36.51976, 36.64259, 36.76533, 36.88797, 
    37.01052, 37.13297, 37.25533, 37.37759, 37.49975, 37.62182, 37.74379, 
    37.86567, 37.98745, 38.10912, 38.2307, 38.35218, 38.47356, 38.59484, 
    38.71603, 38.83711, 38.95809, 39.07896, 39.19974, 39.32042, 39.44099, 
    39.56145, 39.68182,
  -14.421, -14.31124, -14.20136, -14.09135, -13.98121, -13.87096, -13.76058, 
    -13.65007, -13.53945, -13.42869, -13.31782, -13.20683, -13.09571, 
    -12.98446, -12.8731, -12.76161, -12.65, -12.53827, -12.42641, -12.31443, 
    -12.20233, -12.09011, -11.97777, -11.8653, -11.75272, -11.64001, 
    -11.52718, -11.41423, -11.30116, -11.18797, -11.07465, -10.96122, 
    -10.84766, -10.73399, -10.6202, -10.50628, -10.39225, -10.27809, 
    -10.16382, -10.04943, -9.934918, -9.820289, -9.70554, -9.590672, 
    -9.475688, -9.360584, -9.245363, -9.130025, -9.014569, -8.898995, 
    -8.783305, -8.667499, -8.551575, -8.435534, -8.319379, -8.203107, 
    -8.08672, -7.970216, -7.853598, -7.736866, -7.620018, -7.503056, 
    -7.38598, -7.26879, -7.151486, -7.034069, -6.916539, -6.798896, 
    -6.681141, -6.563273, -6.445293, -6.327202, -6.209, -6.090686, -5.972261, 
    -5.853726, -5.735081, -5.616325, -5.49746, -5.378487, -5.259403, 
    -5.140212, -5.020912, -4.901504, -4.781988, -4.662365, -4.542635, 
    -4.422799, -4.302856, -4.182807, -4.062653, -3.942393, -3.822029, 
    -3.70156, -3.580986, -3.46031, -3.339529, -3.218646, -3.09766, -2.976571, 
    -2.855381, -2.734089, -2.612697, -2.491203, -2.369609, -2.247916, 
    -2.126122, -2.00423, -1.882239, -1.76015, -1.637962, -1.515678, 
    -1.393296, -1.270818, -1.148244, -1.025574, -0.9028092, -0.7799492, 
    -0.656995, -0.5339468, -0.4108052, -0.2875706, -0.1642435, -0.04082427, 
    0.08268652, 0.2062884, 0.329981, 0.4537638, 0.5776362, 0.7015978, 
    0.8256481, 0.9497867, 1.074013, 1.198327, 1.322727, 1.447213, 1.571786, 
    1.696443, 1.821185, 1.946012, 2.070922, 2.195915, 2.32099, 2.446148, 
    2.571388, 2.696708, 2.822109, 2.94759, 3.07315, 3.198789, 3.324506, 
    3.450301, 3.576174, 3.702122, 3.828147, 3.954247, 4.080423, 4.206673, 
    4.332996, 4.459393, 4.585862, 4.712403, 4.839015, 4.965699, 5.092453, 
    5.219276, 5.346169, 5.47313, 5.600159, 5.727254, 5.854417, 5.981646, 
    6.10894, 6.236299, 6.363722, 6.491209, 6.618759, 6.74637, 6.874044, 
    7.001779, 7.129574, 7.257428, 7.385342, 7.513315, 7.641345, 7.769432, 
    7.897576, 8.025776, 8.154031, 8.282341, 8.410705, 8.539121, 8.66759, 
    8.796112, 8.924685, 9.053308, 9.18198, 9.310702, 9.439473, 9.568293, 
    9.697158, 9.826071, 9.955029, 10.08403, 10.21308, 10.34217, 10.47131, 
    10.60048, 10.7297, 10.85896, 10.98826, 11.1176, 11.24698, 11.3764, 
    11.50585, 11.63534, 11.76487, 11.89443, 12.02403, 12.15366, 12.28332, 
    12.41302, 12.54275, 12.67251, 12.8023, 12.93211, 13.06196, 13.19184, 
    13.32174, 13.45167, 13.58163, 13.71161, 13.84162, 13.97165, 14.1017, 
    14.23177, 14.36187, 14.49199, 14.62212, 14.75228, 14.88246, 15.01265, 
    15.14286, 15.27309, 15.40333, 15.53359, 15.66386, 15.79414, 15.92444, 
    16.05475, 16.18507, 16.3154, 16.44574, 16.57609, 16.70645, 16.83681, 
    16.96719, 17.09756, 17.22795, 17.35834, 17.48873, 17.61912, 17.74952, 
    17.87992, 18.01031, 18.14071, 18.27111, 18.40151, 18.5319, 18.66229, 
    18.79268, 18.92306, 19.05344, 19.18381, 19.31417, 19.44453, 19.57488, 
    19.70522, 19.83554, 19.96586, 20.09617, 20.22647, 20.35675, 20.48702, 
    20.61727, 20.74751, 20.87774, 21.00795, 21.13814, 21.26831, 21.39846, 
    21.5286, 21.65871, 21.7888, 21.91887, 22.04892, 22.17895, 22.30895, 
    22.43893, 22.56888, 22.69881, 22.82871, 22.95858, 23.08842, 23.21824, 
    23.34802, 23.47778, 23.6075, 23.73719, 23.86685, 23.99648, 24.12607, 
    24.25562, 24.38514, 24.51463, 24.64408, 24.77349, 24.90286, 25.03219, 
    25.16149, 25.29074, 25.41995, 25.54912, 25.67825, 25.80734, 25.93638, 
    26.06537, 26.19432, 26.32323, 26.45209, 26.5809, 26.70966, 26.83838, 
    26.96704, 27.09566, 27.22422, 27.35274, 27.4812, 27.6096, 27.73796, 
    27.86626, 27.99451, 28.1227, 28.25083, 28.37891, 28.50693, 28.6349, 
    28.7628, 28.89065, 29.01843, 29.14616, 29.27382, 29.40142, 29.52896, 
    29.65644, 29.78385, 29.9112, 30.03848, 30.1657, 30.29285, 30.41994, 
    30.54696, 30.67391, 30.80079, 30.9276, 31.05434, 31.18102, 31.30762, 
    31.43415, 31.56061, 31.68699, 31.8133, 31.93954, 32.0657, 32.19179, 
    32.31781, 32.44374, 32.5696, 32.69538, 32.82109, 32.94672, 33.07227, 
    33.19773, 33.32312, 33.44843, 33.57365, 33.6988, 33.82386, 33.94884, 
    34.07374, 34.19855, 34.32328, 34.44793, 34.57248, 34.69696, 34.82134, 
    34.94564, 35.06985, 35.19398, 35.31802, 35.44196, 35.56582, 35.68959, 
    35.81327, 35.93686, 36.06035, 36.18376, 36.30707, 36.43029, 36.55342, 
    36.67645, 36.79939, 36.92223, 37.04499, 37.16764, 37.2902, 37.41266, 
    37.53503, 37.6573, 37.77947, 37.90154, 38.02352, 38.14539, 38.26717, 
    38.38885, 38.51043, 38.6319, 38.75328, 38.87456, 38.99573, 39.11681, 
    39.23777, 39.35864, 39.4794, 39.60007, 39.72062,
  -14.47525, -14.36535, -14.25533, -14.14517, -14.0349, -13.9245, -13.81398, 
    -13.70333, -13.59256, -13.48167, -13.37065, -13.25951, -13.14824, 
    -13.03685, -12.92534, -12.81371, -12.70195, -12.59007, -12.47806, 
    -12.36594, -12.25369, -12.14131, -12.02882, -11.9162, -11.80346, 
    -11.6906, -11.57762, -11.46451, -11.35129, -11.23794, -11.12447, 
    -11.01088, -10.89717, -10.78334, -10.66939, -10.55532, -10.44112, 
    -10.32681, -10.21238, -10.09782, -9.98315, -9.868359, -9.753448, 
    -9.638417, -9.523269, -9.408001, -9.292615, -9.177111, -9.061489, 
    -8.945749, -8.829892, -8.713917, -8.597825, -8.481616, -8.365291, 
    -8.248849, -8.132291, -8.015617, -7.898828, -7.781922, -7.664902, 
    -7.547766, -7.430516, -7.313152, -7.195673, -7.078081, -6.960374, 
    -6.842555, -6.724622, -6.606576, -6.488418, -6.370148, -6.251765, 
    -6.133271, -6.014666, -5.895949, -5.777122, -5.658185, -5.539137, 
    -5.419979, -5.300712, -5.181336, -5.061851, -4.942257, -4.822555, 
    -4.702745, -4.582828, -4.462803, -4.342672, -4.222434, -4.10209, 
    -3.98164, -3.861085, -3.740424, -3.619659, -3.49879, -3.377817, -3.25674, 
    -3.13556, -3.014277, -2.892891, -2.771404, -2.649815, -2.528125, 
    -2.406333, -2.284442, -2.16245, -2.040359, -1.918169, -1.79588, 
    -1.673492, -1.551007, -1.428424, -1.305743, -1.182967, -1.060094, 
    -0.9371251, -0.8140611, -0.6909022, -0.5676489, -0.4443017, -0.320861, 
    -0.1973272, -0.07370089, 0.05001754, 0.1738276, 0.2977288, 0.4217207, 
    0.5458027, 0.6699744, 0.7942354, 0.9185851, 1.043023, 1.167549, 1.292161, 
    1.416861, 1.541647, 1.666518, 1.791475, 1.916516, 2.041641, 2.16685, 
    2.292142, 2.417517, 2.542974, 2.668512, 2.794131, 2.91983, 3.045609, 
    3.171468, 3.297405, 3.42342, 3.549513, 3.675683, 3.80193, 3.928252, 
    4.05465, 4.181123, 4.30767, 4.43429, 4.560983, 4.687749, 4.814587, 
    4.941496, 5.068475, 5.195525, 5.322644, 5.449832, 5.577088, 5.704412, 
    5.831803, 5.95926, 6.086783, 6.214371, 6.342024, 6.469741, 6.597521, 
    6.725364, 6.853268, 6.981235, 7.109261, 7.237348, 7.365495, 7.4937, 
    7.621963, 7.750284, 7.878662, 8.007096, 8.135586, 8.26413, 8.392729, 
    8.52138, 8.650085, 8.778843, 8.907652, 9.036512, 9.165422, 9.294381, 
    9.423389, 9.552446, 9.68155, 9.810701, 9.939898, 10.06914, 10.19843, 
    10.32776, 10.45713, 10.58655, 10.71601, 10.84551, 10.97505, 11.10463, 
    11.23425, 11.36391, 11.4936, 11.62334, 11.75311, 11.88291, 12.01275, 
    12.14262, 12.27253, 12.40247, 12.53244, 12.66244, 12.79247, 12.92254, 
    13.05263, 13.18275, 13.3129, 13.44307, 13.57327, 13.7035, 13.83375, 
    13.96402, 14.09432, 14.22464, 14.35498, 14.48535, 14.61573, 14.74613, 
    14.87655, 15.00699, 15.13745, 15.26792, 15.39841, 15.52892, 15.65943, 
    15.78996, 15.92051, 16.05106, 16.18163, 16.31221, 16.4428, 16.57339, 
    16.704, 16.83461, 16.96523, 17.09585, 17.22648, 17.35712, 17.48776, 
    17.6184, 17.74904, 17.87969, 18.01033, 18.14098, 18.27162, 18.40227, 
    18.53291, 18.66355, 18.79418, 18.92481, 19.05543, 19.18605, 19.31666, 
    19.44727, 19.57786, 19.70845, 19.83902, 19.96959, 20.10014, 20.23068, 
    20.36121, 20.49173, 20.62223, 20.75272, 20.88319, 21.01364, 21.14408, 
    21.2745, 21.4049, 21.53527, 21.66563, 21.79597, 21.92629, 22.05659, 
    22.18686, 22.3171, 22.44732, 22.57752, 22.70769, 22.83784, 22.96795, 
    23.09804, 23.2281, 23.35812, 23.48812, 23.61809, 23.74802, 23.87792, 
    24.00779, 24.13763, 24.26743, 24.39719, 24.52691, 24.6566, 24.78626, 
    24.91587, 25.04544, 25.17498, 25.30447, 25.43393, 25.56334, 25.6927, 
    25.82203, 25.95131, 26.08054, 26.20973, 26.33887, 26.46797, 26.59702, 
    26.72602, 26.85497, 26.98388, 27.11273, 27.24153, 27.37028, 27.49897, 
    27.62762, 27.75621, 27.88474, 28.01322, 28.14165, 28.27002, 28.39833, 
    28.52658, 28.65478, 28.78292, 28.911, 29.03901, 29.16697, 29.29486, 
    29.4227, 29.55047, 29.67817, 29.80581, 29.93339, 30.06091, 30.18835, 
    30.31573, 30.44305, 30.57029, 30.69747, 30.82458, 30.95162, 31.07858, 
    31.20548, 31.33231, 31.45906, 31.58574, 31.71235, 31.83889, 31.96535, 
    32.09174, 32.21804, 32.34428, 32.47044, 32.59652, 32.72252, 32.84845, 
    32.97429, 33.10006, 33.22575, 33.35135, 33.47688, 33.60232, 33.72768, 
    33.85296, 33.97816, 34.10327, 34.2283, 34.35324, 34.4781, 34.60287, 
    34.72755, 34.85215, 34.97667, 35.10109, 35.22543, 35.34967, 35.47383, 
    35.5979, 35.72188, 35.84576, 35.96956, 36.09326, 36.21687, 36.34039, 
    36.46382, 36.58715, 36.71039, 36.83353, 36.95658, 37.07954, 37.2024, 
    37.32516, 37.44782, 37.57039, 37.69286, 37.81523, 37.9375, 38.05968, 
    38.18176, 38.30373, 38.42561, 38.54738, 38.66906, 38.79063, 38.9121, 
    39.03347, 39.15474, 39.2759, 39.39696, 39.51792, 39.63877, 39.75952,
  -14.52961, -14.41957, -14.3094, -14.19911, -14.08869, -13.97815, -13.86749, 
    -13.7567, -13.64578, -13.53475, -13.42358, -13.3123, -13.20089, 
    -13.08935, -12.97769, -12.86591, -12.754, -12.64197, -12.52982, 
    -12.41754, -12.30514, -12.19262, -12.07997, -11.96721, -11.85431, 
    -11.7413, -11.62816, -11.5149, -11.40152, -11.28802, -11.1744, -11.06065, 
    -10.94678, -10.83279, -10.71868, -10.60445, -10.4901, -10.37563, 
    -10.26103, -10.14632, -10.03149, -9.916532, -9.801457, -9.686264, 
    -9.570951, -9.45552, -9.339969, -9.224299, -9.108511, -8.992604, 
    -8.87658, -8.760437, -8.644177, -8.5278, -8.411304, -8.294692, -8.177963, 
    -8.061118, -7.944157, -7.827079, -7.709886, -7.592577, -7.475152, 
    -7.357614, -7.239959, -7.122191, -7.004308, -6.886312, -6.768201, 
    -6.649978, -6.531641, -6.413191, -6.294629, -6.175954, -6.057168, 
    -5.93827, -5.819261, -5.70014, -5.58091, -5.461568, -5.342116, -5.222555, 
    -5.102885, -4.983105, -4.863216, -4.743219, -4.623114, -4.502901, 
    -4.382581, -4.262154, -4.14162, -4.020979, -3.900233, -3.779381, 
    -3.658424, -3.537362, -3.416195, -3.294924, -3.17355, -3.052072, 
    -2.930491, -2.808808, -2.687023, -2.565135, -2.443146, -2.321057, 
    -2.198867, -2.076576, -1.954186, -1.831697, -1.709108, -1.586421, 
    -1.463637, -1.340754, -1.217774, -1.094698, -0.9715255, -0.848257, 
    -0.7248932, -0.6014344, -0.4778811, -0.3542339, -0.2304931, -0.1066592, 
    0.01726721, 0.1412858, 0.265396, 0.3895974, 0.5138896, 0.6382718, 
    0.7627438, 0.887305, 1.011955, 1.136693, 1.261519, 1.386432, 1.511431, 
    1.636517, 1.761689, 1.886945, 2.012287, 2.137712, 2.263221, 2.388813, 
    2.514487, 2.640243, 2.766081, 2.891999, 3.017998, 3.144076, 3.270234, 
    3.39647, 3.522784, 3.649176, 3.775645, 3.90219, 4.028811, 4.155507, 
    4.282277, 4.409122, 4.53604, 4.663031, 4.790094, 4.917229, 5.044435, 
    5.171711, 5.299057, 5.426473, 5.553957, 5.681509, 5.809129, 5.936815, 
    6.064568, 6.192386, 6.320269, 6.448216, 6.576227, 6.704301, 6.832438, 
    6.960636, 7.088895, 7.217215, 7.345594, 7.474032, 7.60253, 7.731085, 
    7.859697, 7.988366, 8.11709, 8.245871, 8.374704, 8.503592, 8.632534, 
    8.761528, 8.890574, 9.019671, 9.148819, 9.278016, 9.407263, 9.536558, 
    9.6659, 9.79529, 9.924726, 10.05421, 10.18373, 10.31331, 10.44292, 
    10.57258, 10.70228, 10.83202, 10.9618, 11.09162, 11.22148, 11.35138, 
    11.48132, 11.6113, 11.74131, 11.87136, 12.00144, 12.13155, 12.26171, 
    12.39189, 12.5221, 12.65235, 12.78263, 12.91293, 13.04327, 13.17364, 
    13.30403, 13.43445, 13.56489, 13.69537, 13.82586, 13.95638, 14.08693, 
    14.21749, 14.34808, 14.47869, 14.60932, 14.73997, 14.87064, 15.00132, 
    15.13202, 15.26274, 15.39348, 15.52423, 15.65499, 15.78577, 15.91656, 
    16.04737, 16.17818, 16.30901, 16.43984, 16.57069, 16.70154, 16.8324, 
    16.96327, 17.09414, 17.22502, 17.3559, 17.48679, 17.61768, 17.74857, 
    17.87946, 18.01035, 18.14125, 18.27214, 18.40303, 18.53392, 18.6648, 
    18.79569, 18.92656, 19.05743, 19.1883, 19.31916, 19.45001, 19.58085, 
    19.71169, 19.84251, 19.97332, 20.10413, 20.23491, 20.36569, 20.49645, 
    20.6272, 20.75793, 20.88865, 21.01935, 21.15004, 21.2807, 21.41135, 
    21.54197, 21.67258, 21.80316, 21.93373, 22.06427, 22.19478, 22.32528, 
    22.45574, 22.58618, 22.7166, 22.84699, 22.97735, 23.10768, 23.23798, 
    23.36826, 23.4985, 23.62871, 23.75888, 23.88903, 24.01914, 24.14922, 
    24.27926, 24.40927, 24.53923, 24.66917, 24.79906, 24.92892, 25.05873, 
    25.18851, 25.31824, 25.44794, 25.57759, 25.70719, 25.83676, 25.96628, 
    26.09575, 26.22518, 26.35456, 26.4839, 26.61319, 26.74242, 26.87161, 
    27.00075, 27.12984, 27.25888, 27.38787, 27.5168, 27.64568, 27.7745, 
    27.90328, 28.03199, 28.16065, 28.28926, 28.4178, 28.54629, 28.67472, 
    28.80309, 28.9314, 29.05965, 29.18784, 29.31596, 29.44403, 29.57203, 
    29.69996, 29.82784, 29.95564, 30.08339, 30.21106, 30.33867, 30.46621, 
    30.59369, 30.72109, 30.84843, 30.97569, 31.10289, 31.23001, 31.35706, 
    31.48404, 31.61095, 31.73778, 31.86454, 31.99122, 32.11783, 32.24437, 
    32.37082, 32.4972, 32.6235, 32.74973, 32.87587, 33.00194, 33.12793, 
    33.25383, 33.37965, 33.5054, 33.63106, 33.75664, 33.88213, 34.00755, 
    34.13287, 34.25812, 34.38327, 34.50835, 34.63334, 34.75823, 34.88305, 
    35.00777, 35.1324, 35.25695, 35.38141, 35.50578, 35.63005, 35.75424, 
    35.87834, 36.00234, 36.12626, 36.25007, 36.3738, 36.49743, 36.62097, 
    36.74442, 36.86776, 36.99102, 37.11417, 37.23724, 37.3602, 37.48307, 
    37.60583, 37.72851, 37.85108, 37.97355, 38.09593, 38.2182, 38.34038, 
    38.46245, 38.58442, 38.7063, 38.82806, 38.94973, 39.0713, 39.19276, 
    39.31411, 39.43537, 39.55652, 39.67756, 39.7985,
  -14.58407, -14.47389, -14.36358, -14.25315, -14.14259, -14.03191, -13.9211, 
    -13.81017, -13.69911, -13.58793, -13.47662, -13.36519, -13.25363, 
    -13.14195, -13.03015, -12.91822, -12.80616, -12.69398, -12.58168, 
    -12.46926, -12.35671, -12.24403, -12.13124, -12.01831, -11.90527, 
    -11.7921, -11.67881, -11.5654, -11.45187, -11.33821, -11.22443, 
    -11.11052, -10.9965, -10.88235, -10.76808, -10.65369, -10.53918, 
    -10.42455, -10.30979, -10.19492, -10.07992, -9.964808, -9.849571, 
    -9.734215, -9.618738, -9.503141, -9.387425, -9.27159, -9.155636, 
    -9.039562, -8.92337, -8.80706, -8.690631, -8.574084, -8.457419, 
    -8.340637, -8.223738, -8.106721, -7.989587, -7.872337, -7.754971, 
    -7.637488, -7.519889, -7.402175, -7.284346, -7.166401, -7.048342, 
    -6.930168, -6.81188, -6.693478, -6.574962, -6.456333, -6.337591, 
    -6.218736, -6.099768, -5.980688, -5.861496, -5.742193, -5.622779, 
    -5.503253, -5.383617, -5.263871, -5.144014, -5.024048, -4.903973, 
    -4.783788, -4.663496, -4.543094, -4.422585, -4.301968, -4.181243, 
    -4.060412, -3.939475, -3.818431, -3.697281, -3.576026, -3.454666, 
    -3.333201, -3.211632, -3.089959, -2.968182, -2.846303, -2.72432, 
    -2.602236, -2.480049, -2.357761, -2.235371, -2.112881, -1.990291, 
    -1.867601, -1.744812, -1.621923, -1.498936, -1.375851, -1.252668, 
    -1.129388, -1.006011, -0.8825375, -0.7589683, -0.6353037, -0.511544, 
    -0.3876899, -0.2637417, -0.1396999, -0.01556499, 0.1086625, 0.2329822, 
    0.3573936, 0.4818961, 0.6064894, 0.7311728, 0.8559459, 0.9808083, 
    1.105759, 1.230798, 1.355925, 1.481139, 1.60644, 1.731827, 1.857299, 
    1.982857, 2.108499, 2.234225, 2.360034, 2.485927, 2.611902, 2.737958, 
    2.864096, 2.990315, 3.116614, 3.242992, 3.36945, 3.495986, 3.6226, 
    3.749291, 3.87606, 4.002904, 4.129824, 4.256819, 4.383888, 4.511032, 
    4.638248, 4.765537, 4.892899, 5.020331, 5.147835, 5.275409, 5.403053, 
    5.530765, 5.658546, 5.786395, 5.914311, 6.042294, 6.170342, 6.298456, 
    6.426634, 6.554877, 6.683183, 6.811551, 6.939982, 7.068474, 7.197027, 
    7.32564, 7.454313, 7.583045, 7.711834, 7.840682, 7.969585, 8.098546, 
    8.227562, 8.356632, 8.485757, 8.614936, 8.744167, 8.87345, 9.002786, 
    9.132171, 9.261607, 9.391092, 9.520626, 9.650208, 9.779838, 9.909513, 
    10.03924, 10.169, 10.29881, 10.42867, 10.55857, 10.68851, 10.81849, 
    10.94852, 11.07858, 11.20868, 11.33883, 11.46901, 11.59923, 11.72948, 
    11.85977, 11.9901, 12.12046, 12.25085, 12.38128, 12.51174, 12.64223, 
    12.77275, 12.90331, 13.03389, 13.1645, 13.29514, 13.4258, 13.55649, 
    13.68721, 13.81795, 13.94872, 14.07951, 14.21032, 14.34116, 14.47201, 
    14.60289, 14.73378, 14.8647, 14.99563, 15.12658, 15.25755, 15.38853, 
    15.51953, 15.65055, 15.78157, 15.91261, 16.04366, 16.17472, 16.3058, 
    16.43688, 16.56797, 16.69907, 16.83018, 16.9613, 17.09242, 17.22355, 
    17.35468, 17.48581, 17.61695, 17.74809, 17.87923, 18.01037, 18.14151, 
    18.27266, 18.4038, 18.53493, 18.66607, 18.7972, 18.92832, 19.05944, 
    19.19056, 19.32166, 19.45276, 19.58385, 19.71494, 19.84601, 19.97707, 
    20.10812, 20.23916, 20.37018, 20.50119, 20.63219, 20.76317, 20.89413, 
    21.02508, 21.15601, 21.28692, 21.41782, 21.54869, 21.67954, 21.81037, 
    21.94118, 22.07197, 22.20273, 22.33347, 22.46418, 22.59487, 22.72553, 
    22.85616, 22.98677, 23.11735, 23.2479, 23.37841, 23.5089, 23.63935, 
    23.76978, 23.90017, 24.03052, 24.16084, 24.29113, 24.42138, 24.55159, 
    24.68176, 24.8119, 24.942, 25.07205, 25.20207, 25.33205, 25.46198, 
    25.59188, 25.72172, 25.85153, 25.98129, 26.111, 26.24067, 26.37029, 
    26.49987, 26.62939, 26.75887, 26.8883, 27.01768, 27.147, 27.27628, 
    27.4055, 27.53467, 27.66379, 27.79285, 27.92186, 28.05081, 28.1797, 
    28.30854, 28.43732, 28.56605, 28.69471, 28.82331, 28.95185, 29.08034, 
    29.20876, 29.33712, 29.46541, 29.59365, 29.72181, 29.84992, 29.97795, 
    30.10593, 30.23383, 30.36167, 30.48944, 30.61714, 30.74478, 30.87234, 
    30.99983, 31.12725, 31.2546, 31.38188, 31.50908, 31.63622, 31.76328, 
    31.89026, 32.01717, 32.144, 32.27076, 32.39743, 32.52404, 32.65056, 
    32.777, 32.90337, 33.02966, 33.15586, 33.28199, 33.40803, 33.53399, 
    33.65987, 33.78567, 33.91138, 34.03701, 34.16256, 34.28801, 34.41339, 
    34.53867, 34.66387, 34.78899, 34.91401, 35.03895, 35.1638, 35.28856, 
    35.41323, 35.5378, 35.66229, 35.78669, 35.911, 36.03521, 36.15933, 
    36.28336, 36.40729, 36.53113, 36.65487, 36.77852, 36.90208, 37.02553, 
    37.1489, 37.27216, 37.39533, 37.5184, 37.64137, 37.76424, 37.88702, 
    38.00969, 38.13226, 38.25474, 38.37711, 38.49938, 38.62156, 38.74362, 
    38.86559, 38.98745, 39.10921, 39.23087, 39.35242, 39.47387, 39.59521, 
    39.71645, 39.83759,
  -14.63863, -14.52831, -14.41787, -14.30729, -14.1966, -14.08577, -13.97482, 
    -13.86375, -13.75255, -13.64122, -13.52977, -13.41819, -13.30649, 
    -13.19466, -13.08271, -12.97063, -12.85843, -12.7461, -12.63365, 
    -12.52108, -12.40837, -12.29555, -12.1826, -12.06953, -11.95633, 
    -11.84301, -11.72957, -11.616, -11.50231, -11.3885, -11.27456, -11.1605, 
    -11.04632, -10.93202, -10.81759, -10.70304, -10.58837, -10.47357, 
    -10.35866, -10.24362, -10.12847, -10.01319, -9.897789, -9.782269, 
    -9.666628, -9.550867, -9.434986, -9.318985, -9.202864, -9.086623, 
    -8.970263, -8.853786, -8.737187, -8.620472, -8.503637, -8.386684, 
    -8.269613, -8.152425, -8.035119, -7.917696, -7.800157, -7.6825, 
    -7.564727, -7.446837, -7.328832, -7.210711, -7.092475, -6.974124, 
    -6.855658, -6.737077, -6.618382, -6.499574, -6.380651, -6.261615, 
    -6.142467, -6.023205, -5.903831, -5.784344, -5.664746, -5.545036, 
    -5.425215, -5.305283, -5.185241, -5.065088, -4.944825, -4.824453, 
    -4.703972, -4.583382, -4.462683, -4.341876, -4.220961, -4.099939, 
    -3.97881, -3.857574, -3.736231, -3.614783, -3.493229, -3.371569, 
    -3.249805, -3.127937, -3.005964, -2.883888, -2.761708, -2.639426, 
    -2.517041, -2.394554, -2.271965, -2.149276, -2.026485, -1.903594, 
    -1.780603, -1.657512, -1.534323, -1.411034, -1.287648, -1.164163, 
    -1.040582, -0.9169032, -0.7931283, -0.6692573, -0.5452909, -0.4212295, 
    -0.2970735, -0.1728233, -0.04847958, 0.07595731, 0.2004869, 0.3251086, 
    0.449822, 0.5746266, 0.6995219, 0.8245074, 0.9495826, 1.074747, 1.2, 
    1.325341, 1.45077, 1.576286, 1.701889, 1.827577, 1.953352, 2.079211, 
    2.205155, 2.331182, 2.457293, 2.583487, 2.709764, 2.836122, 2.962561, 
    3.089081, 3.21568, 3.34236, 3.469118, 3.595955, 3.722869, 3.849861, 
    3.976929, 4.104074, 4.231294, 4.358588, 4.485958, 4.6134, 4.740916, 
    4.868505, 4.996164, 5.123896, 5.251698, 5.37957, 5.507512, 5.635522, 
    5.763601, 5.891747, 6.01996, 6.14824, 6.276585, 6.404995, 6.533469, 
    6.662008, 6.790609, 6.919273, 7.047999, 7.176785, 7.305633, 7.43454, 
    7.563507, 7.692532, 7.821614, 7.950755, 8.079951, 8.209204, 8.338511, 
    8.467874, 8.597289, 8.726759, 8.85628, 8.985853, 9.115478, 9.245152, 
    9.374878, 9.504651, 9.634473, 9.764342, 9.894259, 10.02422, 10.15423, 
    10.28428, 10.41438, 10.54452, 10.6747, 10.80493, 10.9352, 11.0655, 
    11.19585, 11.32623, 11.45666, 11.58712, 11.71762, 11.84816, 11.97873, 
    12.10933, 12.23997, 12.37064, 12.50135, 12.63208, 12.76285, 12.89365, 
    13.02448, 13.15533, 13.28622, 13.41713, 13.54807, 13.67903, 13.81002, 
    13.94103, 14.07207, 14.20313, 14.33421, 14.46532, 14.59644, 14.72758, 
    14.85875, 14.98993, 15.12113, 15.25234, 15.38357, 15.51482, 15.64608, 
    15.77736, 15.90865, 16.03995, 16.17126, 16.30258, 16.43391, 16.56525, 
    16.6966, 16.82796, 16.95932, 17.09069, 17.22207, 17.35345, 17.48483, 
    17.61622, 17.74761, 17.879, 18.01039, 18.14178, 18.27317, 18.40456, 
    18.53595, 18.66733, 18.79871, 18.93009, 19.06146, 19.19282, 19.32417, 
    19.45552, 19.58686, 19.71819, 19.84952, 19.98083, 20.11212, 20.24341, 
    20.37468, 20.50594, 20.63719, 20.76841, 20.89963, 21.03082, 21.162, 
    21.29316, 21.4243, 21.55542, 21.68652, 21.8176, 21.94866, 22.07969, 
    22.2107, 22.34169, 22.47265, 22.60358, 22.73449, 22.86537, 22.99622, 
    23.12704, 23.25784, 23.3886, 23.51933, 23.65003, 23.7807, 23.91133, 
    24.04193, 24.1725, 24.30303, 24.43352, 24.56397, 24.69439, 24.82477, 
    24.95511, 25.08541, 25.21567, 25.34589, 25.47607, 25.6062, 25.73629, 
    25.86634, 25.99634, 26.1263, 26.2562, 26.38607, 26.51588, 26.64565, 
    26.77536, 26.90503, 27.03465, 27.16421, 27.29373, 27.42319, 27.55259, 
    27.68195, 27.81124, 27.94049, 28.06968, 28.19881, 28.32788, 28.4569, 
    28.58586, 28.71475, 28.84359, 28.97237, 29.10108, 29.22974, 29.35833, 
    29.48686, 29.61532, 29.74372, 29.87206, 30.00033, 30.12853, 30.25666, 
    30.38473, 30.51273, 30.64066, 30.76852, 30.89631, 31.02403, 31.15168, 
    31.27926, 31.40676, 31.53419, 31.66155, 31.78884, 31.91604, 32.04317, 
    32.17023, 32.29721, 32.42411, 32.55094, 32.67768, 32.80435, 32.93094, 
    33.05745, 33.18387, 33.31022, 33.43648, 33.56266, 33.68876, 33.81477, 
    33.9407, 34.06655, 34.19231, 34.31799, 34.44357, 34.56908, 34.69449, 
    34.81982, 34.94506, 35.07021, 35.19527, 35.32024, 35.44512, 35.56991, 
    35.69461, 35.81922, 35.94373, 36.06815, 36.19249, 36.31672, 36.44086, 
    36.56491, 36.68886, 36.81271, 36.93647, 37.06014, 37.1837, 37.30717, 
    37.43054, 37.55381, 37.67699, 37.80006, 37.92304, 38.04591, 38.16869, 
    38.29136, 38.41394, 38.53641, 38.65878, 38.78104, 38.90321, 39.02526, 
    39.14722, 39.26907, 39.39082, 39.51246, 39.634, 39.75543, 39.87676,
  -14.69331, -14.58285, -14.47226, -14.36155, -14.25071, -14.13974, 
    -14.02865, -13.91743, -13.80609, -13.69462, -13.58302, -13.4713, 
    -13.35945, -13.24748, -13.13538, -13.02315, -12.9108, -12.79833, 
    -12.68573, -12.573, -12.46015, -12.34717, -12.23407, -12.12085, -12.0075, 
    -11.89403, -11.78043, -11.66671, -11.55286, -11.43889, -11.3248, 
    -11.21059, -11.09625, -10.98178, -10.8672, -10.75249, -10.63766, 
    -10.52271, -10.40763, -10.29243, -10.17711, -10.06167, -9.946112, 
    -9.830427, -9.714622, -9.598697, -9.48265, -9.366483, -9.250196, 
    -9.133788, -9.017261, -8.900614, -8.783848, -8.666962, -8.549957, 
    -8.432834, -8.315592, -8.198232, -8.080753, -7.963158, -7.845444, 
    -7.727613, -7.609666, -7.491601, -7.37342, -7.255123, -7.13671, 
    -7.018181, -6.899537, -6.780777, -6.661903, -6.542914, -6.423811, 
    -6.304594, -6.185264, -6.06582, -5.946262, -5.826593, -5.70681, 
    -5.586916, -5.46691, -5.346793, -5.226564, -5.106224, -4.985774, 
    -4.865214, -4.744544, -4.623765, -4.502876, -4.381879, -4.260774, 
    -4.13956, -4.018239, -3.89681, -3.775275, -3.653633, -3.531885, 
    -3.410031, -3.288071, -3.166007, -3.043838, -2.921565, -2.799187, 
    -2.676707, -2.554123, -2.431437, -2.308649, -2.185759, -2.062768, 
    -1.939675, -1.816482, -1.693189, -1.569797, -1.446305, -1.322714, 
    -1.199025, -1.075239, -0.9513546, -0.8273735, -0.7032959, -0.5791224, 
    -0.4548532, -0.330489, -0.2060301, -0.08147711, 0.04316954, 0.1679094, 
    0.2927419, 0.4176666, 0.5426829, 0.6677905, 0.7929888, 0.9182773, 
    1.043656, 1.169123, 1.294679, 1.420323, 1.546055, 1.671874, 1.797779, 
    1.92377, 2.049847, 2.176009, 2.302256, 2.428586, 2.554999, 2.681495, 
    2.808074, 2.934734, 3.061475, 3.188297, 3.315199, 3.44218, 3.56924, 
    3.696378, 3.823594, 3.950887, 4.078256, 4.205701, 4.333222, 4.460817, 
    4.588487, 4.716229, 4.844046, 4.971933, 5.099893, 5.227924, 5.356026, 
    5.484197, 5.612437, 5.740746, 5.869123, 5.997567, 6.126078, 6.254655, 
    6.383297, 6.512005, 6.640776, 6.769611, 6.898509, 7.027468, 7.15649, 
    7.285572, 7.414714, 7.543916, 7.673177, 7.802496, 7.931873, 8.061306, 
    8.190796, 8.320341, 8.449941, 8.579596, 8.709303, 8.839063, 8.968876, 
    9.09874, 9.228654, 9.358619, 9.488632, 9.618695, 9.748805, 9.878963, 
    10.00917, 10.13942, 10.26971, 10.40005, 10.53043, 10.66086, 10.79133, 
    10.92184, 11.05239, 11.18298, 11.31361, 11.44428, 11.57498, 11.70573, 
    11.83651, 11.96732, 12.09817, 12.22906, 12.35997, 12.49092, 12.62191, 
    12.75292, 12.88397, 13.01504, 13.14614, 13.27727, 13.40843, 13.53962, 
    13.67083, 13.80207, 13.93333, 14.06461, 14.19592, 14.32725, 14.4586, 
    14.58998, 14.72137, 14.85278, 14.98421, 15.11566, 15.24712, 15.3786, 
    15.5101, 15.64161, 15.77313, 15.90467, 16.03622, 16.16778, 16.29935, 
    16.43093, 16.56252, 16.69412, 16.82573, 16.95734, 17.08896, 17.22059, 
    17.35222, 17.48385, 17.61549, 17.74713, 17.87877, 18.01041, 18.14205, 
    18.27369, 18.40533, 18.53697, 18.6686, 18.80023, 18.93186, 19.06347, 
    19.19509, 19.32669, 19.45829, 19.58988, 19.72146, 19.85303, 19.98459, 
    20.11614, 20.24767, 20.3792, 20.5107, 20.6422, 20.77368, 20.90514, 
    21.03658, 21.16801, 21.29942, 21.43081, 21.56218, 21.69352, 21.82485, 
    21.95616, 22.08744, 22.21869, 22.34993, 22.48113, 22.61232, 22.74347, 
    22.8746, 23.0057, 23.13676, 23.26781, 23.39881, 23.52979, 23.66074, 
    23.79165, 23.92253, 24.05337, 24.18418, 24.31496, 24.4457, 24.5764, 
    24.70706, 24.83768, 24.96827, 25.09881, 25.22931, 25.35977, 25.49019, 
    25.62057, 25.7509, 25.88119, 26.01143, 26.14163, 26.27178, 26.40188, 
    26.53194, 26.66194, 26.7919, 26.92181, 27.05166, 27.18147, 27.31122, 
    27.44092, 27.57056, 27.70016, 27.82969, 27.95917, 28.0886, 28.21796, 
    28.34727, 28.47653, 28.60572, 28.73485, 28.86392, 28.99294, 29.12189, 
    29.25077, 29.3796, 29.50836, 29.63706, 29.76569, 29.89425, 30.02275, 
    30.15119, 30.27955, 30.40785, 30.53608, 30.66424, 30.79233, 30.92035, 
    31.0483, 31.17618, 31.30398, 31.43171, 31.55937, 31.68695, 31.81446, 
    31.9419, 32.06926, 32.19653, 32.32374, 32.45086, 32.57791, 32.70488, 
    32.83177, 32.95858, 33.08531, 33.21196, 33.33852, 33.465, 33.5914, 
    33.71772, 33.84395, 33.9701, 34.09616, 34.22214, 34.34803, 34.47384, 
    34.59956, 34.72519, 34.85073, 34.97618, 35.10155, 35.22682, 35.35201, 
    35.4771, 35.6021, 35.72701, 35.85183, 35.97655, 36.10118, 36.22572, 
    36.35017, 36.47452, 36.59877, 36.72293, 36.84699, 36.97096, 37.09483, 
    37.2186, 37.34227, 37.46585, 37.58932, 37.7127, 37.83598, 37.95915, 
    38.08223, 38.2052, 38.32808, 38.45085, 38.57352, 38.69609, 38.81855, 
    38.94091, 39.06317, 39.18532, 39.30737, 39.42931, 39.55115, 39.67288, 
    39.79451, 39.91603,
  -14.74809, -14.63749, -14.52676, -14.41591, -14.30493, -14.19382, 
    -14.08259, -13.97122, -13.85974, -13.74812, -13.63638, -13.52451, 
    -13.41252, -13.3004, -13.18815, -13.07578, -12.96328, -12.85066, 
    -12.73791, -12.62503, -12.51203, -12.39891, -12.28566, -12.17228, 
    -12.05878, -11.94515, -11.8314, -11.71752, -11.60352, -11.4894, 
    -11.37515, -11.26078, -11.14628, -11.03166, -10.91691, -10.80205, 
    -10.68706, -10.57194, -10.45671, -10.34135, -10.22587, -10.11026, 
    -9.994539, -9.878692, -9.762722, -9.646631, -9.530419, -9.414086, 
    -9.297632, -9.181058, -9.064363, -8.947547, -8.830611, -8.713556, 
    -8.596381, -8.479087, -8.361673, -8.244142, -8.126491, -8.008722, 
    -7.890835, -7.77283, -7.654707, -7.536467, -7.41811, -7.299636, 
    -7.181046, -7.062339, -6.943516, -6.824578, -6.705524, -6.586355, 
    -6.467071, -6.347673, -6.22816, -6.108534, -5.988794, -5.86894, 
    -5.748974, -5.628895, -5.508703, -5.3884, -5.267984, -5.147458, -5.02682, 
    -4.906072, -4.785213, -4.664245, -4.543166, -4.421978, -4.300682, 
    -4.179276, -4.057763, -3.936141, -3.814413, -3.692577, -3.570634, 
    -3.448585, -3.32643, -3.20417, -3.081804, -2.959333, -2.836758, 
    -2.714079, -2.591297, -2.468411, -2.345423, -2.222332, -2.09914, 
    -1.975846, -1.85245, -1.728955, -1.605359, -1.481663, -1.357868, 
    -1.233974, -1.109982, -0.9858922, -0.8617046, -0.73742, -0.6130388, 
    -0.4885616, -0.3639887, -0.2393208, -0.1145581, 0.01029872, 0.1352492, 
    0.2602929, 0.3854293, 0.510658, 0.6359783, 0.7613898, 0.886892, 1.012484, 
    1.138166, 1.263938, 1.389798, 1.515746, 1.641781, 1.767904, 1.894113, 
    2.020408, 2.146788, 2.273254, 2.399804, 2.526437, 2.653154, 2.779953, 
    2.906835, 3.033798, 3.160842, 3.287967, 3.415171, 3.542455, 3.669817, 
    3.797257, 3.924775, 4.05237, 4.180041, 4.307788, 4.43561, 4.563507, 
    4.691478, 4.819521, 4.947638, 5.075827, 5.204087, 5.332418, 5.460819, 
    5.58929, 5.71783, 5.846438, 5.975114, 6.103857, 6.232666, 6.361542, 
    6.490482, 6.619487, 6.748556, 6.877688, 7.006883, 7.136139, 7.265457, 
    7.394835, 7.524273, 7.65377, 7.783326, 7.91294, 8.04261, 8.172338, 
    8.302121, 8.43196, 8.561852, 8.691799, 8.821799, 8.951852, 9.081955, 
    9.212111, 9.342316, 9.47257, 9.602874, 9.733226, 9.863626, 9.994071, 
    10.12456, 10.2551, 10.38568, 10.51631, 10.64698, 10.77769, 10.90844, 
    11.03924, 11.17007, 11.30095, 11.43186, 11.56281, 11.6938, 11.82483, 
    11.95589, 12.08698, 12.21811, 12.34928, 12.48047, 12.6117, 12.74296, 
    12.87426, 13.00558, 13.13693, 13.26831, 13.39971, 13.53115, 13.66261, 
    13.79409, 13.9256, 14.05713, 14.18869, 14.32027, 14.45187, 14.58349, 
    14.71513, 14.84679, 14.97847, 15.11017, 15.24188, 15.37361, 15.50536, 
    15.63712, 15.76889, 15.90068, 16.03248, 16.16429, 16.29611, 16.42795, 
    16.55979, 16.69164, 16.8235, 16.95536, 17.08723, 17.21911, 17.35099, 
    17.48287, 17.61476, 17.74665, 17.87854, 18.01043, 18.14232, 18.27421, 
    18.4061, 18.53799, 18.66987, 18.80175, 18.93363, 19.0655, 19.19736, 
    19.32922, 19.46107, 19.59291, 19.72474, 19.85656, 19.98837, 20.12017, 
    20.25195, 20.38372, 20.51548, 20.64722, 20.77895, 20.91066, 21.04236, 
    21.17403, 21.30569, 21.43733, 21.56895, 21.70054, 21.83212, 21.96367, 
    22.0952, 22.22671, 22.35819, 22.48965, 22.62107, 22.75248, 22.88385, 
    23.0152, 23.14651, 23.2778, 23.40906, 23.54028, 23.67147, 23.80263, 
    23.93376, 24.06485, 24.1959, 24.32692, 24.4579, 24.58885, 24.71976, 
    24.85063, 24.98145, 25.11224, 25.24299, 25.37369, 25.50436, 25.63498, 
    25.76555, 25.89608, 26.02657, 26.15701, 26.2874, 26.41774, 26.54804, 
    26.67828, 26.80848, 26.93863, 27.06872, 27.19877, 27.32876, 27.4587, 
    27.58858, 27.71841, 27.84819, 27.97791, 28.10757, 28.23717, 28.36672, 
    28.49621, 28.62564, 28.755, 28.88431, 29.01356, 29.14274, 29.27187, 
    29.40092, 29.52992, 29.65885, 29.78771, 29.91651, 30.04524, 30.17391, 
    30.30251, 30.43104, 30.5595, 30.68789, 30.81621, 30.94446, 31.07263, 
    31.20074, 31.32877, 31.45673, 31.58461, 31.71242, 31.84016, 31.96782, 
    32.0954, 32.22291, 32.35033, 32.47768, 32.60496, 32.73215, 32.85926, 
    32.98629, 33.11324, 33.24011, 33.3669, 33.4936, 33.62022, 33.74676, 
    33.87321, 33.99958, 34.12586, 34.25205, 34.37816, 34.50418, 34.63012, 
    34.75596, 34.88172, 35.00739, 35.13297, 35.25845, 35.38385, 35.50916, 
    35.63437, 35.75949, 35.88452, 36.00946, 36.1343, 36.25905, 36.3837, 
    36.50826, 36.63272, 36.75709, 36.88136, 37.00553, 37.1296, 37.25358, 
    37.37746, 37.50124, 37.62492, 37.7485, 37.87197, 37.99535, 38.11863, 
    38.24181, 38.36488, 38.48786, 38.61073, 38.73349, 38.85616, 38.97871, 
    39.10117, 39.22351, 39.34576, 39.4679, 39.58993, 39.71186, 39.83368, 
    39.95539,
  -14.80298, -14.69224, -14.58137, -14.47038, -14.35926, -14.24801, 
    -14.13663, -14.02513, -13.9135, -13.80174, -13.68985, -13.57784, 
    -13.4657, -13.35343, -13.24104, -13.12852, -13.01587, -12.9031, -12.7902, 
    -12.67717, -12.56402, -12.45075, -12.33734, -12.22381, -12.11016, 
    -11.99638, -11.88247, -11.76844, -11.65429, -11.54001, -11.4256, 
    -11.31107, -11.19642, -11.08164, -10.96674, -10.85171, -10.73656, 
    -10.62129, -10.50589, -10.39037, -10.27473, -10.15896, -10.04307, 
    -9.927061, -9.810927, -9.694672, -9.578294, -9.461795, -9.345174, 
    -9.228432, -9.111568, -8.994584, -8.87748, -8.760255, -8.642909, 
    -8.525444, -8.40786, -8.290155, -8.172332, -8.054389, -7.936328, 
    -7.818149, -7.699851, -7.581435, -7.462902, -7.344251, -7.225483, 
    -7.106598, -6.987597, -6.86848, -6.749246, -6.629897, -6.510432, 
    -6.390852, -6.271157, -6.151348, -6.031425, -5.911387, -5.791236, 
    -5.670972, -5.550595, -5.430106, -5.309504, -5.188789, -5.067964, 
    -4.947027, -4.825979, -4.704821, -4.583552, -4.462173, -4.340686, 
    -4.219089, -4.097383, -3.975568, -3.853645, -3.731615, -3.609478, 
    -3.487233, -3.364882, -3.242425, -3.119863, -2.997194, -2.874421, 
    -2.751544, -2.628562, -2.505476, -2.382288, -2.258996, -2.135602, 
    -2.012106, -1.888508, -1.764809, -1.64101, -1.51711, -1.39311, -1.269011, 
    -1.144813, -1.020517, -0.8961222, -0.7716301, -0.647041, -0.5223553, 
    -0.3975734, -0.2726958, -0.1477231, -0.0226557, 0.1025059, 0.2277612, 
    0.3531098, 0.4785511, 0.6040846, 0.7297097, 0.8554261, 0.9812332, 
    1.10713, 1.233117, 1.359193, 1.485358, 1.611611, 1.737951, 1.864378, 
    1.990892, 2.117491, 2.244176, 2.370946, 2.4978, 2.624738, 2.751759, 
    2.878863, 3.006048, 3.133315, 3.260663, 3.388091, 3.515599, 3.643186, 
    3.770852, 3.898595, 4.026416, 4.154314, 4.282288, 4.410337, 4.538461, 
    4.66666, 4.794932, 4.923278, 5.051696, 5.180186, 5.308747, 5.437379, 
    5.566081, 5.694852, 5.823693, 5.952601, 6.081576, 6.210619, 6.339727, 
    6.468902, 6.598141, 6.727444, 6.856811, 6.986241, 7.115733, 7.245286, 
    7.374901, 7.504576, 7.63431, 7.764103, 7.893955, 8.023864, 8.15383, 
    8.283852, 8.413929, 8.544062, 8.674248, 8.804488, 8.93478, 9.065125, 
    9.19552, 9.325967, 9.456464, 9.587009, 9.717603, 9.848245, 9.978933, 
    10.10967, 10.24045, 10.37127, 10.50214, 10.63306, 10.76401, 10.89501, 
    11.02605, 11.15713, 11.28825, 11.41941, 11.55061, 11.68184, 11.81311, 
    11.94442, 12.07576, 12.20714, 12.33855, 12.47, 12.60147, 12.73298, 
    12.86452, 12.99609, 13.12769, 13.25931, 13.39097, 13.52265, 13.65436, 
    13.78609, 13.91785, 14.04963, 14.18144, 14.31327, 14.44512, 14.57699, 
    14.70888, 14.84079, 14.97272, 15.10467, 15.23663, 15.36861, 15.50061, 
    15.63262, 15.76464, 15.89668, 16.02873, 16.1608, 16.29287, 16.42495, 
    16.55704, 16.68914, 16.82125, 16.95337, 17.08549, 17.21762, 17.34975, 
    17.48189, 17.61403, 17.74617, 17.87831, 18.01045, 18.1426, 18.27474, 
    18.40688, 18.53902, 18.67115, 18.80328, 18.93541, 19.06753, 19.19964, 
    19.33175, 19.46385, 19.59594, 19.72802, 19.8601, 19.99216, 20.1242, 
    20.25624, 20.38826, 20.52027, 20.65227, 20.78424, 20.9162, 21.04815, 
    21.18007, 21.31198, 21.44387, 21.57574, 21.70759, 21.83941, 21.97121, 
    22.10299, 22.23475, 22.36648, 22.49818, 22.62986, 22.76151, 22.89313, 
    23.02472, 23.15629, 23.28782, 23.41933, 23.5508, 23.68224, 23.81364, 
    23.94502, 24.07635, 24.20765, 24.33892, 24.47015, 24.60134, 24.73249, 
    24.86361, 24.99468, 25.12571, 25.2567, 25.38765, 25.51856, 25.64942, 
    25.78024, 25.91101, 26.04174, 26.17242, 26.30306, 26.43365, 26.56418, 
    26.69467, 26.82511, 26.9555, 27.08583, 27.21612, 27.34635, 27.47653, 
    27.60665, 27.73672, 27.86673, 27.99669, 28.12659, 28.25643, 28.38622, 
    28.51594, 28.64561, 28.77521, 28.90475, 29.03424, 29.16366, 29.29301, 
    29.42231, 29.55154, 29.6807, 29.8098, 29.93883, 30.06779, 30.19669, 
    30.32552, 30.45428, 30.58297, 30.71159, 30.84014, 30.96862, 31.09703, 
    31.22536, 31.35362, 31.48181, 31.60992, 31.73796, 31.86592, 31.99381, 
    32.12162, 32.24935, 32.377, 32.50458, 32.63207, 32.75949, 32.88682, 
    33.01408, 33.14125, 33.26834, 33.39535, 33.52227, 33.64911, 33.77587, 
    33.90254, 34.02913, 34.15563, 34.28204, 34.40837, 34.53461, 34.66076, 
    34.78682, 34.91279, 35.03867, 35.16447, 35.29017, 35.41578, 35.5413, 
    35.66673, 35.79206, 35.9173, 36.04245, 36.1675, 36.29246, 36.41732, 
    36.54208, 36.66676, 36.79133, 36.91581, 37.04018, 37.16447, 37.28865, 
    37.41273, 37.53672, 37.6606, 37.78438, 37.90807, 38.03165, 38.15513, 
    38.27851, 38.40178, 38.52495, 38.64802, 38.77099, 38.89385, 39.01661, 
    39.13926, 39.2618, 39.38424, 39.50658, 39.62881, 39.75093, 39.87294, 
    39.99484,
  -14.85798, -14.7471, -14.63609, -14.52496, -14.41369, -14.3023, -14.19078, 
    -14.07914, -13.96736, -13.85546, -13.74343, -13.63127, -13.51898, 
    -13.40657, -13.29403, -13.18136, -13.06857, -12.95565, -12.8426, 
    -12.72942, -12.61612, -12.50269, -12.38914, -12.27546, -12.16165, 
    -12.04772, -11.93366, -11.81947, -11.70516, -11.59073, -11.47617, 
    -11.36148, -11.24667, -11.13173, -11.01667, -10.90148, -10.78617, 
    -10.67074, -10.55518, -10.4395, -10.32369, -10.20777, -10.09171, 
    -9.975537, -9.85924, -9.742818, -9.626275, -9.509609, -9.392821, 
    -9.275911, -9.15888, -9.041727, -8.924453, -8.807058, -8.689543, 
    -8.571906, -8.454149, -8.336273, -8.218277, -8.100161, -7.981925, 
    -7.863571, -7.745098, -7.626507, -7.507797, -7.388969, -7.270023, 
    -7.15096, -7.03178, -6.912483, -6.79307, -6.67354, -6.553894, -6.434132, 
    -6.314255, -6.194263, -6.074156, -5.953935, -5.833599, -5.71315, 
    -5.592587, -5.47191, -5.351121, -5.23022, -5.109206, -4.988081, 
    -4.866843, -4.745495, -4.624035, -4.502466, -4.380786, -4.258996, 
    -4.137098, -4.01509, -3.892973, -3.770749, -3.648416, -3.525976, 
    -3.403429, -3.280775, -3.158015, -3.035149, -2.912177, -2.7891, 
    -2.665919, -2.542634, -2.419244, -2.295751, -2.172155, -2.048457, 
    -1.924656, -1.800754, -1.67675, -1.552645, -1.428441, -1.304136, 
    -1.179732, -1.055228, -0.9306266, -0.8059268, -0.6811293, -0.5562347, 
    -0.4312433, -0.3061559, -0.1809727, -0.05569425, 0.0696789, 0.1951463, 
    0.3207074, 0.4463617, 0.5721088, 0.6979481, 0.8238791, 0.9499013, 
    1.076014, 1.202217, 1.32851, 1.454892, 1.581362, 1.70792, 1.834566, 
    1.961299, 2.088118, 2.215023, 2.342013, 2.469089, 2.596248, 2.723491, 
    2.850817, 2.978225, 3.105716, 3.233287, 3.36094, 3.488672, 3.616484, 
    3.744375, 3.872345, 4.000392, 4.128517, 4.256719, 4.384995, 4.513348, 
    4.641776, 4.770278, 4.898852, 5.027501, 5.156221, 5.285013, 5.413876, 
    5.542809, 5.671813, 5.800886, 5.930027, 6.059236, 6.188511, 6.317854, 
    6.447263, 6.576736, 6.706275, 6.835877, 6.965543, 7.095272, 7.225061, 
    7.354913, 7.484825, 7.614797, 7.744829, 7.874918, 8.005066, 8.135271, 
    8.265532, 8.395849, 8.526222, 8.656649, 8.787129, 8.917663, 9.048248, 
    9.178885, 9.309574, 9.440312, 9.5711, 9.701938, 9.832822, 9.963754, 
    10.09473, 10.22576, 10.35683, 10.48794, 10.6191, 10.7503, 10.88154, 
    11.01283, 11.14415, 11.27552, 11.40692, 11.53837, 11.66985, 11.80137, 
    11.93292, 12.06451, 12.19614, 12.32779, 12.45949, 12.59121, 12.72297, 
    12.85476, 12.98657, 13.11842, 13.2503, 13.3822, 13.51413, 13.64609, 
    13.77807, 13.91008, 14.04211, 14.17417, 14.30625, 14.43835, 14.57047, 
    14.70261, 14.83477, 14.96695, 15.09915, 15.23137, 15.3636, 15.49585, 
    15.62811, 15.76038, 15.89267, 16.02497, 16.15729, 16.28961, 16.42195, 
    16.55429, 16.68665, 16.81901, 16.95137, 17.08375, 17.21613, 17.34851, 
    17.4809, 17.61329, 17.74568, 17.87808, 18.01047, 18.14287, 18.27526, 
    18.40765, 18.54004, 18.67243, 18.80482, 18.93719, 19.06957, 19.20193, 
    19.33429, 19.46664, 19.59899, 19.73132, 19.86364, 19.99595, 20.12825, 
    20.26054, 20.39281, 20.52508, 20.65732, 20.78955, 20.92176, 21.05396, 
    21.18613, 21.31829, 21.45043, 21.58255, 21.71465, 21.84672, 21.97877, 
    22.1108, 22.24281, 22.37479, 22.50674, 22.63867, 22.77057, 22.90244, 
    23.03428, 23.16609, 23.29788, 23.42963, 23.56135, 23.69304, 23.82469, 
    23.95631, 24.08789, 24.21944, 24.35095, 24.48243, 24.61386, 24.74526, 
    24.87662, 25.00794, 25.13922, 25.27046, 25.40165, 25.5328, 25.66391, 
    25.79497, 25.92599, 26.05696, 26.18789, 26.31876, 26.44959, 26.58037, 
    26.7111, 26.84178, 26.97241, 27.10299, 27.23351, 27.36399, 27.4944, 
    27.62477, 27.75508, 27.88533, 28.01553, 28.14566, 28.27574, 28.40577, 
    28.53573, 28.66563, 28.79547, 28.92525, 29.05497, 29.18463, 29.31422, 
    29.44375, 29.57321, 29.70261, 29.83194, 29.96121, 30.09041, 30.21954, 
    30.3486, 30.47759, 30.60651, 30.73536, 30.86415, 30.99286, 31.12149, 
    31.25006, 31.37854, 31.50696, 31.6353, 31.76357, 31.89176, 32.01987, 
    32.1479, 32.27586, 32.40374, 32.53154, 32.65926, 32.7869, 32.91446, 
    33.04193, 33.16933, 33.29664, 33.42387, 33.55102, 33.67808, 33.80506, 
    33.93195, 34.05875, 34.18547, 34.31211, 34.43865, 34.56511, 34.69147, 
    34.81775, 34.94394, 35.07004, 35.19605, 35.32196, 35.44779, 35.57352, 
    35.69916, 35.82471, 35.95016, 36.07552, 36.20078, 36.32595, 36.45102, 
    36.576, 36.70088, 36.82566, 36.95034, 37.07493, 37.19942, 37.32381, 
    37.44809, 37.57228, 37.69637, 37.82036, 37.94424, 38.06803, 38.19171, 
    38.31529, 38.43877, 38.56214, 38.68541, 38.80857, 38.93164, 39.05459, 
    39.17744, 39.30018, 39.42282, 39.54535, 39.66777, 39.79009, 39.9123, 
    40.0344,
  -14.91309, -14.80207, -14.69092, -14.57965, -14.46824, -14.35671, 
    -14.24505, -14.13326, -14.02134, -13.90929, -13.79712, -13.68481, 
    -13.57238, -13.45982, -13.34713, -13.23432, -13.12138, -13.00831, 
    -12.89511, -12.78178, -12.66833, -12.55475, -12.44104, -12.32721, 
    -12.21325, -12.09916, -11.98495, -11.87061, -11.75615, -11.64155, 
    -11.52684, -11.41199, -11.29702, -11.18193, -11.06671, -10.95136, 
    -10.83589, -10.7203, -10.60458, -10.48874, -10.37277, -10.25668, 
    -10.14046, -10.02412, -9.907658, -9.791072, -9.674362, -9.557529, 
    -9.440575, -9.323498, -9.206298, -9.088976, -8.971533, -8.853968, 
    -8.73628, -8.618473, -8.500545, -8.382496, -8.264326, -8.146037, 
    -8.027627, -7.909098, -7.79045, -7.671682, -7.552795, -7.43379, 
    -7.314667, -7.195426, -7.076066, -6.95659, -6.836996, -6.717285, 
    -6.597458, -6.477514, -6.357455, -6.237279, -6.116989, -5.996583, 
    -5.876062, -5.755427, -5.634678, -5.513815, -5.392838, -5.271749, 
    -5.150547, -5.029232, -4.907805, -4.786267, -4.664617, -4.542856, 
    -4.420984, -4.299002, -4.17691, -4.054708, -3.932398, -3.809978, 
    -3.68745, -3.564814, -3.44207, -3.319219, -3.196261, -3.073197, 
    -2.950027, -2.82675, -2.703369, -2.579883, -2.456292, -2.332598, -2.2088, 
    -2.084898, -1.960894, -1.836788, -1.71258, -1.588271, -1.46386, 
    -1.339349, -1.214739, -1.090028, -0.9652187, -0.8403106, -0.7153043, 
    -0.5902004, -0.4649993, -0.3397014, -0.2143073, -0.08881748, 0.03676761, 
    0.1624475, 0.2882216, 0.4140894, 0.5400505, 0.6661043, 0.7922504, 
    0.9184881, 1.044817, 1.171237, 1.297746, 1.424346, 1.551034, 1.677811, 
    1.804676, 1.931628, 2.058668, 2.185793, 2.313004, 2.440301, 2.567683, 
    2.695148, 2.822697, 2.950328, 3.078043, 3.205839, 3.333716, 3.461674, 
    3.589712, 3.717829, 3.846025, 3.9743, 4.102652, 4.231081, 4.359587, 
    4.488168, 4.616825, 4.745556, 4.874362, 5.00324, 5.132191, 5.261215, 
    5.39031, 5.519475, 5.648711, 5.778017, 5.907391, 6.036834, 6.166344, 
    6.295921, 6.425565, 6.555274, 6.685048, 6.814887, 6.944789, 7.074754, 
    7.204782, 7.33487, 7.465021, 7.595231, 7.725501, 7.855829, 7.986217, 
    8.116661, 8.247162, 8.37772, 8.508333, 8.639001, 8.769722, 8.900497, 
    9.031325, 9.162205, 9.293136, 9.424117, 9.555148, 9.686228, 9.817356, 
    9.948532, 10.07976, 10.21102, 10.34234, 10.4737, 10.6051, 10.73655, 
    10.86804, 10.99957, 11.13114, 11.26275, 11.3944, 11.52609, 11.65782, 
    11.78959, 11.92139, 12.05323, 12.1851, 12.31701, 12.44895, 12.58092, 
    12.71293, 12.84496, 12.97703, 13.10913, 13.24125, 13.37341, 13.50559, 
    13.6378, 13.77003, 13.90229, 14.03457, 14.16688, 14.29921, 14.43156, 
    14.56393, 14.69633, 14.82874, 14.96117, 15.09362, 15.22609, 15.35857, 
    15.49107, 15.62358, 15.75611, 15.88865, 16.02121, 16.15377, 16.28635, 
    16.41894, 16.55153, 16.68414, 16.81675, 16.94937, 17.082, 17.21463, 
    17.34727, 17.47991, 17.61255, 17.7452, 17.87784, 18.01049, 18.14314, 
    18.27579, 18.40843, 18.54107, 18.67372, 18.80635, 18.93898, 19.07161, 
    19.20423, 19.33684, 19.46944, 19.60204, 19.73462, 19.8672, 19.99976, 
    20.13231, 20.26485, 20.39738, 20.52989, 20.66239, 20.79487, 20.92733, 
    21.05978, 21.19221, 21.32462, 21.45701, 21.58938, 21.72173, 21.85405, 
    21.98635, 22.11863, 22.25089, 22.38312, 22.51532, 22.6475, 22.77965, 
    22.91177, 23.04386, 23.17592, 23.30796, 23.43996, 23.57193, 23.70386, 
    23.83576, 23.96763, 24.09946, 24.23126, 24.36302, 24.49474, 24.62642, 
    24.75807, 24.88968, 25.02124, 25.15277, 25.28425, 25.41569, 25.54708, 
    25.67844, 25.80974, 25.94101, 26.07222, 26.20339, 26.33451, 26.46558, 
    26.59661, 26.72758, 26.8585, 26.98937, 27.12019, 27.25096, 27.38167, 
    27.51233, 27.64294, 27.77349, 27.90398, 28.03441, 28.16479, 28.29511, 
    28.42537, 28.55557, 28.68571, 28.81579, 28.94581, 29.07576, 29.20566, 
    29.33548, 29.46525, 29.59495, 29.72458, 29.85415, 29.98365, 30.11308, 
    30.24244, 30.37174, 30.50096, 30.63012, 30.7592, 30.88821, 31.01715, 
    31.14602, 31.27481, 31.40353, 31.53218, 31.66075, 31.78924, 31.91766, 
    32.046, 32.17426, 32.30244, 32.43055, 32.55857, 32.68652, 32.81438, 
    32.94217, 33.06987, 33.19749, 33.32502, 33.45247, 33.57984, 33.70712, 
    33.83432, 33.96143, 34.08846, 34.2154, 34.34225, 34.46901, 34.59569, 
    34.72227, 34.84877, 34.97517, 35.10149, 35.22771, 35.35384, 35.47988, 
    35.60583, 35.73168, 35.85744, 35.9831, 36.10867, 36.23415, 36.35953, 
    36.48481, 36.61, 36.73508, 36.86008, 36.98497, 37.10976, 37.23446, 
    37.35905, 37.48355, 37.60794, 37.73223, 37.85643, 37.98052, 38.1045, 
    38.22839, 38.35217, 38.47585, 38.59942, 38.72289, 38.84626, 38.96952, 
    39.09267, 39.21572, 39.33866, 39.46149, 39.58422, 39.70684, 39.82935, 
    39.95175, 40.07405,
  -14.96831, -14.85715, -14.74586, -14.63444, -14.5229, -14.41122, -14.29942, 
    -14.18749, -14.07543, -13.96323, -13.85091, -13.73847, -13.62589, 
    -13.51318, -13.40035, -13.28738, -13.17429, -13.06108, -12.94773, 
    -12.83425, -12.72065, -12.60692, -12.49306, -12.37907, -12.26496, 
    -12.15072, -12.03635, -11.92186, -11.80724, -11.69249, -11.57762, 
    -11.46262, -11.34749, -11.23224, -11.11686, -11.00135, -10.88572, 
    -10.76997, -10.65409, -10.53808, -10.42195, -10.3057, -10.18932, 
    -10.07281, -9.956184, -9.839433, -9.722557, -9.605557, -9.488436, 
    -9.37119, -9.253822, -9.136332, -9.018718, -8.900983, -8.783126, 
    -8.665147, -8.547046, -8.428824, -8.310481, -8.192018, -8.073434, 
    -7.95473, -7.835906, -7.716962, -7.597898, -7.478716, -7.359415, 
    -7.239995, -7.120456, -7.000799, -6.881025, -6.761133, -6.641124, 
    -6.520998, -6.400756, -6.280397, -6.159923, -6.039332, -5.918626, 
    -5.797805, -5.67687, -5.55582, -5.434656, -5.313378, -5.191987, 
    -5.070483, -4.948866, -4.827137, -4.705296, -4.583344, -4.461279, 
    -4.339105, -4.216819, -4.094424, -3.971918, -3.849303, -3.72658, 
    -3.603747, -3.480807, -3.357758, -3.234602, -3.111339, -2.98797, 
    -2.864494, -2.740912, -2.617225, -2.493433, -2.369537, -2.245536, 
    -2.121431, -1.997224, -1.872913, -1.7485, -1.623986, -1.499369, 
    -1.374652, -1.249834, -1.124916, -0.9998989, -0.8747821, -0.7495667, 
    -0.624253, -0.4988416, -0.373333, -0.2477276, -0.1220259, 0.003771531, 
    0.1296643, 0.2556518, 0.3817336, 0.5079092, 0.634178, 0.7605395, 
    0.8869933, 1.013539, 1.140175, 1.266903, 1.39372, 1.520627, 1.647623, 
    1.774707, 1.90188, 2.02914, 2.156486, 2.283919, 2.411438, 2.539042, 
    2.66673, 2.794502, 2.922358, 3.050296, 3.178317, 3.30642, 3.434603, 
    3.562867, 3.691211, 3.819635, 3.948137, 4.076717, 4.205375, 4.334109, 
    4.46292, 4.591806, 4.720768, 4.849804, 4.978914, 5.108097, 5.237352, 
    5.366679, 5.496078, 5.625547, 5.755086, 5.884694, 6.014371, 6.144116, 
    6.273929, 6.403808, 6.533753, 6.663763, 6.793839, 6.923978, 7.05418, 
    7.184445, 7.314773, 7.445161, 7.57561, 7.70612, 7.836688, 7.967315, 
    8.098, 8.228742, 8.35954, 8.490395, 8.621304, 8.752267, 8.883285, 
    9.014355, 9.145477, 9.276651, 9.407876, 9.53915, 9.670475, 9.801847, 
    9.933269, 10.06474, 10.19625, 10.32781, 10.45942, 10.59106, 10.72276, 
    10.85449, 10.98627, 11.11809, 11.24995, 11.38185, 11.51379, 11.64576, 
    11.77777, 11.90983, 12.04191, 12.17403, 12.30619, 12.43838, 12.5706, 
    12.70286, 12.83514, 12.96746, 13.09981, 13.23218, 13.36459, 13.49702, 
    13.62948, 13.76196, 13.89447, 14.02701, 14.15957, 14.29215, 14.42475, 
    14.55737, 14.69002, 14.82268, 14.95537, 15.08807, 15.22079, 15.35353, 
    15.48628, 15.61904, 15.75182, 15.88462, 16.01743, 16.15025, 16.28308, 
    16.41592, 16.54877, 16.68162, 16.81449, 16.94736, 17.08024, 17.21313, 
    17.34602, 17.47891, 17.61181, 17.74471, 17.87761, 18.01051, 18.14341, 
    18.27631, 18.40921, 18.54211, 18.675, 18.80789, 18.94078, 19.07366, 
    19.20653, 19.33939, 19.47225, 19.6051, 19.73794, 19.87077, 20.00358, 
    20.13639, 20.26918, 20.40196, 20.53472, 20.66747, 20.80021, 20.93292, 
    21.06562, 21.1983, 21.33096, 21.46361, 21.59623, 21.72883, 21.8614, 
    21.99396, 22.12649, 22.259, 22.39148, 22.52393, 22.65636, 22.78876, 
    22.92113, 23.05347, 23.18578, 23.31807, 23.45032, 23.58253, 23.71472, 
    23.84687, 23.97898, 24.11106, 24.24311, 24.37512, 24.50709, 24.63902, 
    24.77091, 24.90277, 25.03458, 25.16635, 25.29808, 25.42976, 25.56141, 
    25.693, 25.82456, 25.95606, 26.08752, 26.21894, 26.3503, 26.48162, 
    26.61288, 26.7441, 26.87527, 27.00638, 27.13744, 27.26845, 27.39941, 
    27.53031, 27.66115, 27.79194, 27.92268, 28.05335, 28.18397, 28.31453, 
    28.44503, 28.57547, 28.70585, 28.83616, 28.96642, 29.09661, 29.22674, 
    29.35681, 29.48681, 29.61674, 29.74661, 29.87641, 30.00615, 30.13581, 
    30.26541, 30.39494, 30.52439, 30.65378, 30.7831, 30.91234, 31.04151, 
    31.17061, 31.29964, 31.42859, 31.55746, 31.68626, 31.81498, 31.94363, 
    32.0722, 32.20068, 32.32909, 32.45743, 32.58568, 32.71385, 32.84194, 
    32.96995, 33.09787, 33.22572, 33.35347, 33.48115, 33.60874, 33.73624, 
    33.86366, 33.991, 34.11824, 34.2454, 34.37247, 34.49945, 34.62635, 
    34.75315, 34.87986, 35.00648, 35.13301, 35.25946, 35.3858, 35.51205, 
    35.63822, 35.76428, 35.89025, 36.01613, 36.14192, 36.2676, 36.39319, 
    36.51869, 36.64408, 36.76938, 36.89458, 37.01968, 37.14468, 37.26958, 
    37.39439, 37.51909, 37.64369, 37.76819, 37.89259, 38.01688, 38.14107, 
    38.26516, 38.38914, 38.51302, 38.6368, 38.76047, 38.88403, 39.00749, 
    39.13084, 39.25409, 39.37723, 39.50026, 39.62318, 39.746, 39.86871, 
    39.9913, 40.11379,
  -15.02363, -14.91234, -14.80091, -14.68935, -14.57767, -14.46585, -14.3539, 
    -14.24183, -14.12962, -14.01729, -13.90482, -13.79223, -13.67951, 
    -13.56665, -13.45367, -13.34056, -13.22732, -13.11395, -13.00046, 
    -12.88683, -12.77308, -12.6592, -12.54519, -12.43105, -12.31678, 
    -12.20239, -12.08787, -11.97322, -11.85844, -11.74354, -11.62851, 
    -11.51335, -11.39806, -11.28265, -11.16711, -11.05145, -10.93566, 
    -10.81974, -10.7037, -10.58753, -10.47124, -10.35482, -10.23828, 
    -10.12161, -10.00482, -9.887901, -9.77086, -9.653693, -9.536404, 
    -9.418991, -9.301454, -9.183794, -9.06601, -8.948105, -8.830077, 
    -8.711926, -8.593654, -8.475259, -8.356743, -8.238105, -8.119347, 
    -8.000467, -7.881467, -7.762347, -7.643106, -7.523746, -7.404266, 
    -7.284667, -7.164949, -7.045113, -6.925158, -6.805085, -6.684894, 
    -6.564586, -6.44416, -6.323617, -6.202959, -6.082183, -5.961292, 
    -5.840285, -5.719163, -5.597926, -5.476574, -5.355108, -5.233528, 
    -5.111834, -4.990027, -4.868107, -4.746075, -4.62393, -4.501674, 
    -4.379305, -4.256826, -4.134236, -4.011536, -3.888726, -3.765806, 
    -3.642777, -3.519639, -3.396393, -3.273039, -3.149577, -3.026008, 
    -2.902332, -2.778549, -2.654661, -2.530667, -2.406568, -2.282365, 
    -2.158057, -2.033645, -1.90913, -1.784512, -1.659791, -1.534969, 
    -1.410045, -1.28502, -1.159894, -1.034668, -0.9093419, -0.7839169, 
    -0.6583931, -0.5327711, -0.4070512, -0.2812341, -0.1553202, -0.0293099, 
    0.09679617, 0.2229975, 0.3492937, 0.4756842, 0.6021684, 0.728746, 
    0.8554162, 0.9821787, 1.109033, 1.235978, 1.363014, 1.49014, 1.617355, 
    1.74466, 1.872053, 1.999534, 2.127102, 2.254757, 2.382498, 2.510324, 
    2.638236, 2.766232, 2.894312, 3.022476, 3.150722, 3.279051, 3.40746, 
    3.535951, 3.664523, 3.793174, 3.921904, 4.050713, 4.179599, 4.308563, 
    4.437604, 4.56672, 4.695913, 4.82518, 4.954522, 5.083936, 5.213424, 
    5.342984, 5.472616, 5.602319, 5.732092, 5.861935, 5.991847, 6.121828, 
    6.251875, 6.381991, 6.512172, 6.64242, 6.772732, 6.903109, 7.03355, 
    7.164053, 7.29462, 7.425247, 7.555936, 7.686685, 7.817493, 7.94836, 
    8.079287, 8.21027, 8.34131, 8.472405, 8.603558, 8.734763, 8.866023, 
    8.997337, 9.128703, 9.26012, 9.391589, 9.523108, 9.654677, 9.786295, 
    9.917961, 10.04967, 10.18143, 10.31324, 10.44509, 10.57699, 10.70893, 
    10.84091, 10.97294, 11.105, 11.23711, 11.36926, 11.50144, 11.63367, 
    11.76593, 11.89823, 12.03057, 12.16294, 12.29534, 12.42778, 12.56026, 
    12.69276, 12.8253, 12.95786, 13.09046, 13.22309, 13.35575, 13.48843, 
    13.62114, 13.75388, 13.88664, 14.01942, 14.15223, 14.28507, 14.41792, 
    14.5508, 14.6837, 14.81661, 14.94955, 15.08251, 15.21548, 15.34847, 
    15.48147, 15.61449, 15.74753, 15.88058, 16.01364, 16.14671, 16.27979, 
    16.41289, 16.54599, 16.6791, 16.81222, 16.94535, 17.07848, 17.21162, 
    17.34477, 17.47792, 17.61107, 17.74422, 17.87738, 18.01053, 18.14369, 
    18.27684, 18.41, 18.54315, 18.67629, 18.80944, 18.94258, 19.07571, 
    19.20884, 19.34196, 19.47507, 19.60817, 19.74126, 19.87434, 20.00741, 
    20.14047, 20.27352, 20.40655, 20.53957, 20.67257, 20.80556, 20.93853, 
    21.07148, 21.20441, 21.33733, 21.47022, 21.60309, 21.73595, 21.86878, 
    22.00158, 22.13437, 22.26712, 22.39986, 22.53256, 22.66524, 22.79789, 
    22.93051, 23.06311, 23.19567, 23.3282, 23.4607, 23.59317, 23.72561, 
    23.85801, 23.99037, 24.1227, 24.255, 24.38725, 24.51947, 24.65165, 
    24.78379, 24.91589, 25.04795, 25.17997, 25.31194, 25.44388, 25.57577, 
    25.70761, 25.83941, 25.97116, 26.10287, 26.23453, 26.36614, 26.4977, 
    26.62921, 26.76067, 26.89208, 27.02344, 27.15474, 27.286, 27.41719, 
    27.54834, 27.67942, 27.81045, 27.94143, 28.07234, 28.2032, 28.334, 
    28.46474, 28.59542, 28.72604, 28.85659, 28.98709, 29.11752, 29.24788, 
    29.37819, 29.50842, 29.6386, 29.7687, 29.89874, 30.02871, 30.15861, 
    30.28844, 30.4182, 30.54789, 30.67752, 30.80706, 30.93654, 31.06594, 
    31.19527, 31.32453, 31.45371, 31.58281, 31.71184, 31.84079, 31.96967, 
    32.09846, 32.22718, 32.35582, 32.48438, 32.61286, 32.74125, 32.86957, 
    32.9978, 33.12595, 33.25402, 33.382, 33.5099, 33.63771, 33.76544, 
    33.89308, 34.02064, 34.14811, 34.27548, 34.40277, 34.52998, 34.65709, 
    34.78411, 34.91104, 35.03788, 35.16463, 35.29128, 35.41785, 35.54432, 
    35.67069, 35.79697, 35.92316, 36.04925, 36.17524, 36.30114, 36.42694, 
    36.55265, 36.67826, 36.80376, 36.92917, 37.05448, 37.1797, 37.3048, 
    37.42981, 37.55472, 37.67953, 37.80423, 37.92883, 38.05333, 38.17773, 
    38.30202, 38.4262, 38.55029, 38.67427, 38.79814, 38.9219, 39.04556, 
    39.16911, 39.29256, 39.4159, 39.53912, 39.66225, 39.78526, 39.90816, 
    40.03095, 40.15364,
  -15.07908, -14.96764, -14.85607, -14.74438, -14.63255, -14.52059, -14.4085, 
    -14.29628, -14.18393, -14.07145, -13.95884, -13.8461, -13.73323, 
    -13.62024, -13.50711, -13.39385, -13.28046, -13.16694, -13.0533, 
    -12.93952, -12.82562, -12.71159, -12.59742, -12.48313, -12.36871, 
    -12.25417, -12.13949, -12.02468, -11.90975, -11.79469, -11.67951, 
    -11.56419, -11.44875, -11.33318, -11.21748, -11.10166, -10.98571, 
    -10.86963, -10.75343, -10.6371, -10.52064, -10.40406, -10.28735, 
    -10.17052, -10.05356, -9.936479, -9.819271, -9.701938, -9.584481, 
    -9.466899, -9.349194, -9.231364, -9.113411, -8.995335, -8.877135, 
    -8.758813, -8.640368, -8.5218, -8.403111, -8.284299, -8.165365, -8.04631, 
    -7.927134, -7.807837, -7.688419, -7.568882, -7.449224, -7.329445, 
    -7.209548, -7.089531, -6.969395, -6.84914, -6.728767, -6.608276, 
    -6.487668, -6.366941, -6.246098, -6.125137, -6.00406, -5.882867, 
    -5.761558, -5.640133, -5.518593, -5.396938, -5.275169, -5.153286, 
    -5.031288, -4.909177, -4.786953, -4.664616, -4.542167, -4.419605, 
    -4.296932, -4.174148, -4.051252, -3.928246, -3.80513, -3.681904, 
    -3.558568, -3.435124, -3.311571, -3.18791, -3.064141, -2.940264, 
    -2.816281, -2.692191, -2.567995, -2.443693, -2.319287, -2.194775, 
    -2.070159, -1.945439, -1.820615, -1.695688, -1.570659, -1.445528, 
    -1.320295, -1.194961, -1.069526, -0.9439905, -0.8183555, -0.6926212, 
    -0.5667881, -0.4408567, -0.3148274, -0.1887007, -0.06247725, 0.06384259, 
    0.1902583, 0.3167693, 0.4433751, 0.5700752, 0.6968691, 0.8237563, 
    0.9507362, 1.077808, 1.204972, 1.332227, 1.459572, 1.587008, 1.714533, 
    1.842147, 1.969849, 2.097639, 2.225517, 2.353481, 2.481531, 2.609666, 
    2.737887, 2.866192, 2.994581, 3.123053, 3.251608, 3.380244, 3.508963, 
    3.637762, 3.766641, 3.8956, 4.024638, 4.153754, 4.282948, 4.412219, 
    4.541567, 4.67099, 4.800489, 4.930063, 5.059711, 5.189431, 5.319225, 
    5.44909, 5.579028, 5.709035, 5.839114, 5.969261, 6.099477, 6.229762, 
    6.360114, 6.490532, 6.621017, 6.751568, 6.882183, 7.012862, 7.143605, 
    7.27441, 7.405278, 7.536206, 7.667196, 7.798245, 7.929354, 8.060521, 
    8.191746, 8.323029, 8.454367, 8.585761, 8.717211, 8.848714, 8.980271, 
    9.111881, 9.243544, 9.375257, 9.507022, 9.638836, 9.7707, 9.902612, 
    10.03457, 10.16658, 10.29863, 10.43073, 10.56287, 10.69506, 10.82729, 
    10.95956, 11.09188, 11.22423, 11.35663, 11.48906, 11.62154, 11.75405, 
    11.8866, 12.01919, 12.15181, 12.28446, 12.41715, 12.54988, 12.68263, 
    12.81542, 12.94824, 13.08109, 13.21397, 13.34688, 13.47981, 13.61277, 
    13.74576, 13.87878, 14.01182, 14.14488, 14.27797, 14.41107, 14.5442, 
    14.67736, 14.81053, 14.94372, 15.07693, 15.21015, 15.3434, 15.47665, 
    15.60993, 15.74322, 15.87652, 16.00983, 16.14316, 16.2765, 16.40985, 
    16.54321, 16.67657, 16.80995, 16.94333, 17.07672, 17.21011, 17.34351, 
    17.47692, 17.61032, 17.74373, 17.87714, 18.01055, 18.14396, 18.27737, 
    18.41078, 18.54419, 18.67759, 18.81099, 18.94438, 19.07777, 19.21115, 
    19.34452, 19.47789, 19.61125, 19.74459, 19.87793, 20.01126, 20.14457, 
    20.27787, 20.41115, 20.54443, 20.67768, 20.81092, 20.94415, 21.07735, 
    21.21054, 21.34371, 21.47686, 21.60998, 21.74309, 21.87617, 22.00923, 
    22.14227, 22.27527, 22.40826, 22.54122, 22.67415, 22.80705, 22.93993, 
    23.07277, 23.20559, 23.33837, 23.47112, 23.60384, 23.73652, 23.86917, 
    24.00179, 24.13437, 24.26691, 24.39942, 24.53189, 24.66432, 24.79671, 
    24.92906, 25.06136, 25.19363, 25.32585, 25.45803, 25.59017, 25.72226, 
    25.85431, 25.98631, 26.11826, 26.25016, 26.38202, 26.51382, 26.64558, 
    26.77729, 26.90894, 27.04054, 27.17209, 27.30359, 27.43503, 27.56641, 
    27.69774, 27.82902, 27.96023, 28.09139, 28.22249, 28.35353, 28.48451, 
    28.61543, 28.74628, 28.87708, 29.00781, 29.13848, 29.26909, 29.39963, 
    29.5301, 29.66051, 29.79085, 29.92113, 30.05133, 30.18147, 30.31153, 
    30.44153, 30.57146, 30.70131, 30.83109, 30.9608, 31.09044, 31.22, 
    31.34949, 31.4789, 31.60823, 31.73749, 31.86668, 31.99578, 32.12481, 
    32.25375, 32.38262, 32.5114, 32.64011, 32.76873, 32.89727, 33.02573, 
    33.15411, 33.2824, 33.41061, 33.53873, 33.66677, 33.79472, 33.92258, 
    34.05036, 34.17805, 34.30564, 34.43316, 34.56058, 34.68791, 34.81515, 
    34.9423, 35.06936, 35.19632, 35.32319, 35.44997, 35.57666, 35.70325, 
    35.82975, 35.95615, 36.08245, 36.20866, 36.33477, 36.46078, 36.5867, 
    36.71252, 36.83823, 36.96386, 37.08937, 37.21479, 37.34011, 37.46533, 
    37.59044, 37.71546, 37.84037, 37.96518, 38.08988, 38.21448, 38.33897, 
    38.46336, 38.58765, 38.71183, 38.8359, 38.95987, 39.08372, 39.20748, 
    39.33112, 39.45466, 39.57809, 39.7014, 39.82461, 39.94771, 40.0707, 
    40.19358,
  -15.13463, -15.02306, -14.91135, -14.79951, -14.68754, -14.57544, 
    -14.46321, -14.35085, -14.23835, -14.12573, -14.01297, -13.90009, 
    -13.78708, -13.67393, -13.56065, -13.44725, -13.33371, -13.22005, 
    -13.10625, -12.99232, -12.87827, -12.76408, -12.64977, -12.53533, 
    -12.42076, -12.30605, -12.19122, -12.07627, -11.96118, -11.84596, 
    -11.73062, -11.61514, -11.49954, -11.38382, -11.26796, -11.15198, 
    -11.03587, -10.91963, -10.80326, -10.68677, -10.57015, -10.45341, 
    -10.33654, -10.21954, -10.10242, -9.985166, -9.867791, -9.750292, 
    -9.632667, -9.514916, -9.397042, -9.279043, -9.16092, -9.042673, 
    -8.924302, -8.805808, -8.68719, -8.568449, -8.449586, -8.3306, -8.211491, 
    -8.09226, -7.972908, -7.853434, -7.733839, -7.614123, -7.494286, 
    -7.374329, -7.254251, -7.134054, -7.013737, -6.893301, -6.772745, 
    -6.652071, -6.531279, -6.410368, -6.28934, -6.168194, -6.046931, 
    -5.925551, -5.804055, -5.682443, -5.560715, -5.438871, -5.316912, 
    -5.194838, -5.07265, -4.950347, -4.827931, -4.705402, -4.582759, 
    -4.460004, -4.337137, -4.214157, -4.091066, -3.967864, -3.844551, 
    -3.721128, -3.597594, -3.473952, -3.350199, -3.226339, -3.10237, 
    -2.978292, -2.854108, -2.729816, -2.605417, -2.480913, -2.356302, 
    -2.231586, -2.106765, -1.98184, -1.85681, -1.731677, -1.606441, 
    -1.481102, -1.355661, -1.230118, -1.104474, -0.9787285, -0.8528832, 
    -0.7269379, -0.6008933, -0.4747498, -0.348508, -0.2221682, -0.09573106, 
    0.03080298, 0.1574334, 0.2841597, 0.4109813, 0.5378978, 0.6649085, 
    0.792013, 0.9192109, 1.046501, 1.173884, 1.301358, 1.428924, 1.55658, 
    1.684326, 1.812161, 1.940085, 2.068098, 2.196198, 2.324386, 2.45266, 
    2.58102, 2.709466, 2.837996, 2.966611, 3.095309, 3.224091, 3.352955, 
    3.481901, 3.610928, 3.740036, 3.869224, 3.998492, 4.127838, 4.257263, 
    4.386765, 4.516344, 4.645999, 4.775731, 4.905537, 5.035418, 5.165372, 
    5.2954, 5.4255, 5.555672, 5.685915, 5.816229, 5.946613, 6.077066, 
    6.207587, 6.338176, 6.468833, 6.599556, 6.730345, 6.861199, 6.992117, 
    7.123099, 7.254145, 7.385252, 7.516422, 7.647653, 7.778944, 7.910294, 
    8.041703, 8.173171, 8.304696, 8.436277, 8.567916, 8.699609, 8.831357, 
    8.963159, 9.095014, 9.22692, 9.358879, 9.49089, 9.62295, 9.755059, 
    9.887218, 10.01942, 10.15168, 10.28398, 10.41632, 10.54872, 10.68115, 
    10.81363, 10.94615, 11.07872, 11.21132, 11.34397, 11.47665, 11.60938, 
    11.74214, 11.87494, 12.00777, 12.14065, 12.27355, 12.4065, 12.53947, 
    12.67248, 12.80552, 12.93859, 13.07169, 13.20482, 13.33798, 13.47117, 
    13.60439, 13.73763, 13.8709, 14.00419, 14.13751, 14.27085, 14.40421, 
    14.53759, 14.671, 14.80442, 14.93787, 15.07133, 15.20481, 15.33831, 
    15.47182, 15.60535, 15.73889, 15.87245, 16.00602, 16.1396, 16.2732, 
    16.4068, 16.54041, 16.67404, 16.80767, 16.94131, 17.07495, 17.2086, 
    17.34225, 17.47591, 17.60958, 17.74324, 17.87691, 18.01057, 18.14424, 
    18.2779, 18.41157, 18.54523, 18.67889, 18.81254, 18.94619, 19.07983, 
    19.21347, 19.3471, 19.48072, 19.61433, 19.74794, 19.88153, 20.01511, 
    20.14868, 20.28223, 20.41577, 20.5493, 20.68281, 20.81631, 20.94978, 
    21.08324, 21.21668, 21.35011, 21.48351, 21.61689, 21.75025, 21.88358, 
    22.0169, 22.15019, 22.28345, 22.41669, 22.5499, 22.68308, 22.81624, 
    22.94937, 23.08246, 23.21553, 23.34856, 23.48157, 23.61454, 23.74747, 
    23.88037, 24.01324, 24.14607, 24.27887, 24.41162, 24.54434, 24.67702, 
    24.80966, 24.94226, 25.07481, 25.20733, 25.3398, 25.47223, 25.60461, 
    25.73695, 25.86925, 26.00149, 26.13369, 26.26584, 26.39794, 26.52999, 
    26.662, 26.79395, 26.92585, 27.05769, 27.18949, 27.32123, 27.45291, 
    27.58454, 27.71611, 27.84763, 27.97909, 28.11049, 28.24183, 28.37311, 
    28.50433, 28.63549, 28.76659, 28.89762, 29.0286, 29.1595, 29.29035, 
    29.42113, 29.55184, 29.68249, 29.81306, 29.94357, 30.07402, 30.20439, 
    30.33469, 30.46492, 30.59509, 30.72517, 30.85519, 30.98513, 31.115, 
    31.24479, 31.37452, 31.50416, 31.63373, 31.76322, 31.89263, 32.02196, 
    32.15121, 32.28039, 32.40949, 32.5385, 32.66743, 32.79629, 32.92505, 
    33.05374, 33.18234, 33.31086, 33.43929, 33.56764, 33.6959, 33.82407, 
    33.95216, 34.08015, 34.20807, 34.33589, 34.46362, 34.59126, 34.71881, 
    34.84627, 34.97364, 35.10092, 35.2281, 35.35519, 35.48219, 35.60909, 
    35.73589, 35.8626, 35.98922, 36.11574, 36.24216, 36.36848, 36.49471, 
    36.62084, 36.74687, 36.8728, 36.99863, 37.12436, 37.24998, 37.37551, 
    37.50093, 37.62626, 37.75148, 37.87659, 38.00161, 38.12652, 38.25132, 
    38.37602, 38.50061, 38.6251, 38.74949, 38.87376, 38.99792, 39.12199, 
    39.24594, 39.36978, 39.49352, 39.61714, 39.74066, 39.86406, 39.98736, 
    40.11055, 40.23362,
  -15.1903, -15.07858, -14.96673, -14.85476, -14.74265, -14.6304, -14.51803, 
    -14.40552, -14.29289, -14.18012, -14.06722, -13.95419, -13.84103, 
    -13.72774, -13.61431, -13.50076, -13.38708, -13.27326, -13.15932, 
    -13.04524, -12.93103, -12.8167, -12.70223, -12.58764, -12.47291, 
    -12.35806, -12.24307, -12.12796, -12.01271, -11.89734, -11.78184, 
    -11.66621, -11.55045, -11.43456, -11.31855, -11.20241, -11.08613, 
    -10.96974, -10.85321, -10.73655, -10.61977, -10.50286, -10.38583, 
    -10.26867, -10.15138, -10.03396, -9.916422, -9.798755, -9.680963, 
    -9.563044, -9.445001, -9.326832, -9.208538, -9.09012, -8.971578, 
    -8.852911, -8.73412, -8.615207, -8.496169, -8.377008, -8.257725, 
    -8.138318, -8.018789, -7.899138, -7.779366, -7.659471, -7.539455, 
    -7.419319, -7.299061, -7.178683, -7.058185, -6.937566, -6.816828, 
    -6.695971, -6.574995, -6.4539, -6.332687, -6.211355, -6.089906, 
    -5.968339, -5.846656, -5.724855, -5.602939, -5.480906, -5.358757, 
    -5.236492, -5.114113, -4.991619, -4.869011, -4.746288, -4.623452, 
    -4.500503, -4.377441, -4.254266, -4.13098, -4.007581, -3.884071, 
    -3.76045, -3.636719, -3.512877, -3.388925, -3.264865, -3.140695, 
    -3.016417, -2.89203, -2.767536, -2.642935, -2.518226, -2.393412, 
    -2.268491, -2.143465, -2.018334, -1.893098, -1.767758, -1.642315, 
    -1.516768, -1.391118, -1.265366, -1.139512, -1.013557, -0.8875004, 
    -0.7613438, -0.6350873, -0.5087313, -0.3822764, -0.2557231, -0.1290719, 
    -0.002323223, 0.1245224, 0.2514644, 0.3785022, 0.5056354, 0.6328635, 
    0.7601859, 0.8876021, 1.015111, 1.142714, 1.270408, 1.398194, 1.526071, 
    1.654038, 1.782095, 1.910242, 2.038478, 2.166802, 2.295213, 2.423712, 
    2.552297, 2.680968, 2.809724, 2.938565, 3.067491, 3.1965, 3.325592, 
    3.454766, 3.584022, 3.713359, 3.842777, 3.972275, 4.101852, 4.231508, 
    4.361241, 4.491053, 4.620941, 4.750905, 4.880944, 5.011059, 5.141247, 
    5.27151, 5.401845, 5.532252, 5.662732, 5.793282, 5.923902, 6.054592, 
    6.185351, 6.316178, 6.447073, 6.578034, 6.709063, 6.840156, 6.971314, 
    7.102537, 7.233823, 7.365171, 7.496583, 7.628055, 7.759588, 7.891181, 
    8.022833, 8.154543, 8.286312, 8.418138, 8.550019, 8.681957, 8.81395, 
    8.945996, 9.078097, 9.21025, 9.342455, 9.474711, 9.607018, 9.739375, 
    9.871781, 10.00424, 10.13674, 10.26929, 10.40188, 10.53452, 10.6672, 
    10.79993, 10.9327, 11.06552, 11.19837, 11.33127, 11.4642, 11.59718, 
    11.73019, 11.86324, 11.99633, 12.12945, 12.26261, 12.39581, 12.52903, 
    12.66229, 12.79559, 12.92891, 13.06227, 13.19565, 13.32906, 13.46251, 
    13.59597, 13.72947, 13.86299, 13.99654, 14.13011, 14.2637, 14.39732, 
    14.53096, 14.66462, 14.7983, 14.932, 15.06572, 15.19945, 15.33321, 
    15.46698, 15.60076, 15.73456, 15.86837, 16.0022, 16.13604, 16.26989, 
    16.40375, 16.53762, 16.6715, 16.80538, 16.93928, 17.07318, 17.20708, 
    17.34099, 17.47491, 17.60883, 17.74275, 17.87667, 18.01059, 18.14452, 
    18.27844, 18.41236, 18.54627, 18.68019, 18.8141, 18.94801, 19.08191, 
    19.2158, 19.34968, 19.48356, 19.61743, 19.75129, 19.88514, 20.01897, 
    20.1528, 20.28661, 20.4204, 20.55419, 20.68795, 20.8217, 20.95544, 
    21.08915, 21.22285, 21.35653, 21.49018, 21.62382, 21.75743, 21.89102, 
    22.02459, 22.15813, 22.29165, 22.42514, 22.55861, 22.69204, 22.82545, 
    22.95883, 23.09218, 23.2255, 23.35879, 23.49204, 23.62527, 23.75845, 
    23.89161, 24.02472, 24.15781, 24.29085, 24.42386, 24.55683, 24.68976, 
    24.82265, 24.9555, 25.0883, 25.22107, 25.35379, 25.48647, 25.6191, 
    25.75168, 25.88423, 26.01672, 26.14917, 26.28156, 26.41391, 26.54621, 
    26.67846, 26.81066, 26.9428, 27.07489, 27.20693, 27.33892, 27.47085, 
    27.60272, 27.73454, 27.86629, 27.998, 28.12964, 28.26122, 28.39275, 
    28.52421, 28.65561, 28.78695, 28.91822, 29.04944, 29.18059, 29.31167, 
    29.44269, 29.57364, 29.70452, 29.83534, 29.96609, 30.09677, 30.22737, 
    30.35791, 30.48838, 30.61878, 30.7491, 30.87935, 31.00953, 31.13963, 
    31.26966, 31.39961, 31.52949, 31.65929, 31.78901, 31.91865, 32.04821, 
    32.1777, 32.30711, 32.43643, 32.56567, 32.69484, 32.82391, 32.95291, 
    33.08182, 33.21065, 33.33939, 33.46805, 33.59662, 33.72511, 33.8535, 
    33.98181, 34.11003, 34.23817, 34.36621, 34.49416, 34.62202, 34.7498, 
    34.87748, 35.00507, 35.13256, 35.25996, 35.38727, 35.51448, 35.6416, 
    35.76862, 35.89555, 36.02238, 36.14911, 36.27575, 36.40229, 36.52872, 
    36.65507, 36.78131, 36.90745, 37.03349, 37.15943, 37.28526, 37.411, 
    37.53663, 37.66217, 37.78759, 37.91291, 38.03814, 38.16325, 38.28826, 
    38.41316, 38.53796, 38.66265, 38.78724, 38.91171, 39.03608, 39.16034, 
    39.2845, 39.40854, 39.53247, 39.6563, 39.78001, 39.90361, 40.02711, 
    40.15049, 40.27376,
  -15.24608, -15.13422, -15.02224, -14.91012, -14.79786, -14.68548, 
    -14.57296, -14.46031, -14.34754, -14.23462, -14.12158, -14.0084, 
    -13.8951, -13.78166, -13.66809, -13.55439, -13.44055, -13.32659, 
    -13.21249, -13.09827, -12.98391, -12.86942, -12.75481, -12.64006, 
    -12.52518, -12.41017, -12.29503, -12.17976, -12.06436, -11.94883, 
    -11.83318, -11.71739, -11.60147, -11.48543, -11.36925, -11.25295, 
    -11.13652, -11.01996, -10.90327, -10.78645, -10.66951, -10.55243, 
    -10.43523, -10.31791, -10.20045, -10.08287, -9.965163, -9.847329, 
    -9.729368, -9.611281, -9.493069, -9.37473, -9.256266, -9.137677, 
    -9.018963, -8.900124, -8.78116, -8.662073, -8.542861, -8.423526, 
    -8.304067, -8.184484, -8.064778, -7.94495, -7.824999, -7.704926, 
    -7.584732, -7.464415, -7.343977, -7.223418, -7.102738, -6.981938, 
    -6.861017, -6.739976, -6.618816, -6.497537, -6.376138, -6.254621, 
    -6.132985, -6.011231, -5.88936, -5.767371, -5.645266, -5.523043, 
    -5.400704, -5.278249, -5.155678, -5.032992, -4.910192, -4.787276, 
    -4.664246, -4.541102, -4.417846, -4.294475, -4.170992, -4.047397, 
    -3.92369, -3.799871, -3.675941, -3.5519, -3.427749, -3.303488, -3.179117, 
    -3.054637, -2.930049, -2.805352, -2.680547, -2.555635, -2.430617, 
    -2.305491, -2.180259, -2.054922, -1.92948, -1.803932, -1.678281, 
    -1.552525, -1.426667, -1.300705, -1.174641, -1.048475, -0.9222078, 
    -0.7958394, -0.6693705, -0.5428017, -0.4161334, -0.2893661, -0.1625003, 
    -0.03553658, 0.09152463, 0.2186828, 0.3459373, 0.4732878, 0.6007336, 
    0.7282743, 0.8559093, 0.9836381, 1.11146, 1.239375, 1.367381, 1.49548, 
    1.623669, 1.751949, 1.880319, 2.008778, 2.137326, 2.265962, 2.394685, 
    2.523496, 2.652393, 2.781376, 2.910444, 3.039597, 3.168834, 3.298154, 
    3.427557, 3.557043, 3.68661, 3.816258, 3.945986, 4.075794, 4.205682, 
    4.335648, 4.465692, 4.595812, 4.72601, 4.856284, 4.986632, 5.117056, 
    5.247553, 5.378124, 5.508768, 5.639483, 5.77027, 5.901128, 6.032056, 
    6.163053, 6.294118, 6.425252, 6.556453, 6.687721, 6.819055, 6.950453, 
    7.081917, 7.213444, 7.345034, 7.476687, 7.608402, 7.740178, 7.872014, 
    8.003909, 8.135863, 8.267876, 8.399946, 8.532073, 8.664256, 8.796494, 
    8.928786, 9.061133, 9.193532, 9.325984, 9.458488, 9.591042, 9.723646, 
    9.8563, 9.989002, 10.12175, 10.25455, 10.38739, 10.52028, 10.65322, 
    10.78619, 10.91922, 11.05228, 11.18539, 11.31853, 11.45172, 11.58494, 
    11.71821, 11.85151, 11.98485, 12.11823, 12.25164, 12.38509, 12.51857, 
    12.65208, 12.78563, 12.9192, 13.05281, 13.18645, 13.32012, 13.45381, 
    13.58754, 13.72129, 13.85506, 13.98887, 14.12269, 14.25654, 14.39041, 
    14.52431, 14.65822, 14.79216, 14.92611, 15.06009, 15.19408, 15.32809, 
    15.46212, 15.59616, 15.73021, 15.86428, 15.99836, 16.13246, 16.26657, 
    16.40068, 16.53481, 16.66894, 16.80309, 16.93724, 17.0714, 17.20556, 
    17.33973, 17.4739, 17.60808, 17.74225, 17.87643, 18.01061, 18.14479, 
    18.27897, 18.41315, 18.54732, 18.6815, 18.81566, 18.94983, 19.08398, 
    19.21813, 19.35227, 19.48641, 19.62053, 19.75465, 19.88875, 20.02285, 
    20.15693, 20.29099, 20.42505, 20.55909, 20.69311, 20.82712, 20.96111, 
    21.09508, 21.22903, 21.36296, 21.49687, 21.63076, 21.76463, 21.89848, 
    22.0323, 22.1661, 22.29987, 22.43362, 22.56734, 22.70103, 22.83469, 
    22.96832, 23.10193, 23.2355, 23.36904, 23.50255, 23.63602, 23.76947, 
    23.90287, 24.03624, 24.16958, 24.30287, 24.43613, 24.56935, 24.70253, 
    24.83567, 24.96877, 25.10183, 25.23484, 25.36782, 25.50074, 25.63362, 
    25.76646, 25.89925, 26.03199, 26.16469, 26.29733, 26.42993, 26.56248, 
    26.69497, 26.82742, 26.95981, 27.09214, 27.22443, 27.35666, 27.48883, 
    27.62095, 27.75301, 27.88501, 28.01696, 28.14885, 28.28067, 28.41244, 
    28.54414, 28.67579, 28.80737, 28.93888, 29.07034, 29.20173, 29.33305, 
    29.46431, 29.5955, 29.72662, 29.85767, 29.98866, 30.11958, 30.25042, 
    30.3812, 30.5119, 30.64253, 30.77309, 30.90358, 31.03399, 31.16433, 
    31.29459, 31.42478, 31.55488, 31.68492, 31.81487, 31.94474, 32.07454, 
    32.20425, 32.33389, 32.46344, 32.59292, 32.72231, 32.85162, 32.98084, 
    33.10998, 33.23903, 33.368, 33.49689, 33.62568, 33.75439, 33.88301, 
    34.01155, 34.13999, 34.26835, 34.39661, 34.52479, 34.65287, 34.78086, 
    34.90876, 35.03657, 35.16429, 35.29191, 35.41943, 35.54686, 35.6742, 
    35.80144, 35.92858, 36.05563, 36.18258, 36.30943, 36.43618, 36.56283, 
    36.68938, 36.81583, 36.94219, 37.06844, 37.19459, 37.32064, 37.44658, 
    37.57243, 37.69816, 37.8238, 37.94933, 38.07476, 38.20008, 38.32529, 
    38.4504, 38.5754, 38.7003, 38.82508, 38.94976, 39.07434, 39.1988, 
    39.32315, 39.4474, 39.57153, 39.69555, 39.81947, 39.94326, 40.06696, 
    40.19053, 40.314,
  -15.30197, -15.18998, -15.07785, -14.96559, -14.8532, -14.74067, -14.62801, 
    -14.51522, -14.4023, -14.28924, -14.17605, -14.06273, -13.94928, 
    -13.83569, -13.72197, -13.60812, -13.49414, -13.38003, -13.26579, 
    -13.15141, -13.0369, -12.92226, -12.80749, -12.69259, -12.57756, 
    -12.4624, -12.3471, -12.23168, -12.11612, -12.00044, -11.88462, 
    -11.76868, -11.6526, -11.5364, -11.42006, -11.3036, -11.18701, -11.07029, 
    -10.95344, -10.83646, -10.71935, -10.60211, -10.48475, -10.36726, 
    -10.24964, -10.13189, -10.01402, -9.896013, -9.777884, -9.659629, 
    -9.541247, -9.422738, -9.304104, -9.185344, -9.066458, -8.947446, 
    -8.82831, -8.709048, -8.589663, -8.470152, -8.350517, -8.230759, 
    -8.110876, -7.99087, -7.870742, -7.75049, -7.630116, -7.509619, 
    -7.389001, -7.26826, -7.147399, -7.026416, -6.905312, -6.784088, 
    -6.662744, -6.541279, -6.419695, -6.297992, -6.176169, -6.054228, 
    -5.932169, -5.809991, -5.687696, -5.565284, -5.442755, -5.320109, 
    -5.197347, -5.074468, -4.951475, -4.828366, -4.705142, -4.581803, 
    -4.458351, -4.334785, -4.211105, -4.087313, -3.963408, -3.839391, 
    -3.715262, -3.591022, -3.466671, -3.342209, -3.217637, -3.092956, 
    -2.968165, -2.843265, -2.718257, -2.593141, -2.467917, -2.342586, 
    -2.217148, -2.091604, -1.965955, -1.8402, -1.71434, -1.588376, -1.462308, 
    -1.336136, -1.209862, -1.083485, -0.9570059, -0.8304253, -0.7037437, 
    -0.5769616, -0.4500794, -0.3230977, -0.1960169, -0.06883766, 0.05843962, 
    0.1858144, 0.3132861, 0.4408543, 0.5685183, 0.6962778, 0.8241321, 
    0.9520807, 1.080123, 1.208259, 1.336487, 1.464807, 1.593219, 1.721722, 
    1.850315, 1.978998, 2.10777, 2.236631, 2.36558, 2.494617, 2.62374, 
    2.75295, 2.882246, 3.011627, 3.141092, 3.270641, 3.400274, 3.529989, 
    3.659787, 3.789665, 3.919625, 4.049665, 4.179785, 4.309983, 4.44026, 
    4.570615, 4.701046, 4.831554, 4.962138, 5.092797, 5.22353, 5.354338, 
    5.485218, 5.61617, 5.747195, 5.878291, 6.009457, 6.140692, 6.271997, 
    6.40337, 6.534811, 6.666319, 6.797894, 6.929533, 7.061238, 7.193007, 
    7.32484, 7.456736, 7.588693, 7.720712, 7.852792, 7.984931, 8.11713, 
    8.249388, 8.381703, 8.514075, 8.646504, 8.778988, 8.911528, 9.044121, 
    9.176767, 9.309466, 9.442218, 9.57502, 9.707872, 9.840775, 9.973726, 
    10.10673, 10.23977, 10.37287, 10.50601, 10.63919, 10.77242, 10.90569, 
    11.03901, 11.17236, 11.30576, 11.4392, 11.57268, 11.70619, 11.83975, 
    11.97334, 12.10697, 12.24064, 12.37434, 12.50807, 12.64184, 12.77564, 
    12.90947, 13.04333, 13.17722, 13.31115, 13.4451, 13.57908, 13.71308, 
    13.84711, 13.98117, 14.11525, 14.24936, 14.38349, 14.51764, 14.65181, 
    14.786, 14.92021, 15.05444, 15.18869, 15.32296, 15.45724, 15.59154, 
    15.72585, 15.86018, 15.99452, 16.12887, 16.26324, 16.39761, 16.53199, 
    16.66639, 16.80079, 16.9352, 17.06961, 17.20403, 17.33846, 17.47289, 
    17.60732, 17.74176, 17.8762, 18.01063, 18.14507, 18.27951, 18.41394, 
    18.54838, 18.68281, 18.81723, 18.95165, 19.08607, 19.22047, 19.35487, 
    19.48927, 19.62365, 19.75802, 19.89238, 20.02673, 20.16107, 20.29539, 
    20.42971, 20.564, 20.69828, 20.83254, 20.96679, 21.10102, 21.23523, 
    21.36942, 21.50359, 21.63773, 21.77186, 21.90596, 22.04004, 22.17409, 
    22.30812, 22.44212, 22.57609, 22.71004, 22.84396, 22.97785, 23.1117, 
    23.24553, 23.37932, 23.51309, 23.64682, 23.78051, 23.91417, 24.04779, 
    24.18138, 24.31493, 24.44844, 24.58191, 24.71534, 24.84874, 24.98209, 
    25.11539, 25.24866, 25.38188, 25.51506, 25.64819, 25.78128, 25.91432, 
    26.04731, 26.18025, 26.31315, 26.44599, 26.57878, 26.71153, 26.84422, 
    26.97686, 27.10944, 27.24197, 27.37445, 27.50687, 27.63923, 27.77154, 
    27.90379, 28.03597, 28.1681, 28.30017, 28.43218, 28.56413, 28.69602, 
    28.82784, 28.9596, 29.09129, 29.22292, 29.35449, 29.48598, 29.61741, 
    29.74878, 29.88007, 30.0113, 30.14245, 30.27354, 30.40455, 30.53549, 
    30.66636, 30.79716, 30.92788, 31.05852, 31.18909, 31.31959, 31.45001, 
    31.58035, 31.71062, 31.8408, 31.97091, 32.10094, 32.23088, 32.36075, 
    32.49054, 32.62024, 32.74986, 32.87939, 33.00885, 33.13821, 33.26749, 
    33.39669, 33.5258, 33.65482, 33.78376, 33.91261, 34.04136, 34.17003, 
    34.29861, 34.4271, 34.5555, 34.6838, 34.81202, 34.94014, 35.06816, 
    35.1961, 35.32394, 35.45168, 35.57933, 35.70689, 35.83434, 35.9617, 
    36.08896, 36.21613, 36.34319, 36.47016, 36.59702, 36.72379, 36.85046, 
    36.97702, 37.10348, 37.22984, 37.3561, 37.48226, 37.60831, 37.73426, 
    37.8601, 37.98584, 38.11147, 38.237, 38.36242, 38.48773, 38.61294, 
    38.73804, 38.86303, 38.98791, 39.11269, 39.23735, 39.3619, 39.48635, 
    39.61068, 39.73491, 39.85902, 39.98302, 40.1069, 40.23068, 40.35434,
  -15.35798, -15.24585, -15.13358, -15.02118, -14.90864, -14.79598, 
    -14.68318, -14.57024, -14.45717, -14.34397, -14.23064, -14.11717, 
    -14.00357, -13.88984, -13.77598, -13.66198, -13.54785, -13.43359, 
    -13.31919, -13.20467, -13.09001, -12.97522, -12.86029, -12.74524, 
    -12.63006, -12.51474, -12.39929, -12.28371, -12.168, -12.05216, 
    -11.93619, -11.82008, -11.70385, -11.58749, -11.47099, -11.35437, 
    -11.23762, -11.12073, -11.00372, -10.88658, -10.76931, -10.65191, 
    -10.53438, -10.41672, -10.29894, -10.18102, -10.06298, -9.94481, 
    -9.826513, -9.708089, -9.589537, -9.470859, -9.352053, -9.233121, 
    -9.114063, -8.99488, -8.875569, -8.756134, -8.636574, -8.516888, 
    -8.397078, -8.277143, -8.157083, -8.0369, -7.916593, -7.796162, 
    -7.675608, -7.554932, -7.434133, -7.313211, -7.192167, -7.071002, 
    -6.949715, -6.828306, -6.706778, -6.585128, -6.463358, -6.341468, 
    -6.219459, -6.09733, -5.975083, -5.852716, -5.730232, -5.60763, -5.48491, 
    -5.362072, -5.239118, -5.116047, -4.99286, -4.869558, -4.74614, 
    -4.622606, -4.498958, -4.375196, -4.25132, -4.12733, -4.003227, 
    -3.879011, -3.754683, -3.630243, -3.505692, -3.381029, -3.256255, 
    -3.131371, -3.006378, -2.881275, -2.756063, -2.630742, -2.505313, 
    -2.379776, -2.254133, -2.128382, -2.002525, -1.876562, -1.750493, 
    -1.62432, -1.498042, -1.37166, -1.245175, -1.118586, -0.9918953, 
    -0.8651021, -0.7382073, -0.6112115, -0.484115, -0.3569184, -0.2296223, 
    -0.102227, 0.02526676, 0.1528586, 0.2805479, 0.4083342, 0.536217, 
    0.6641957, 0.7922697, 0.9204386, 1.048702, 1.177059, 1.305509, 1.434052, 
    1.562686, 1.691412, 1.82023, 1.949137, 2.078135, 2.207221, 2.336396, 
    2.465659, 2.59501, 2.724447, 2.853971, 2.98358, 3.113275, 3.243053, 
    3.372916, 3.502861, 3.63289, 3.763, 3.893192, 4.023464, 4.153816, 
    4.284248, 4.414759, 4.545348, 4.676013, 4.806757, 4.937576, 5.068471, 
    5.19944, 5.330484, 5.461602, 5.592792, 5.724055, 5.855389, 5.986794, 
    6.118269, 6.249814, 6.381427, 6.513109, 6.644857, 6.776673, 6.908555, 
    7.040502, 7.172513, 7.304589, 7.436728, 7.568929, 7.701192, 7.833516, 
    7.9659, 8.098345, 8.230847, 8.363408, 8.496027, 8.628701, 8.761433, 
    8.894218, 9.02706, 9.159954, 9.292901, 9.4259, 9.558951, 9.692054, 
    9.825205, 9.958406, 10.09166, 10.22495, 10.3583, 10.49169, 10.62512, 
    10.7586, 10.89213, 11.02569, 11.1593, 11.29295, 11.42664, 11.56037, 
    11.69414, 11.82795, 11.9618, 12.09568, 12.2296, 12.36355, 12.49754, 
    12.63156, 12.76562, 12.89971, 13.03382, 13.16797, 13.30215, 13.43636, 
    13.57059, 13.70485, 13.83914, 13.97345, 14.10779, 14.24215, 14.37654, 
    14.51095, 14.64538, 14.77982, 14.91429, 15.04878, 15.18329, 15.31781, 
    15.45235, 15.58691, 15.72148, 15.85606, 15.99066, 16.12527, 16.25989, 
    16.39453, 16.52917, 16.66382, 16.79848, 16.93315, 17.06782, 17.2025, 
    17.33719, 17.47187, 17.60657, 17.74126, 17.87596, 18.01065, 18.14535, 
    18.28005, 18.41474, 18.54943, 18.68412, 18.8188, 18.95348, 19.08815, 
    19.22282, 19.35748, 19.49213, 19.62677, 19.7614, 19.89602, 20.03063, 
    20.16523, 20.29981, 20.43438, 20.56893, 20.70347, 20.83799, 20.97249, 
    21.10698, 21.24144, 21.37589, 21.51032, 21.64472, 21.7791, 21.91346, 
    22.04779, 22.1821, 22.31639, 22.45065, 22.58488, 22.71908, 22.85325, 
    22.98739, 23.12151, 23.25559, 23.38964, 23.52365, 23.65764, 23.79159, 
    23.9255, 24.05938, 24.19322, 24.32702, 24.46078, 24.59451, 24.72819, 
    24.86184, 24.99544, 25.129, 25.26252, 25.39599, 25.52942, 25.6628, 
    25.79614, 25.92943, 26.06267, 26.19586, 26.329, 26.4621, 26.59514, 
    26.72813, 26.86107, 26.99396, 27.12679, 27.25957, 27.39229, 27.52496, 
    27.65756, 27.79012, 27.92261, 28.05504, 28.18742, 28.31973, 28.45199, 
    28.58418, 28.71631, 28.84837, 28.98038, 29.11231, 29.24418, 29.37599, 
    29.50773, 29.6394, 29.771, 29.90253, 30.034, 30.16539, 30.29671, 
    30.42797, 30.55914, 30.69025, 30.82128, 30.95224, 31.08312, 31.21393, 
    31.34466, 31.47532, 31.60589, 31.73639, 31.86681, 31.99715, 32.12741, 
    32.25759, 32.38768, 32.5177, 32.64763, 32.77748, 32.90725, 33.03693, 
    33.16652, 33.29603, 33.42546, 33.55479, 33.68404, 33.81321, 33.94228, 
    34.07126, 34.20015, 34.32896, 34.45767, 34.58629, 34.71482, 34.84325, 
    34.97159, 35.09984, 35.228, 35.35606, 35.48402, 35.61189, 35.73966, 
    35.86733, 35.99491, 36.12239, 36.24976, 36.37704, 36.50423, 36.63131, 
    36.75829, 36.88517, 37.01194, 37.13862, 37.26519, 37.39166, 37.51802, 
    37.64429, 37.77044, 37.8965, 38.02244, 38.14828, 38.27401, 38.39964, 
    38.52516, 38.65057, 38.77588, 38.90107, 39.02616, 39.15113, 39.276, 
    39.40076, 39.5254, 39.64994, 39.77436, 39.89867, 40.02287, 40.14695, 
    40.27092, 40.39478,
  -15.41411, -15.30183, -15.18943, -15.07688, -14.96421, -14.8514, -14.73845, 
    -14.62538, -14.51217, -14.39882, -14.28534, -14.17173, -14.05799, 
    -13.94411, -13.83009, -13.71595, -13.60167, -13.48726, -13.37271, 
    -13.25804, -13.14323, -13.02829, -12.91321, -12.798, -12.68267, 
    -12.56719, -12.45159, -12.33586, -12.21999, -12.10399, -11.98786, 
    -11.8716, -11.75521, -11.63869, -11.52203, -11.40525, -11.28834, 
    -11.17129, -11.05412, -10.93681, -10.81938, -10.70181, -10.58412, 
    -10.4663, -10.34835, -10.23027, -10.11206, -9.99372, -9.875254, -9.75666, 
    -9.637939, -9.519091, -9.400114, -9.281011, -9.16178, -9.042423, 
    -8.92294, -8.80333, -8.683596, -8.563734, -8.443748, -8.323636, -8.2034, 
    -8.083038, -7.962553, -7.841943, -7.72121, -7.600353, -7.479373, 
    -7.358269, -7.237043, -7.115695, -6.994225, -6.872633, -6.750918, 
    -6.629084, -6.507128, -6.385051, -6.262855, -6.140538, -6.018102, 
    -5.895547, -5.772872, -5.65008, -5.527169, -5.40414, -5.280993, -5.15773, 
    -5.03435, -4.910853, -4.78724, -4.663512, -4.539668, -4.415709, 
    -4.291636, -4.167448, -4.043147, -3.918732, -3.794204, -3.669564, 
    -3.544812, -3.419948, -3.294973, -3.169886, -3.044689, -2.919383, 
    -2.793966, -2.66844, -2.542806, -2.417063, -2.291213, -2.165255, 
    -2.03919, -1.913018, -1.786741, -1.660358, -1.53387, -1.407277, 
    -1.280581, -1.15378, -1.026877, -0.8998705, -0.7727621, -0.645552, 
    -0.5182408, -0.3908289, -0.2633169, -0.1357053, -0.007994519, 0.1198148, 
    0.2477222, 0.3757271, 0.5038291, 0.6320274, 0.7603217, 0.8887114, 
    1.017196, 1.145775, 1.274447, 1.403213, 1.532071, 1.661021, 1.790063, 
    1.919195, 2.048418, 2.177731, 2.307132, 2.436622, 2.5662, 2.695866, 
    2.825618, 2.955456, 3.08538, 3.215389, 3.345482, 3.475659, 3.605919, 
    3.736261, 3.866685, 3.99719, 4.127776, 4.258441, 4.389186, 4.52001, 
    4.650911, 4.78189, 4.912945, 5.044076, 5.175283, 5.306565, 5.43792, 
    5.569348, 5.70085, 5.832423, 5.964067, 6.095783, 6.227568, 6.359422, 
    6.491344, 6.623335, 6.755393, 6.887516, 7.019707, 7.151961, 7.28428, 
    7.416663, 7.549109, 7.681616, 7.814185, 7.946815, 8.079505, 8.212254, 
    8.345061, 8.477926, 8.610848, 8.743827, 8.876861, 9.00995, 9.143092, 
    9.276288, 9.409537, 9.542837, 9.676188, 9.80959, 9.943042, 10.07654, 
    10.21009, 10.34368, 10.47733, 10.61101, 10.74474, 10.87852, 11.01234, 
    11.1462, 11.28011, 11.41405, 11.54803, 11.68206, 11.81612, 11.95022, 
    12.08436, 12.21853, 12.35274, 12.48698, 12.62126, 12.75557, 12.88991, 
    13.02429, 13.15869, 13.29313, 13.42759, 13.56208, 13.6966, 13.83114, 
    13.96571, 14.10031, 14.23493, 14.36957, 14.50424, 14.63892, 14.77363, 
    14.90836, 15.0431, 15.17787, 15.31265, 15.44745, 15.58226, 15.71709, 
    15.85194, 15.98679, 16.12166, 16.25654, 16.39144, 16.52634, 16.66125, 
    16.79617, 16.93109, 17.06603, 17.20097, 17.33591, 17.47086, 17.60581, 
    17.74076, 17.87572, 18.01067, 18.14563, 18.28058, 18.41554, 18.55049, 
    18.68544, 18.82038, 18.95532, 19.09025, 19.22518, 19.36009, 19.495, 
    19.6299, 19.76479, 19.89967, 20.03454, 20.16939, 20.30424, 20.43906, 
    20.57388, 20.70867, 20.84345, 20.97821, 21.11296, 21.24768, 21.38238, 
    21.51707, 21.65173, 21.78637, 21.92098, 22.05557, 22.19014, 22.32468, 
    22.4592, 22.59368, 22.72814, 22.86257, 22.99697, 23.13134, 23.26568, 
    23.39998, 23.53425, 23.66849, 23.80269, 23.93686, 24.07099, 24.20509, 
    24.33915, 24.47316, 24.60714, 24.74108, 24.87498, 25.00883, 25.14264, 
    25.27641, 25.41014, 25.54382, 25.67745, 25.81104, 25.94458, 26.07807, 
    26.21152, 26.34491, 26.47825, 26.61154, 26.74479, 26.87797, 27.01111, 
    27.14419, 27.27721, 27.41018, 27.54309, 27.67595, 27.80875, 27.94149, 
    28.07417, 28.20679, 28.33935, 28.47185, 28.60428, 28.73665, 28.86896, 
    29.00121, 29.13339, 29.2655, 29.39755, 29.52953, 29.66144, 29.79328, 
    29.92506, 30.05676, 30.18839, 30.31996, 30.45145, 30.58286, 30.71421, 
    30.84548, 30.97667, 31.10779, 31.23883, 31.3698, 31.50069, 31.6315, 
    31.76223, 31.89289, 32.02346, 32.15395, 32.28436, 32.41469, 32.54494, 
    32.6751, 32.80518, 32.93518, 33.06509, 33.19491, 33.32465, 33.4543, 
    33.58387, 33.71334, 33.84273, 33.97203, 34.10124, 34.23035, 34.35938, 
    34.48832, 34.61716, 34.74591, 34.87457, 35.00314, 35.1316, 35.25998, 
    35.38826, 35.51644, 35.64453, 35.77252, 35.90041, 36.0282, 36.1559, 
    36.28349, 36.41099, 36.53839, 36.66568, 36.79288, 36.91997, 37.04696, 
    37.17384, 37.30063, 37.42731, 37.55389, 37.68036, 37.80672, 37.93298, 
    38.05914, 38.18519, 38.31113, 38.43696, 38.56269, 38.6883, 38.81381, 
    38.93921, 39.0645, 39.18968, 39.31475, 39.43971, 39.56455, 39.68929, 
    39.81391, 39.93842, 40.06282, 40.1871, 40.31127, 40.43533,
  -15.47035, -15.35794, -15.24539, -15.13271, -15.01989, -14.90694, 
    -14.79385, -14.68063, -14.56728, -14.45378, -14.34016, -14.2264, 
    -14.11251, -13.99849, -13.88433, -13.77003, -13.65561, -13.54105, 
    -13.42635, -13.31153, -13.19656, -13.08147, -12.96624, -12.85088, 
    -12.73539, -12.61977, -12.50401, -12.38812, -12.2721, -12.15594, 
    -12.03965, -11.92324, -11.80669, -11.69, -11.57319, -11.45625, -11.33917, 
    -11.22196, -11.10463, -10.98716, -10.86956, -10.75183, -10.63398, 
    -10.51599, -10.39787, -10.27962, -10.16125, -10.04274, -9.924108, 
    -9.805346, -9.686454, -9.567434, -9.448287, -9.329012, -9.209609, 
    -9.090079, -8.970423, -8.850639, -8.730729, -8.610692, -8.49053, 
    -8.370241, -8.249827, -8.129288, -8.008624, -7.887835, -7.766922, 
    -7.645884, -7.524722, -7.403437, -7.282029, -7.160497, -7.038843, 
    -6.917066, -6.795167, -6.673147, -6.551005, -6.428741, -6.306357, 
    -6.183853, -6.061228, -5.938483, -5.815619, -5.692636, -5.569533, 
    -5.446313, -5.322974, -5.199517, -5.075943, -4.952252, -4.828444, 
    -4.70452, -4.58048, -4.456325, -4.332054, -4.207668, -4.083168, 
    -3.958554, -3.833827, -3.708986, -3.584033, -3.458967, -3.333789, 
    -3.2085, -3.0831, -2.957589, -2.831968, -2.706237, -2.580396, -2.454447, 
    -2.328389, -2.202224, -2.075951, -1.949571, -1.823084, -1.696491, 
    -1.569792, -1.442988, -1.31608, -1.189067, -1.061951, -0.9347309, 
    -0.8074085, -0.6799838, -0.5524574, -0.4248298, -0.2971015, -0.169273, 
    -0.04134479, 0.08668252, 0.2148084, 0.3430324, 0.471354, 0.5997726, 
    0.7282876, 0.8568985, 0.9856048, 1.114406, 1.243301, 1.37229, 1.501372, 
    1.630547, 1.759814, 1.889172, 2.01862, 2.14816, 2.277788, 2.407506, 
    2.537312, 2.667206, 2.797188, 2.927255, 3.057409, 3.187649, 3.317973, 
    3.448381, 3.578873, 3.709447, 3.840105, 3.970843, 4.101663, 4.232563, 
    4.363543, 4.494601, 4.625739, 4.756953, 4.888246, 5.019614, 5.151058, 
    5.282578, 5.414171, 5.545839, 5.677579, 5.809392, 5.941277, 6.073233, 
    6.205258, 6.337354, 6.469519, 6.601751, 6.734052, 6.866419, 6.998852, 
    7.131351, 7.263914, 7.396541, 7.529232, 7.661984, 7.794799, 7.927675, 
    8.060611, 8.193606, 8.326661, 8.459774, 8.592944, 8.726171, 8.859453, 
    8.99279, 9.126183, 9.259628, 9.393126, 9.526677, 9.660278, 9.793931, 
    9.927633, 10.06138, 10.19518, 10.32903, 10.46292, 10.59686, 10.73085, 
    10.86488, 10.99895, 11.13306, 11.26722, 11.40142, 11.53566, 11.66994, 
    11.80425, 11.93861, 12.073, 12.20743, 12.3419, 12.4764, 12.61093, 
    12.74549, 12.88009, 13.01472, 13.14939, 13.28408, 13.4188, 13.55354, 
    13.68832, 13.82312, 13.95795, 14.0928, 14.22768, 14.36258, 14.49751, 
    14.63245, 14.76742, 14.9024, 15.03741, 15.17243, 15.30747, 15.44253, 
    15.57761, 15.71269, 15.8478, 15.98291, 16.11804, 16.25318, 16.38833, 
    16.5235, 16.65867, 16.79385, 16.92903, 17.06423, 17.19942, 17.33463, 
    17.46984, 17.60505, 17.74026, 17.87548, 18.01069, 18.14591, 18.28113, 
    18.41634, 18.55155, 18.68676, 18.82196, 18.95716, 19.09235, 19.22754, 
    19.36271, 19.49788, 19.63305, 19.76819, 19.90333, 20.03846, 20.17357, 
    20.30868, 20.44376, 20.57883, 20.71389, 20.84893, 20.98395, 21.11895, 
    21.25393, 21.3889, 21.52384, 21.65876, 21.79366, 21.92853, 22.06338, 
    22.1982, 22.333, 22.46777, 22.60252, 22.73723, 22.87192, 23.00657, 
    23.1412, 23.27579, 23.41035, 23.54488, 23.67938, 23.81384, 23.94826, 
    24.08265, 24.217, 24.35131, 24.48558, 24.61981, 24.754, 24.88815, 
    25.02226, 25.15633, 25.29035, 25.42433, 25.55826, 25.69214, 25.82598, 
    25.95978, 26.09352, 26.22721, 26.36086, 26.49445, 26.62799, 26.76148, 
    26.89492, 27.02831, 27.16163, 27.29491, 27.42813, 27.56129, 27.69439, 
    27.82743, 27.96042, 28.09335, 28.22621, 28.35902, 28.49176, 28.62444, 
    28.75706, 28.88961, 29.0221, 29.15452, 29.28688, 29.41917, 29.55139, 
    29.68355, 29.81563, 29.94765, 30.07959, 30.21146, 30.34327, 30.47499, 
    30.60665, 30.73823, 30.86974, 31.00117, 31.13253, 31.26381, 31.39501, 
    31.52614, 31.65718, 31.78815, 31.91904, 32.04984, 32.18057, 32.31121, 
    32.44178, 32.57225, 32.70265, 32.83296, 32.96318, 33.09333, 33.22338, 
    33.35335, 33.48323, 33.61302, 33.74272, 33.87234, 34.00186, 34.1313, 
    34.26064, 34.38989, 34.51905, 34.64812, 34.7771, 34.90598, 35.03476, 
    35.16345, 35.29205, 35.42055, 35.54895, 35.67726, 35.80547, 35.93357, 
    36.06159, 36.1895, 36.31731, 36.44503, 36.57264, 36.70015, 36.82756, 
    36.95486, 37.08207, 37.20916, 37.33616, 37.46305, 37.58984, 37.71652, 
    37.8431, 37.96957, 38.09593, 38.22219, 38.34834, 38.47438, 38.60031, 
    38.72613, 38.85184, 38.97745, 39.10294, 39.22832, 39.3536, 39.47876, 
    39.60381, 39.72874, 39.85357, 39.97828, 40.10287, 40.22735, 40.35172, 
    40.47597,
  -15.52671, -15.41416, -15.30147, -15.18864, -15.07569, -14.96259, 
    -14.84936, -14.736, -14.6225, -14.50887, -14.3951, -14.28119, -14.16716, 
    -14.05298, -13.93868, -13.82424, -13.70966, -13.59495, -13.48011, 
    -13.36513, -13.25002, -13.13477, -13.01939, -12.90388, -12.78823, 
    -12.67245, -12.55654, -12.4405, -12.32432, -12.20801, -12.09156, 
    -11.97499, -11.85828, -11.74144, -11.62446, -11.50736, -11.39012, 
    -11.27275, -11.15525, -11.03762, -10.91986, -10.80197, -10.68395, 
    -10.56579, -10.44751, -10.3291, -10.21055, -10.09188, -9.973076, 
    -9.854143, -9.735082, -9.615892, -9.496573, -9.377127, -9.257551, 
    -9.137848, -9.018018, -8.89806, -8.777974, -8.657762, -8.537423, 
    -8.416958, -8.296366, -8.175649, -8.054806, -7.933837, -7.812743, 
    -7.691525, -7.570182, -7.448715, -7.327124, -7.205409, -7.08357, 
    -6.961609, -6.839525, -6.717319, -6.59499, -6.47254, -6.349968, 
    -6.227275, -6.104461, -5.981527, -5.858472, -5.735298, -5.612004, 
    -5.488591, -5.365059, -5.241409, -5.117641, -4.993755, -4.869752, 
    -4.745632, -4.621396, -4.497043, -4.372574, -4.247991, -4.123292, 
    -3.998478, -3.873551, -3.748509, -3.623354, -3.498086, -3.372706, 
    -3.247214, -3.121609, -2.995894, -2.870068, -2.744131, -2.618085, 
    -2.491929, -2.365664, -2.23929, -2.112808, -1.986219, -1.859522, 
    -1.732718, -1.605809, -1.478794, -1.351673, -1.224447, -1.097118, 
    -0.9696839, -0.8421471, -0.7145073, -0.5867653, -0.4589216, -0.3309765, 
    -0.2029307, -0.07478464, 0.0534611, 0.181806, 0.3102496, 0.4387912, 
    0.5674304, 0.6961666, 0.8249993, 0.9539279, 1.082952, 1.21207, 1.341283, 
    1.47059, 1.59999, 1.729482, 1.859066, 1.988741, 2.118507, 2.248363, 
    2.378309, 2.508344, 2.638467, 2.768678, 2.898976, 3.029361, 3.159831, 
    3.290387, 3.421027, 3.551752, 3.682559, 3.81345, 3.944422, 4.075477, 
    4.206612, 4.337827, 4.469121, 4.600495, 4.731947, 4.863476, 4.995082, 
    5.126765, 5.258523, 5.390356, 5.522263, 5.654243, 5.786296, 5.918422, 
    6.050619, 6.182886, 6.315224, 6.447631, 6.580106, 6.71265, 6.845261, 
    6.977938, 7.110681, 7.243489, 7.376361, 7.509297, 7.642296, 7.775357, 
    7.90848, 8.041663, 8.174906, 8.308208, 8.441569, 8.574987, 8.708463, 
    8.841994, 8.975581, 9.109223, 9.242919, 9.376668, 9.510469, 9.644321, 
    9.778226, 9.912179, 10.04618, 10.18023, 10.31433, 10.44848, 10.58267, 
    10.71691, 10.85119, 10.98552, 11.11989, 11.2543, 11.38875, 11.52325, 
    11.65778, 11.79235, 11.92696, 12.06161, 12.1963, 12.33102, 12.46578, 
    12.60056, 12.73539, 12.87024, 13.00513, 13.14005, 13.275, 13.40998, 
    13.54498, 13.68002, 13.81508, 13.95017, 14.08528, 14.22042, 14.35557, 
    14.49076, 14.62596, 14.76119, 14.89643, 15.0317, 15.16698, 15.30228, 
    15.4376, 15.57293, 15.70828, 15.84365, 15.97902, 16.11441, 16.24981, 
    16.38523, 16.52065, 16.65608, 16.79152, 16.92697, 17.06242, 17.19788, 
    17.33335, 17.46881, 17.60429, 17.73976, 17.87524, 18.01072, 18.14619, 
    18.28167, 18.41714, 18.55262, 18.68808, 18.82355, 18.95901, 19.09446, 
    19.22991, 19.36535, 19.50077, 19.6362, 19.77161, 19.90701, 20.04239, 
    20.17777, 20.31313, 20.44847, 20.58381, 20.71912, 20.85442, 20.9897, 
    21.12496, 21.2602, 21.39543, 21.53063, 21.66581, 21.80096, 21.9361, 
    22.0712, 22.20629, 22.34134, 22.47637, 22.61138, 22.74635, 22.88129, 
    23.01621, 23.15109, 23.28594, 23.42076, 23.55554, 23.69029, 23.82501, 
    23.95969, 24.09433, 24.22894, 24.3635, 24.49803, 24.63252, 24.76696, 
    24.90137, 25.03573, 25.17005, 25.30433, 25.43856, 25.57274, 25.70688, 
    25.84097, 25.97502, 26.10901, 26.24296, 26.37686, 26.5107, 26.64449, 
    26.77823, 26.91192, 27.04555, 27.17913, 27.31265, 27.44612, 27.57953, 
    27.71288, 27.84617, 27.97941, 28.11258, 28.2457, 28.37875, 28.51174, 
    28.64466, 28.77752, 28.91032, 29.04305, 29.17572, 29.30832, 29.44085, 
    29.57332, 29.70572, 29.83804, 29.9703, 30.10248, 30.2346, 30.36664, 
    30.49861, 30.6305, 30.76233, 30.89407, 31.02574, 31.15734, 31.28885, 
    31.42029, 31.55165, 31.68293, 31.81414, 31.94526, 32.0763, 32.20726, 
    32.33814, 32.46893, 32.59964, 32.73027, 32.86081, 32.99127, 33.12164, 
    33.25193, 33.38212, 33.51223, 33.64225, 33.77218, 33.90203, 34.03178, 
    34.16144, 34.29101, 34.42049, 34.54987, 34.67916, 34.80836, 34.93747, 
    35.06647, 35.19538, 35.3242, 35.45293, 35.58155, 35.71008, 35.8385, 
    35.96683, 36.09506, 36.22319, 36.35122, 36.47915, 36.60698, 36.7347, 
    36.86233, 36.98985, 37.11727, 37.24458, 37.37179, 37.49889, 37.62589, 
    37.75278, 37.87957, 38.00625, 38.13282, 38.25929, 38.38564, 38.51189, 
    38.63803, 38.76406, 38.88998, 39.01579, 39.14149, 39.26707, 39.39255, 
    39.51791, 39.64316, 39.7683, 39.89332, 40.01823, 40.14302, 40.2677, 
    40.39227, 40.51672,
  -15.58318, -15.47049, -15.35766, -15.2447, -15.1316, -15.01836, -14.90499, 
    -14.79149, -14.67784, -14.56406, -14.45015, -14.3361, -14.22192, 
    -14.1076, -13.99314, -13.87856, -13.76383, -13.64897, -13.53398, 
    -13.41885, -13.30359, -13.18819, -13.07266, -12.95699, -12.84119, 
    -12.72526, -12.60919, -12.49299, -12.37666, -12.26019, -12.14359, 
    -12.02685, -11.90998, -11.79298, -11.67585, -11.55859, -11.44119, 
    -11.32366, -11.206, -11.0882, -10.97028, -10.85222, -10.73403, -10.61571, 
    -10.49726, -10.37868, -10.25997, -10.14113, -10.02216, -9.903056, 
    -9.783824, -9.664464, -9.544973, -9.425355, -9.305607, -9.18573, 
    -9.065725, -8.945593, -8.825333, -8.704944, -8.584429, -8.463786, 
    -8.343017, -8.22212, -8.101098, -7.97995, -7.858676, -7.737277, 
    -7.615752, -7.494102, -7.372328, -7.25043, -7.128407, -7.006261, 
    -6.883992, -6.7616, -6.639084, -6.516447, -6.393686, -6.270805, 
    -6.147802, -6.024677, -5.901433, -5.778067, -5.654581, -5.530976, 
    -5.407251, -5.283407, -5.159445, -5.035364, -4.911165, -4.786849, 
    -4.662416, -4.537866, -4.413199, -4.288416, -4.163518, -4.038505, 
    -3.913377, -3.788134, -3.662777, -3.537307, -3.411724, -3.286028, 
    -3.160219, -3.034299, -2.908267, -2.782125, -2.655872, -2.529508, 
    -2.403035, -2.276453, -2.149762, -2.022963, -1.896056, -1.769042, 
    -1.641921, -1.514694, -1.38736, -1.259922, -1.132378, -1.00473, 
    -0.8769786, -0.7491233, -0.6211653, -0.4931049, -0.3649426, -0.236679, 
    -0.1083147, 0.02014998, 0.1487144, 0.2773779, 0.4061401, 0.5350005, 
    0.6639584, 0.7930133, 0.9221646, 1.051412, 1.180754, 1.310192, 1.439723, 
    1.569348, 1.699066, 1.828877, 1.958779, 2.088773, 2.218858, 2.349032, 
    2.479296, 2.609649, 2.74009, 2.870618, 3.001234, 3.131936, 3.262724, 
    3.393597, 3.524554, 3.655596, 3.786721, 3.917928, 4.049217, 4.180588, 
    4.312039, 4.44357, 4.575181, 4.70687, 4.838637, 4.970481, 5.102402, 
    5.2344, 5.366472, 5.498619, 5.63084, 5.763134, 5.895501, 6.02794, 
    6.16045, 6.29303, 6.42568, 6.558399, 6.691186, 6.824042, 6.956964, 
    7.089952, 7.223005, 7.356123, 7.489305, 7.622551, 7.755859, 7.889229, 
    8.02266, 8.156151, 8.289701, 8.423311, 8.556979, 8.690704, 8.824486, 
    8.958323, 9.092215, 9.226161, 9.360162, 9.494214, 9.628319, 9.762475, 
    9.896681, 10.03094, 10.16524, 10.29959, 10.43399, 10.56844, 10.70293, 
    10.83747, 10.97205, 11.10668, 11.24134, 11.37605, 11.5108, 11.64559, 
    11.78042, 11.91529, 12.05019, 12.18513, 12.32011, 12.45512, 12.59017, 
    12.72525, 12.86037, 12.99551, 13.13069, 13.2659, 13.40113, 13.5364, 
    13.67169, 13.80701, 13.94236, 14.07773, 14.21313, 14.34855, 14.48399, 
    14.61945, 14.75494, 14.89044, 15.02597, 15.16151, 15.29707, 15.43265, 
    15.56825, 15.70386, 15.83948, 15.97512, 16.11077, 16.24643, 16.38211, 
    16.51779, 16.65348, 16.78918, 16.92489, 17.06061, 17.19633, 17.33206, 
    17.46779, 17.60352, 17.73926, 17.875, 18.01074, 18.14647, 18.28221, 
    18.41795, 18.55368, 18.68941, 18.82514, 18.96086, 19.09657, 19.23228, 
    19.36798, 19.50367, 19.63935, 19.77503, 19.91069, 20.04634, 20.18197, 
    20.31759, 20.4532, 20.58879, 20.72437, 20.85993, 20.99547, 21.13099, 
    21.26649, 21.40198, 21.53744, 21.67288, 21.80829, 21.94369, 22.07905, 
    22.2144, 22.34971, 22.485, 22.62026, 22.75549, 22.8907, 23.02587, 
    23.16101, 23.29612, 23.43119, 23.56623, 23.70124, 23.83622, 23.97115, 
    24.10605, 24.24091, 24.37573, 24.51052, 24.64526, 24.77996, 24.91462, 
    25.04924, 25.18382, 25.31834, 25.45283, 25.58727, 25.72166, 25.85601, 
    25.9903, 26.12455, 26.25875, 26.3929, 26.52699, 26.66104, 26.79503, 
    26.92897, 27.06285, 27.19668, 27.33045, 27.46417, 27.59783, 27.73143, 
    27.86497, 27.99845, 28.13187, 28.26523, 28.39853, 28.53176, 28.66494, 
    28.79805, 28.93109, 29.06407, 29.19698, 29.32982, 29.4626, 29.59531, 
    29.72795, 29.86052, 29.99302, 30.12544, 30.2578, 30.39008, 30.52229, 
    30.65442, 30.78649, 30.91847, 31.05038, 31.18221, 31.31397, 31.44564, 
    31.57724, 31.70876, 31.8402, 31.97156, 32.10283, 32.23403, 32.36514, 
    32.49617, 32.62711, 32.75797, 32.88874, 33.01943, 33.15004, 33.28055, 
    33.41098, 33.54132, 33.67157, 33.80173, 33.9318, 34.06178, 34.19166, 
    34.32146, 34.45116, 34.58077, 34.71029, 34.83971, 34.96904, 35.09827, 
    35.22741, 35.35645, 35.48539, 35.61423, 35.74298, 35.87163, 36.00018, 
    36.12863, 36.25697, 36.38522, 36.51337, 36.64141, 36.76936, 36.89719, 
    37.02493, 37.15256, 37.28009, 37.40751, 37.53482, 37.66204, 37.78914, 
    37.91614, 38.04303, 38.16981, 38.29648, 38.42305, 38.5495, 38.67585, 
    38.80209, 38.92821, 39.05423, 39.18013, 39.30592, 39.43159, 39.55716, 
    39.68261, 39.80795, 39.93318, 40.05829, 40.18328, 40.30816, 40.43293, 
    40.55758,
  -15.63978, -15.52695, -15.41398, -15.30087, -15.18763, -15.07425, 
    -14.96074, -14.84709, -14.7333, -14.61938, -14.50532, -14.39113, 
    -14.2768, -14.16233, -14.04773, -13.93299, -13.81812, -13.70311, 
    -13.58797, -13.47269, -13.35728, -13.24173, -13.12604, -13.01022, 
    -12.89427, -12.77818, -12.66196, -12.5456, -12.42911, -12.31249, 
    -12.19573, -12.07883, -11.96181, -11.84465, -11.72736, -11.60993, 
    -11.49237, -11.37468, -11.25686, -11.1389, -11.02081, -10.90259, 
    -10.78423, -10.66575, -10.54713, -10.42838, -10.30951, -10.1905, 
    -10.07135, -9.952083, -9.832682, -9.71315, -9.593488, -9.473697, 
    -9.353776, -9.233727, -9.113547, -8.993239, -8.872804, -8.752239, 
    -8.631547, -8.510727, -8.38978, -8.268705, -8.147504, -8.026175, 
    -7.904721, -7.78314, -7.661434, -7.539602, -7.417645, -7.295562, 
    -7.173355, -7.051024, -6.928569, -6.80599, -6.683288, -6.560462, 
    -6.437514, -6.314444, -6.191251, -6.067936, -5.9445, -5.820943, 
    -5.697266, -5.573468, -5.44955, -5.325511, -5.201355, -5.077078, 
    -4.952684, -4.828171, -4.703541, -4.578793, -4.453928, -4.328946, 
    -4.203848, -4.078635, -3.953305, -3.827861, -3.702302, -3.57663, 
    -3.450843, -3.324943, -3.19893, -3.072804, -2.946567, -2.820218, 
    -2.693758, -2.567187, -2.440506, -2.313715, -2.186814, -2.059805, 
    -1.932688, -1.805462, -1.678129, -1.55069, -1.423143, -1.295491, 
    -1.167733, -1.039871, -0.9119035, -0.7838324, -0.6556578, -0.5273803, 
    -0.3990004, -0.2705186, -0.1419354, -0.01325142, 0.1155329, 0.2444169, 
    0.3734002, 0.5024821, 0.6316622, 0.7609398, 0.8903144, 1.019786, 
    1.149352, 1.279015, 1.408772, 1.538623, 1.668567, 1.798605, 1.928735, 
    2.058957, 2.18927, 2.319673, 2.450167, 2.58075, 2.711421, 2.842181, 
    2.973029, 3.103963, 3.234984, 3.36609, 3.497281, 3.628557, 3.759916, 
    3.891359, 4.022883, 4.15449, 4.286178, 4.417946, 4.549794, 4.681721, 
    4.813727, 4.94581, 5.077971, 5.210208, 5.342521, 5.474908, 5.607371, 
    5.739906, 5.872515, 6.005197, 6.137949, 6.270773, 6.403666, 6.53663, 
    6.669662, 6.802762, 6.935929, 7.069163, 7.202463, 7.335827, 7.469256, 
    7.602749, 7.736305, 7.869923, 8.003602, 8.137342, 8.271142, 8.405001, 
    8.538918, 8.672894, 8.806926, 8.941013, 9.075157, 9.209355, 9.343607, 
    9.477912, 9.612268, 9.746677, 9.881137, 10.01565, 10.1502, 10.28481, 
    10.41947, 10.55417, 10.68891, 10.82371, 10.95854, 11.09342, 11.22834, 
    11.36331, 11.49832, 11.63336, 11.76845, 11.90357, 12.03873, 12.17393, 
    12.30917, 12.44444, 12.57975, 12.71509, 12.85046, 12.98586, 13.1213, 
    13.25677, 13.39226, 13.52779, 13.66334, 13.79892, 13.93453, 14.07016, 
    14.20581, 14.34149, 14.4772, 14.61292, 14.74867, 14.88444, 15.02022, 
    15.15603, 15.29185, 15.42769, 15.56355, 15.69942, 15.83531, 15.97121, 
    16.10712, 16.24304, 16.37898, 16.51493, 16.65088, 16.78684, 16.92281, 
    17.05879, 17.19478, 17.33076, 17.46676, 17.60275, 17.73875, 17.87476, 
    18.01076, 18.14676, 18.28276, 18.41876, 18.55475, 18.69075, 18.82673, 
    18.96272, 19.09869, 19.23466, 19.37063, 19.50658, 19.64252, 19.77846, 
    19.91438, 20.05029, 20.18619, 20.32207, 20.45794, 20.5938, 20.72964, 
    20.86546, 21.00126, 21.13704, 21.2728, 21.40855, 21.54427, 21.67997, 
    21.81565, 21.9513, 22.08693, 22.22253, 22.3581, 22.49365, 22.62917, 
    22.76467, 22.90013, 23.03556, 23.17096, 23.30632, 23.44166, 23.57696, 
    23.71222, 23.84745, 23.98265, 24.11781, 24.25292, 24.388, 24.52304, 
    24.65804, 24.793, 24.92792, 25.06279, 25.19762, 25.33241, 25.46714, 
    25.60184, 25.73648, 25.87108, 26.00563, 26.14014, 26.27459, 26.40899, 
    26.54334, 26.67763, 26.81188, 26.94607, 27.0802, 27.21428, 27.3483, 
    27.48227, 27.61618, 27.75003, 27.88382, 28.01755, 28.15122, 28.28483, 
    28.41837, 28.55186, 28.68527, 28.81863, 28.95192, 29.08514, 29.2183, 
    29.35139, 29.48441, 29.61736, 29.75024, 29.88305, 30.0158, 30.14847, 
    30.28106, 30.41359, 30.54604, 30.67841, 30.81071, 30.94294, 31.07509, 
    31.20716, 31.33915, 31.47107, 31.6029, 31.73466, 31.86633, 31.99793, 
    32.12944, 32.26087, 32.39222, 32.52348, 32.65466, 32.78575, 32.91676, 
    33.04768, 33.17851, 33.30925, 33.43991, 33.57048, 33.70096, 33.83135, 
    33.96165, 34.09185, 34.22197, 34.35199, 34.48192, 34.61176, 34.7415, 
    34.87115, 35.0007, 35.13016, 35.25952, 35.38878, 35.51794, 35.64701, 
    35.77598, 35.90485, 36.03362, 36.16228, 36.29085, 36.41932, 36.54768, 
    36.67594, 36.8041, 36.93215, 37.0601, 37.18795, 37.31569, 37.44333, 
    37.57085, 37.69828, 37.8256, 37.9528, 38.0799, 38.20689, 38.33378, 
    38.46055, 38.58722, 38.71377, 38.84021, 38.96654, 39.09276, 39.21887, 
    39.34486, 39.47075, 39.59652, 39.72217, 39.84771, 39.97314, 40.09845, 
    40.22364, 40.34872, 40.47369, 40.59853,
  -15.69649, -15.58352, -15.47041, -15.35717, -15.24378, -15.13026, 
    -15.01661, -14.90281, -14.78888, -14.67482, -14.56061, -14.44627, 
    -14.3318, -14.21719, -14.10244, -13.98755, -13.87253, -13.75737, 
    -13.64208, -13.52665, -13.41108, -13.29538, -13.17954, -13.06357, 
    -12.94746, -12.83122, -12.71484, -12.59833, -12.48168, -12.3649, 
    -12.24799, -12.13094, -12.01375, -11.89643, -11.77898, -11.66139, 
    -11.54367, -11.42582, -11.30783, -11.18971, -11.07146, -10.95307, 
    -10.83455, -10.7159, -10.59712, -10.4782, -10.35916, -10.23998, 
    -10.12067, -10.00123, -9.881654, -9.761951, -9.642118, -9.522154, 
    -9.402061, -9.281837, -9.161484, -9.041001, -8.920389, -8.799649, 
    -8.67878, -8.557782, -8.436656, -8.315403, -8.194022, -8.072514, 
    -7.950878, -7.829116, -7.707227, -7.585213, -7.463072, -7.340806, 
    -7.218414, -7.095898, -6.973257, -6.850491, -6.727601, -6.604588, 
    -6.481451, -6.358191, -6.234809, -6.111304, -5.987677, -5.863928, 
    -5.740058, -5.616067, -5.491955, -5.367723, -5.243371, -5.118899, 
    -4.994308, -4.869599, -4.744771, -4.619825, -4.494761, -4.36958, 
    -4.244282, -4.118868, -3.993338, -3.867692, -3.74193, -3.616055, 
    -3.490064, -3.36396, -3.237742, -3.111411, -2.984967, -2.858411, 
    -2.731744, -2.604965, -2.478075, -2.351075, -2.223964, -2.096745, 
    -1.969416, -1.841979, -1.714434, -1.586782, -1.459022, -1.331156, 
    -1.203183, -1.075105, -0.9469225, -0.818635, -0.6902435, -0.5617485, 
    -0.4331505, -0.30445, -0.1756475, -0.04674372, 0.08226098, 0.211366, 
    0.3405708, 0.4698748, 0.5992776, 0.7287784, 0.8583767, 0.9880721, 
    1.117864, 1.247751, 1.377734, 1.507812, 1.637984, 1.768249, 1.898607, 
    2.029058, 2.1596, 2.290233, 2.420957, 2.55177, 2.682673, 2.813665, 
    2.944745, 3.075912, 3.207165, 3.338506, 3.469931, 3.601441, 3.733036, 
    3.864714, 3.996475, 4.128319, 4.260244, 4.39225, 4.524336, 4.656502, 
    4.788746, 4.921069, 5.05347, 5.185947, 5.318501, 5.45113, 5.583834, 
    5.716612, 5.849463, 5.982388, 6.115384, 6.248452, 6.381589, 6.514798, 
    6.648075, 6.78142, 6.914834, 7.048314, 7.18186, 7.315472, 7.449149, 
    7.58289, 7.716694, 7.85056, 7.984489, 8.118478, 8.252528, 8.386637, 
    8.520805, 8.655031, 8.789314, 8.923654, 9.058049, 9.192499, 9.327003, 
    9.461561, 9.596171, 9.730834, 9.865547, 10.00031, 10.13512, 10.26998, 
    10.40489, 10.53985, 10.67485, 10.8099, 10.94499, 11.08013, 11.21531, 
    11.35053, 11.48579, 11.6211, 11.75644, 11.89182, 12.02724, 12.1627, 
    12.2982, 12.43373, 12.56929, 12.70489, 12.84052, 12.97619, 13.11188, 
    13.24761, 13.38336, 13.51915, 13.65496, 13.7908, 13.92667, 14.06256, 
    14.19848, 14.33442, 14.47039, 14.60637, 14.74238, 14.87841, 15.01446, 
    15.15053, 15.28661, 15.42272, 15.55884, 15.69497, 15.83112, 15.96728, 
    16.10345, 16.23964, 16.37584, 16.51205, 16.64827, 16.78449, 16.92073, 
    17.05697, 17.19322, 17.32947, 17.46573, 17.60199, 17.73825, 17.87451, 
    18.01078, 18.14704, 18.28331, 18.41957, 18.55583, 18.69208, 18.82833, 
    18.96458, 19.10082, 19.23705, 19.37328, 19.5095, 19.6457, 19.7819, 
    19.91809, 20.05426, 20.19042, 20.32657, 20.4627, 20.59881, 20.73491, 
    20.871, 21.00706, 21.14311, 21.27913, 21.41514, 21.55112, 21.68708, 
    21.82302, 21.95893, 22.09482, 22.23069, 22.36652, 22.50233, 22.63811, 
    22.77386, 22.90959, 23.04528, 23.18093, 23.31656, 23.45216, 23.58772, 
    23.72324, 23.85873, 23.99418, 24.12959, 24.26497, 24.40031, 24.5356, 
    24.67086, 24.80608, 24.94125, 25.07638, 25.21146, 25.34651, 25.4815, 
    25.61645, 25.75135, 25.88621, 26.02101, 26.15577, 26.29047, 26.42513, 
    26.55973, 26.69428, 26.82877, 26.96321, 27.0976, 27.23193, 27.36621, 
    27.50042, 27.63458, 27.76868, 27.90272, 28.0367, 28.17062, 28.30448, 
    28.43827, 28.572, 28.70567, 28.83927, 28.97281, 29.10628, 29.23968, 
    29.37301, 29.50628, 29.63947, 29.7726, 29.90566, 30.03864, 30.17156, 
    30.3044, 30.43716, 30.56985, 30.70247, 30.83501, 30.96748, 31.09987, 
    31.23218, 31.36441, 31.49656, 31.62864, 31.76063, 31.89254, 32.02437, 
    32.15612, 32.28778, 32.41937, 32.55087, 32.68228, 32.8136, 32.94484, 
    33.076, 33.20706, 33.33804, 33.46893, 33.59973, 33.73044, 33.86106, 
    33.99158, 34.12202, 34.25237, 34.38261, 34.51277, 34.64283, 34.7728, 
    34.90267, 35.03245, 35.16213, 35.29171, 35.4212, 35.55059, 35.67987, 
    35.80906, 35.93815, 36.06714, 36.19603, 36.32481, 36.4535, 36.58208, 
    36.71056, 36.83894, 36.96721, 37.09537, 37.22343, 37.35139, 37.47924, 
    37.60698, 37.73462, 37.86214, 37.98957, 38.11687, 38.24408, 38.37117, 
    38.49815, 38.62503, 38.75179, 38.87844, 39.00497, 39.1314, 39.25771, 
    39.38391, 39.51, 39.63597, 39.76183, 39.88757, 40.0132, 40.13871, 
    40.26411, 40.38939, 40.51455, 40.6396,
  -15.75332, -15.64021, -15.52696, -15.41358, -15.30005, -15.18639, 
    -15.07259, -14.95866, -14.84458, -14.73037, -14.61602, -14.50154, 
    -14.38692, -14.27216, -14.15726, -14.04223, -13.92706, -13.81175, 
    -13.6963, -13.58072, -13.46501, -13.34915, -13.23317, -13.11704, 
    -13.00078, -12.88438, -12.76785, -12.65118, -12.53438, -12.41744, 
    -12.30036, -12.18316, -12.06581, -11.94833, -11.83072, -11.71297, 
    -11.59509, -11.47707, -11.35892, -11.24064, -11.12222, -11.00367, 
    -10.88499, -10.76617, -10.64722, -10.52814, -10.40892, -10.28958, 
    -10.1701, -10.05049, -9.930742, -9.810868, -9.690864, -9.570727, 
    -9.45046, -9.330063, -9.209535, -9.088878, -8.96809, -8.847173, 
    -8.726127, -8.604951, -8.483647, -8.362214, -8.240654, -8.118965, 
    -7.997149, -7.875205, -7.753134, -7.630936, -7.508612, -7.386161, 
    -7.263585, -7.140882, -7.018055, -6.895103, -6.772026, -6.648824, 
    -6.525498, -6.40205, -6.278477, -6.154781, -6.030962, -5.907022, 
    -5.782959, -5.658774, -5.534469, -5.410042, -5.285495, -5.160828, 
    -5.03604, -4.911133, -4.786108, -4.660963, -4.5357, -4.41032, -4.284822, 
    -4.159206, -4.033474, -3.907626, -3.781662, -3.655583, -3.529388, 
    -3.403079, -3.276656, -3.150119, -3.023468, -2.896705, -2.76983, 
    -2.642843, -2.515744, -2.388534, -2.261214, -2.133783, -2.006243, 
    -1.878594, -1.750836, -1.62297, -1.494997, -1.366916, -1.238729, 
    -1.110435, -0.9820362, -0.8535319, -0.724923, -0.59621, -0.4673934, 
    -0.3384738, -0.2094516, -0.08032748, 0.04889809, 0.1782245, 0.3076514, 
    0.437178, 0.5668038, 0.6965283, 0.826351, 0.9562712, 1.086288, 1.216402, 
    1.346611, 1.476916, 1.607315, 1.737808, 1.868395, 1.999075, 2.129847, 
    2.26071, 2.391665, 2.52271, 2.653844, 2.785068, 2.916381, 3.047781, 
    3.179269, 3.310843, 3.442504, 3.574249, 3.70608, 3.837994, 3.969992, 
    4.102073, 4.234236, 4.36648, 4.498805, 4.63121, 4.763694, 4.896257, 
    5.028898, 5.161617, 5.294412, 5.427283, 5.56023, 5.693251, 5.826345, 
    5.959513, 6.092753, 6.226066, 6.359449, 6.492902, 6.626425, 6.760017, 
    6.893677, 7.027404, 7.161198, 7.295058, 7.428983, 7.562973, 7.697025, 
    7.831141, 7.96532, 8.099559, 8.233859, 8.368219, 8.502639, 8.637116, 
    8.771651, 8.906243, 9.040891, 9.175594, 9.310351, 9.445163, 9.580028, 
    9.714944, 9.849912, 9.98493, 10.12, 10.25511, 10.39028, 10.52549, 
    10.66075, 10.79605, 10.93141, 11.0668, 11.20224, 11.33771, 11.47324, 
    11.6088, 11.7444, 11.88004, 12.01572, 12.15144, 12.28719, 12.42298, 
    12.5588, 12.69466, 12.83055, 12.96648, 13.10244, 13.23842, 13.37444, 
    13.51049, 13.64656, 13.78266, 13.91879, 14.05495, 14.19113, 14.32733, 
    14.46356, 14.59981, 14.73608, 14.87237, 15.00868, 15.14501, 15.28136, 
    15.41772, 15.55411, 15.6905, 15.82692, 15.96334, 16.09978, 16.23623, 
    16.37269, 16.50917, 16.64565, 16.78214, 16.91864, 17.05514, 17.19165, 
    17.32817, 17.46469, 17.60122, 17.73774, 17.87427, 18.0108, 18.14733, 
    18.28386, 18.42038, 18.55691, 18.69342, 18.82994, 18.96645, 19.10295, 
    19.23945, 19.37594, 19.51242, 19.64889, 19.78535, 19.9218, 20.05824, 
    20.19466, 20.33107, 20.46747, 20.60385, 20.74021, 20.87656, 21.01288, 
    21.14919, 21.28548, 21.42175, 21.55799, 21.69422, 21.83042, 21.96659, 
    22.10274, 22.23887, 22.37497, 22.51104, 22.64708, 22.78309, 22.91907, 
    23.05502, 23.19094, 23.32683, 23.46268, 23.5985, 23.73429, 23.87004, 
    24.00574, 24.14142, 24.27705, 24.41265, 24.5482, 24.68372, 24.81919, 
    24.95462, 25.09001, 25.22535, 25.36065, 25.4959, 25.63111, 25.76626, 
    25.90137, 26.03643, 26.17144, 26.3064, 26.44131, 26.57617, 26.71097, 
    26.84572, 26.98041, 27.11505, 27.24963, 27.38416, 27.51863, 27.65304, 
    27.78739, 27.92168, 28.05591, 28.19008, 28.32418, 28.45823, 28.59221, 
    28.72612, 28.85997, 28.99375, 29.12747, 29.26112, 29.3947, 29.52821, 
    29.66166, 29.79503, 29.92833, 30.06156, 30.19471, 30.3278, 30.46081, 
    30.59374, 30.7266, 30.85938, 30.99209, 31.12472, 31.25727, 31.38974, 
    31.52213, 31.65444, 31.78668, 31.91883, 32.05089, 32.18288, 32.31478, 
    32.4466, 32.57833, 32.70998, 32.84154, 32.97301, 33.1044, 33.23569, 
    33.36691, 33.49802, 33.62906, 33.76, 33.89085, 34.0216, 34.15227, 
    34.28284, 34.41332, 34.5437, 34.67399, 34.80419, 34.93428, 35.06429, 
    35.19419, 35.324, 35.45371, 35.58332, 35.71283, 35.84224, 35.97155, 
    36.10076, 36.22987, 36.35888, 36.48778, 36.61658, 36.74527, 36.87387, 
    37.00235, 37.13074, 37.25901, 37.38718, 37.51525, 37.6432, 37.77105, 
    37.89879, 38.02642, 38.15395, 38.28136, 38.40866, 38.53586, 38.66294, 
    38.78991, 38.91676, 39.04351, 39.17014, 39.29666, 39.42307, 39.54936, 
    39.67553, 39.80159, 39.92754, 40.05337, 40.17908, 40.30468, 40.43016, 
    40.55552, 40.68077,
  -15.81028, -15.69703, -15.58364, -15.47011, -15.35645, -15.24264, -15.1287, 
    -15.01462, -14.9004, -14.78605, -14.67155, -14.55692, -14.44215, 
    -14.32725, -14.2122, -14.09702, -13.9817, -13.86625, -13.75065, 
    -13.63492, -13.51905, -13.40305, -13.28691, -13.17063, -13.05421, 
    -12.93766, -12.82097, -12.70415, -12.58719, -12.47009, -12.35286, 
    -12.23549, -12.11799, -12.00035, -11.88258, -11.76467, -11.64663, 
    -11.52845, -11.41014, -11.29169, -11.17311, -11.05439, -10.93554, 
    -10.81656, -10.69744, -10.57819, -10.45881, -10.33929, -10.21964, 
    -10.09986, -9.979948, -9.859902, -9.739725, -9.619416, -9.498976, 
    -9.378405, -9.257702, -9.136869, -9.015905, -8.894812, -8.773588, 
    -8.652235, -8.530752, -8.409141, -8.2874, -8.16553, -8.043532, -7.921407, 
    -7.799154, -7.676773, -7.554265, -7.43163, -7.308868, -7.18598, 
    -7.062966, -6.939826, -6.816562, -6.693172, -6.569657, -6.446018, 
    -6.322255, -6.198368, -6.074358, -5.950225, -5.825969, -5.701591, 
    -5.577091, -5.45247, -5.327727, -5.202863, -5.077879, -4.952775, 
    -4.827551, -4.702208, -4.576746, -4.451165, -4.325466, -4.19965, 
    -4.073716, -3.947665, -3.821498, -3.695214, -3.568815, -3.442301, 
    -3.315672, -3.188929, -3.062072, -2.935101, -2.808018, -2.680821, 
    -2.553513, -2.426093, -2.298563, -2.170921, -2.043169, -1.915307, 
    -1.787336, -1.659257, -1.531069, -1.402773, -1.274371, -1.145861, 
    -1.017245, -0.8885237, -0.7596969, -0.6307654, -0.5017298, -0.3725906, 
    -0.2433482, -0.1140033, 0.01544359, 0.144992, 0.2746413, 0.404391, 
    0.5342404, 0.6641892, 0.7942365, 0.924382, 1.054625, 1.184965, 1.315401, 
    1.445934, 1.576561, 1.707283, 1.838099, 1.969008, 2.10001, 2.231104, 
    2.36229, 2.493567, 2.624934, 2.756391, 2.887937, 3.019571, 3.151293, 
    3.283103, 3.414998, 3.54698, 3.679047, 3.811198, 3.943434, 4.075752, 
    4.208153, 4.340636, 4.473201, 4.605845, 4.73857, 4.871374, 5.004256, 
    5.137217, 5.270254, 5.403368, 5.536557, 5.669821, 5.80316, 5.936573, 
    6.070058, 6.203615, 6.337244, 6.470943, 6.604712, 6.738552, 6.872458, 
    7.006433, 7.140476, 7.274584, 7.408758, 7.542997, 7.677299, 7.811666, 
    7.946094, 8.080585, 8.215136, 8.349748, 8.484419, 8.619148, 8.753936, 
    8.888781, 9.023682, 9.158639, 9.293651, 9.428717, 9.563835, 9.699006, 
    9.834229, 9.969503, 10.10483, 10.2402, 10.37562, 10.51109, 10.64661, 
    10.78217, 10.91778, 11.05343, 11.18912, 11.32486, 11.46064, 11.59646, 
    11.73232, 11.86822, 12.00416, 12.14014, 12.27615, 12.4122, 12.54829, 
    12.68441, 12.82056, 12.95674, 13.09296, 13.22921, 13.36549, 13.5018, 
    13.63813, 13.7745, 13.91089, 14.04731, 14.18375, 14.32022, 14.45671, 
    14.59322, 14.72975, 14.86631, 15.00288, 15.13948, 15.27609, 15.41272, 
    15.54937, 15.68603, 15.8227, 15.95939, 16.0961, 16.23281, 16.36954, 
    16.50628, 16.64302, 16.77978, 16.91654, 17.05331, 17.19009, 17.32687, 
    17.46365, 17.60044, 17.73723, 17.87403, 18.01082, 18.14761, 18.28441, 
    18.4212, 18.55799, 18.69477, 18.83155, 18.96833, 19.10509, 19.24186, 
    19.37861, 19.51536, 19.65209, 19.78882, 19.92553, 20.06223, 20.19892, 
    20.33559, 20.47225, 20.60889, 20.74552, 20.88213, 21.01872, 21.15529, 
    21.29185, 21.42838, 21.56489, 21.70137, 21.83784, 21.97427, 22.11069, 
    22.24707, 22.38343, 22.51977, 22.65607, 22.79234, 22.92859, 23.0648, 
    23.20098, 23.33713, 23.47324, 23.60932, 23.74537, 23.88137, 24.01735, 
    24.15328, 24.28917, 24.42503, 24.56084, 24.69662, 24.83235, 24.96803, 
    25.10368, 25.23928, 25.37483, 25.51034, 25.6458, 25.78122, 25.91658, 
    26.0519, 26.18716, 26.32238, 26.45754, 26.59265, 26.72771, 26.86271, 
    26.99766, 27.13255, 27.26739, 27.40217, 27.53689, 27.67155, 27.80615, 
    27.94069, 28.07517, 28.20959, 28.34395, 28.47824, 28.61247, 28.74663, 
    28.88073, 29.01476, 29.14873, 29.28263, 29.41645, 29.55021, 29.6839, 
    29.81752, 29.95106, 30.08454, 30.21794, 30.35126, 30.48452, 30.61769, 
    30.7508, 30.88382, 31.01677, 31.14964, 31.28243, 31.41514, 31.54778, 
    31.68033, 31.8128, 31.94518, 32.07749, 32.20971, 32.34185, 32.4739, 
    32.60587, 32.73775, 32.86955, 33.00126, 33.13288, 33.26441, 33.39585, 
    33.52721, 33.65847, 33.78964, 33.92072, 34.0517, 34.1826, 34.3134, 
    34.44411, 34.57472, 34.70524, 34.83566, 34.96598, 35.09621, 35.22634, 
    35.35637, 35.48631, 35.61614, 35.74587, 35.87551, 36.00504, 36.13447, 
    36.2638, 36.39302, 36.52215, 36.65117, 36.78008, 36.90889, 37.0376, 
    37.16619, 37.29469, 37.42308, 37.55135, 37.67952, 37.80759, 37.93554, 
    38.06339, 38.19112, 38.31874, 38.44626, 38.57366, 38.70095, 38.82813, 
    38.95519, 39.08215, 39.20898, 39.33571, 39.46232, 39.58882, 39.7152, 
    39.84146, 39.96761, 40.09364, 40.21956, 40.34536, 40.47104, 40.5966, 
    40.72204,
  -15.86735, -15.75396, -15.64043, -15.52676, -15.41296, -15.29901, 
    -15.18493, -15.07071, -14.95634, -14.84184, -14.72721, -14.61243, 
    -14.49751, -14.38246, -14.26727, -14.15194, -14.03647, -13.92086, 
    -13.80512, -13.68924, -13.57322, -13.45706, -13.34077, -13.22434, 
    -13.10777, -12.99106, -12.87422, -12.75724, -12.64012, -12.52287, 
    -12.40548, -12.28795, -12.17029, -12.05249, -11.93456, -11.81649, 
    -11.69828, -11.57994, -11.46147, -11.34285, -11.22411, -11.10523, 
    -10.98621, -10.86706, -10.74778, -10.62836, -10.50881, -10.38913, 
    -10.26931, -10.14936, -10.02927, -9.909055, -9.788705, -9.668223, 
    -9.547609, -9.426864, -9.305986, -9.184978, -9.063838, -8.942567, 
    -8.821166, -8.699635, -8.577973, -8.456182, -8.334261, -8.212211, 
    -8.090032, -7.967724, -7.845288, -7.722723, -7.600031, -7.477211, 
    -7.354264, -7.23119, -7.107989, -6.984663, -6.86121, -6.737631, 
    -6.613927, -6.490098, -6.366145, -6.242066, -6.117865, -5.993539, 
    -5.86909, -5.744518, -5.619823, -5.495007, -5.370068, -5.245008, 
    -5.119826, -4.994524, -4.869102, -4.74356, -4.617898, -4.492117, 
    -4.366217, -4.240199, -4.114063, -3.987809, -3.861438, -3.734951, 
    -3.608347, -3.481627, -3.354792, -3.227842, -3.100778, -2.973599, 
    -2.846307, -2.718902, -2.591384, -2.463753, -2.336011, -2.208158, 
    -2.080194, -1.952119, -1.823935, -1.695641, -1.567239, -1.438728, 
    -1.310109, -1.181383, -1.05255, -0.9236109, -0.7945658, -0.6654155, 
    -0.5361603, -0.406801, -0.277338, -0.1477719, -0.01810312, 0.1116677, 
    0.24154, 0.3715132, 0.5015868, 0.6317602, 0.7620329, 0.8924042, 1.022874, 
    1.15344, 1.284104, 1.414865, 1.54572, 1.676672, 1.807717, 1.938857, 
    2.07009, 2.201415, 2.332833, 2.464342, 2.595942, 2.727632, 2.859412, 
    2.991281, 3.123238, 3.255283, 3.387415, 3.519633, 3.651937, 3.784326, 
    3.916799, 4.049356, 4.181996, 4.314719, 4.447523, 4.580408, 4.713374, 
    4.846419, 4.979543, 5.112746, 5.246026, 5.379383, 5.512816, 5.646324, 
    5.779908, 5.913565, 6.047296, 6.181099, 6.314974, 6.44892, 6.582937, 
    6.717023, 6.851178, 6.985402, 7.119693, 7.25405, 7.388474, 7.522962, 
    7.657516, 7.792132, 7.926812, 8.061554, 8.196357, 8.331221, 8.466145, 
    8.601128, 8.736169, 8.871267, 9.006422, 9.141633, 9.2769, 9.412221, 
    9.547595, 9.683022, 9.818501, 9.954031, 10.08961, 10.22524, 10.36092, 
    10.49665, 10.63242, 10.76824, 10.90411, 11.04002, 11.17597, 11.31197, 
    11.44801, 11.58409, 11.72021, 11.85637, 11.99257, 12.1288, 12.26508, 
    12.40139, 12.53774, 12.67412, 12.81053, 12.94698, 13.08346, 13.21997, 
    13.35651, 13.49308, 13.62968, 13.76631, 13.90296, 14.03965, 14.17635, 
    14.31308, 14.44983, 14.58661, 14.72341, 14.86023, 14.99707, 15.13393, 
    15.2708, 15.4077, 15.54461, 15.68153, 15.81848, 15.95543, 16.0924, 
    16.22938, 16.36637, 16.50337, 16.64039, 16.77741, 16.91444, 17.05147, 
    17.18851, 17.32556, 17.46261, 17.59966, 17.73672, 17.87378, 18.01084, 
    18.1479, 18.28496, 18.42202, 18.55907, 18.69612, 18.83317, 18.97021, 
    19.10724, 19.24427, 19.38129, 19.5183, 19.6553, 19.79229, 19.92927, 
    20.06623, 20.20319, 20.34013, 20.47705, 20.61396, 20.75085, 20.88772, 
    21.02458, 21.16142, 21.29823, 21.43503, 21.5718, 21.70855, 21.84528, 
    21.98198, 22.11865, 22.2553, 22.39193, 22.52852, 22.66509, 22.80163, 
    22.93813, 23.07461, 23.21105, 23.34746, 23.48383, 23.62017, 23.75648, 
    23.89275, 24.02898, 24.16517, 24.30133, 24.43744, 24.57352, 24.70955, 
    24.84554, 24.98149, 25.11739, 25.25325, 25.38906, 25.52483, 25.66055, 
    25.79622, 25.93184, 26.06741, 26.20293, 26.3384, 26.47382, 26.60919, 
    26.7445, 26.87976, 27.01496, 27.15011, 27.2852, 27.42023, 27.5552, 
    27.69012, 27.82497, 27.95976, 28.0945, 28.22917, 28.36377, 28.49832, 
    28.6328, 28.76721, 28.90155, 29.03584, 29.17005, 29.30419, 29.43827, 
    29.57227, 29.70621, 29.84007, 29.97386, 30.10758, 30.24123, 30.3748, 
    30.5083, 30.64172, 30.77506, 30.90833, 31.04152, 31.17463, 31.30766, 
    31.44062, 31.57349, 31.70628, 31.83899, 31.97162, 32.10416, 32.23662, 
    32.369, 32.50129, 32.63349, 32.76561, 32.89764, 33.02958, 33.16144, 
    33.29321, 33.42488, 33.55647, 33.68796, 33.81937, 33.95068, 34.08189, 
    34.21302, 34.34405, 34.47499, 34.60583, 34.73657, 34.86722, 34.99777, 
    35.12822, 35.25858, 35.38884, 35.519, 35.64905, 35.77901, 35.90887, 
    36.03862, 36.16827, 36.29782, 36.42727, 36.55661, 36.68585, 36.81499, 
    36.94402, 37.07294, 37.20175, 37.33046, 37.45906, 37.58756, 37.71594, 
    37.84422, 37.97239, 38.10044, 38.22839, 38.35622, 38.48395, 38.61156, 
    38.73906, 38.86645, 38.99372, 39.12088, 39.24793, 39.37486, 39.50168, 
    39.62838, 39.75497, 39.88144, 40.00779, 40.13402, 40.26014, 40.38614, 
    40.51202, 40.63778, 40.76343,
  -15.92455, -15.81102, -15.69735, -15.58354, -15.46959, -15.3555, -15.24128, 
    -15.12691, -15.01241, -14.89776, -14.78298, -14.66806, -14.553, 
    -14.43779, -14.32246, -14.20698, -14.09136, -13.9756, -13.85971, 
    -13.74368, -13.62751, -13.5112, -13.39475, -13.27817, -13.16144, 
    -13.04458, -12.92758, -12.81045, -12.69317, -12.57576, -12.45822, 
    -12.34053, -12.22271, -12.10475, -11.98666, -11.86843, -11.75006, 
    -11.63156, -11.51292, -11.39414, -11.27523, -11.15619, -11.037, 
    -10.91769, -10.79824, -10.67865, -10.55893, -10.43908, -10.31909, 
    -10.19897, -10.07871, -9.958324, -9.837802, -9.717147, -9.596359, 
    -9.47544, -9.354387, -9.233203, -9.111887, -8.990439, -8.86886, -8.74715, 
    -8.62531, -8.503339, -8.381238, -8.259007, -8.136646, -8.014155, 
    -7.891537, -7.768788, -7.645912, -7.522907, -7.399775, -7.276514, 
    -7.153127, -7.029612, -6.905971, -6.782203, -6.658309, -6.53429, 
    -6.410146, -6.285876, -6.161482, -6.036963, -5.912321, -5.787555, 
    -5.662665, -5.537653, -5.412518, -5.287261, -5.161882, -5.036382, 
    -4.910761, -4.785019, -4.659157, -4.533176, -4.407074, -4.280854, 
    -4.154516, -4.028059, -3.901484, -3.774792, -3.647983, -3.521058, 
    -3.394016, -3.266859, -3.139587, -3.0122, -2.884699, -2.757084, 
    -2.629356, -2.501515, -2.373561, -2.245496, -2.117319, -1.989031, 
    -1.860633, -1.732125, -1.603507, -1.47478, -1.345945, -1.217002, 
    -1.087952, -0.9587942, -0.8295304, -0.7001606, -0.5706856, -0.4411057, 
    -0.3114216, -0.1816337, -0.05174263, 0.07825106, 0.2083468, 0.3385441, 
    0.4688423, 0.599241, 0.7297394, 0.860337, 0.9910333, 1.121828, 1.25272, 
    1.383708, 1.514793, 1.645974, 1.77725, 1.90862, 2.040085, 2.171642, 
    2.303292, 2.435034, 2.566868, 2.698792, 2.830806, 2.96291, 3.095103, 
    3.227384, 3.359752, 3.492207, 3.624749, 3.757376, 3.890088, 4.022884, 
    4.155764, 4.288726, 4.421771, 4.554897, 4.688105, 4.821392, 4.954759, 
    5.088204, 5.221727, 5.355328, 5.489006, 5.622759, 5.756588, 5.890491, 
    6.024467, 6.158517, 6.292639, 6.426833, 6.561097, 6.695432, 6.829835, 
    6.964308, 7.098848, 7.233456, 7.36813, 7.502869, 7.637673, 7.772542, 
    7.907473, 8.042467, 8.177523, 8.312639, 8.447817, 8.583054, 8.718349, 
    8.853702, 8.989111, 9.124578, 9.260099, 9.395676, 9.531306, 9.666989, 
    9.802725, 9.938512, 10.07435, 10.21024, 10.34617, 10.48216, 10.61819, 
    10.75427, 10.89039, 11.02656, 11.16278, 11.29903, 11.43533, 11.57167, 
    11.70806, 11.84448, 11.98094, 12.11744, 12.25397, 12.39055, 12.52715, 
    12.6638, 12.80048, 12.93719, 13.07393, 13.2107, 13.34751, 13.48434, 
    13.6212, 13.7581, 13.89501, 14.03196, 14.16893, 14.30592, 14.44294, 
    14.57998, 14.71705, 14.85413, 14.99124, 15.12836, 15.2655, 15.40266, 
    15.53984, 15.67703, 15.81424, 15.95146, 16.08869, 16.22594, 16.3632, 
    16.50047, 16.63774, 16.77503, 16.91232, 17.04963, 17.18694, 17.32425, 
    17.46157, 17.59889, 17.73621, 17.87354, 18.01086, 18.14819, 18.28551, 
    18.42284, 18.56016, 18.69747, 18.83479, 18.97209, 19.10939, 19.24669, 
    19.38397, 19.52125, 19.65852, 19.79577, 19.93302, 20.07025, 20.20747, 
    20.34467, 20.48186, 20.61904, 20.75619, 20.89333, 21.03045, 21.16755, 
    21.30464, 21.4417, 21.57873, 21.71575, 21.85274, 21.9897, 22.12665, 
    22.26356, 22.40045, 22.53731, 22.67414, 22.81094, 22.9477, 23.08444, 
    23.22115, 23.35782, 23.49446, 23.63106, 23.76763, 23.90416, 24.04065, 
    24.1771, 24.31352, 24.4499, 24.58623, 24.72252, 24.85877, 24.99498, 
    25.13114, 25.26726, 25.40333, 25.53935, 25.67533, 25.81126, 25.94714, 
    26.08297, 26.21875, 26.35448, 26.49015, 26.62577, 26.76134, 26.89685, 
    27.03231, 27.16771, 27.30306, 27.43834, 27.57357, 27.70874, 27.84385, 
    27.97889, 28.11387, 28.2488, 28.38366, 28.51845, 28.65318, 28.78784, 
    28.92244, 29.05697, 29.19143, 29.32582, 29.46015, 29.5944, 29.72858, 
    29.86269, 29.99673, 30.1307, 30.26459, 30.3984, 30.53214, 30.66581, 
    30.7994, 30.93291, 31.06634, 31.1997, 31.33297, 31.46617, 31.59928, 
    31.73231, 31.86526, 31.99813, 32.13091, 32.26361, 32.39622, 32.52875, 
    32.66119, 32.79355, 32.92582, 33.05799, 33.19008, 33.32208, 33.45399, 
    33.58581, 33.71754, 33.84917, 33.98072, 34.11217, 34.24352, 34.37478, 
    34.50595, 34.63702, 34.76799, 34.89887, 35.02965, 35.16033, 35.29091, 
    35.42139, 35.55178, 35.68206, 35.81224, 35.94232, 36.0723, 36.20217, 
    36.33194, 36.46161, 36.59118, 36.72063, 36.84998, 36.97923, 37.10837, 
    37.23741, 37.36633, 37.49515, 37.62386, 37.75246, 37.88095, 38.00933, 
    38.1376, 38.26576, 38.39381, 38.52174, 38.64957, 38.77728, 38.90488, 
    39.03236, 39.15973, 39.28698, 39.41412, 39.54114, 39.66805, 39.79484, 
    39.92151, 40.04807, 40.17451, 40.30083, 40.42703, 40.55311, 40.67907, 
    40.80492,
  -15.98186, -15.86819, -15.75439, -15.64044, -15.52635, -15.41212, 
    -15.29775, -15.18324, -15.06859, -14.9538, -14.83887, -14.72381, 
    -14.6086, -14.49325, -14.37776, -14.26214, -14.14637, -14.03047, 
    -13.91442, -13.79824, -13.68192, -13.56546, -13.44886, -13.33212, 
    -13.21524, -13.09822, -12.98107, -12.86378, -12.74635, -12.62878, 
    -12.51108, -12.39323, -12.27525, -12.15713, -12.03888, -11.92049, 
    -11.80196, -11.68329, -11.56449, -11.44555, -11.32647, -11.20726, 
    -11.08792, -10.96843, -10.84882, -10.72906, -10.60917, -10.48915, 
    -10.36899, -10.2487, -10.12827, -10.00771, -9.887018, -9.766191, 
    -9.645228, -9.524134, -9.402906, -9.281547, -9.160053, -9.038429, 
    -8.916672, -8.794784, -8.672764, -8.550613, -8.428331, -8.305919, 
    -8.183376, -8.060703, -7.937901, -7.814969, -7.691908, -7.568718, 
    -7.445399, -7.321952, -7.198378, -7.074675, -6.950845, -6.826889, 
    -6.702805, -6.578595, -6.454259, -6.329798, -6.205211, -6.0805, 
    -5.955663, -5.830702, -5.705618, -5.58041, -5.455079, -5.329624, 
    -5.204048, -5.07835, -4.952529, -4.826588, -4.700525, -4.574343, 
    -4.44804, -4.321617, -4.195076, -4.068415, -3.941636, -3.814739, 
    -3.687725, -3.560593, -3.433345, -3.30598, -3.1785, -3.050905, -2.923194, 
    -2.795369, -2.66743, -2.539378, -2.411212, -2.282935, -2.154545, 
    -2.026043, -1.897431, -1.768707, -1.639874, -1.510931, -1.381879, 
    -1.252719, -1.12345, -0.9940742, -0.8645912, -0.7350016, -0.6053061, 
    -0.4755053, -0.3455995, -0.2155894, -0.08547557, 0.0447415, 0.1750612, 
    0.305483, 0.4360064, 0.5666307, 0.6973554, 0.82818, 0.9591036, 1.090126, 
    1.221246, 1.352464, 1.483779, 1.61519, 1.746697, 1.878298, 2.009995, 
    2.141784, 2.273667, 2.405643, 2.53771, 2.669869, 2.802119, 2.934458, 
    3.066887, 3.199404, 3.33201, 3.464703, 3.597483, 3.730349, 3.8633, 
    3.996336, 4.129456, 4.262659, 4.395945, 4.529313, 4.662762, 4.796292, 
    4.929902, 5.063591, 5.197358, 5.331203, 5.465126, 5.599124, 5.733199, 
    5.867348, 6.001572, 6.135869, 6.270238, 6.40468, 6.539193, 6.673777, 
    6.80843, 6.943152, 7.077942, 7.212801, 7.347725, 7.482716, 7.617772, 
    7.752892, 7.888076, 8.023323, 8.158632, 8.294003, 8.429434, 8.564925, 
    8.700475, 8.836082, 8.971748, 9.107471, 9.243248, 9.379081, 9.514968, 
    9.650908, 9.786901, 9.922947, 10.05904, 10.19519, 10.33138, 10.46763, 
    10.60392, 10.74026, 10.87664, 11.01307, 11.14955, 11.28606, 11.42262, 
    11.55923, 11.69587, 11.83255, 11.96927, 12.10604, 12.24283, 12.37967, 
    12.51654, 12.65345, 12.79039, 12.92736, 13.06437, 13.20141, 13.33847, 
    13.47557, 13.6127, 13.74986, 13.88704, 14.02425, 14.16149, 14.29875, 
    14.43603, 14.57334, 14.71066, 14.84801, 14.98538, 15.12277, 15.26018, 
    15.39761, 15.53505, 15.67251, 15.80998, 15.94747, 16.08497, 16.22249, 
    16.36001, 16.49755, 16.63509, 16.77265, 16.91021, 17.04778, 17.18535, 
    17.32293, 17.46052, 17.59811, 17.7357, 17.87329, 18.01088, 18.14848, 
    18.28607, 18.42366, 18.56125, 18.69883, 18.83641, 18.97399, 19.11155, 
    19.24911, 19.38667, 19.52421, 19.66174, 19.79927, 19.93678, 20.07428, 
    20.21176, 20.34924, 20.48669, 20.62413, 20.76155, 20.89896, 21.03635, 
    21.17371, 21.31106, 21.44839, 21.58569, 21.72297, 21.86023, 21.99746, 
    22.13466, 22.27184, 22.40899, 22.54612, 22.68321, 22.82027, 22.95731, 
    23.09431, 23.23128, 23.36821, 23.50511, 23.64198, 23.77881, 23.9156, 
    24.05236, 24.18907, 24.32575, 24.46239, 24.59898, 24.73553, 24.87205, 
    25.00851, 25.14494, 25.28131, 25.41764, 25.55393, 25.69016, 25.82635, 
    25.96249, 26.09858, 26.23461, 26.3706, 26.50653, 26.64241, 26.77823, 
    26.914, 27.04972, 27.18537, 27.32097, 27.45651, 27.59199, 27.72742, 
    27.86278, 27.99808, 28.13331, 28.26849, 28.4036, 28.53864, 28.67362, 
    28.80854, 28.94338, 29.07816, 29.21288, 29.34752, 29.48209, 29.61659, 
    29.75102, 29.88538, 30.01966, 30.15388, 30.28802, 30.42208, 30.55606, 
    30.68997, 30.82381, 30.95756, 31.09124, 31.22484, 31.35835, 31.49179, 
    31.62514, 31.75842, 31.89161, 32.02472, 32.15774, 32.29068, 32.42353, 
    32.55629, 32.68897, 32.82156, 32.95407, 33.08648, 33.21881, 33.35104, 
    33.48318, 33.61524, 33.7472, 33.87907, 34.01085, 34.14252, 34.27411, 
    34.40561, 34.537, 34.6683, 34.7995, 34.93061, 35.06161, 35.19252, 
    35.32333, 35.45404, 35.58465, 35.71515, 35.84556, 35.97586, 36.10606, 
    36.23616, 36.36615, 36.49604, 36.62583, 36.75551, 36.88508, 37.01455, 
    37.14391, 37.27316, 37.4023, 37.53133, 37.66026, 37.78908, 37.91778, 
    38.04638, 38.17486, 38.30323, 38.4315, 38.55964, 38.68768, 38.8156, 
    38.94341, 39.07109, 39.19867, 39.32613, 39.45348, 39.58071, 39.70782, 
    39.83482, 39.9617, 40.08846, 40.2151, 40.34163, 40.46803, 40.59431, 
    40.72047, 40.84652,
  -16.0393, -15.9255, -15.81155, -15.69746, -15.58323, -15.46886, -15.35435, 
    -15.23969, -15.1249, -15.00997, -14.89489, -14.77968, -14.66433, 
    -14.54883, -14.4332, -14.31742, -14.20151, -14.08545, -13.96926, 
    -13.85292, -13.73645, -13.61984, -13.50308, -13.38619, -13.26916, 
    -13.15199, -13.03468, -12.91723, -12.79965, -12.68192, -12.56406, 
    -12.44605, -12.32791, -12.20964, -12.09122, -11.97267, -11.85398, 
    -11.73515, -11.61618, -11.49708, -11.37784, -11.25846, -11.13895, 
    -11.0193, -10.89951, -10.77959, -10.65954, -10.53934, -10.41901, 
    -10.29855, -10.17795, -10.05722, -9.936354, -9.815352, -9.694217, 
    -9.572948, -9.451545, -9.330009, -9.208339, -9.086536, -8.964602, 
    -8.842535, -8.720335, -8.598004, -8.475542, -8.352948, -8.230223, 
    -8.107368, -7.984382, -7.861266, -7.738019, -7.614644, -7.491139, 
    -7.367506, -7.243743, -7.119853, -6.995834, -6.871688, -6.747415, 
    -6.623014, -6.498487, -6.373833, -6.249053, -6.124148, -5.999117, 
    -5.873962, -5.748682, -5.623278, -5.49775, -5.372098, -5.246324, 
    -5.120426, -4.994407, -4.868265, -4.742002, -4.615618, -4.489113, 
    -4.362488, -4.235743, -4.108879, -3.981895, -3.854793, -3.727572, 
    -3.600234, -3.472779, -3.345206, -3.217518, -3.089713, -2.961793, 
    -2.833757, -2.705608, -2.577344, -2.448966, -2.320475, -2.191872, 
    -2.063156, -1.934329, -1.80539, -1.676341, -1.547181, -1.417912, 
    -1.288534, -1.159047, -1.029452, -0.8997489, -0.7699391, -0.6400227, 
    -0.5100003, -0.3798724, -0.2496397, -0.1193025, 0.01113839, 0.1416826, 
    0.2723294, 0.4030784, 0.5339289, 0.6648805, 0.7959324, 0.927084, 
    1.058335, 1.189684, 1.321132, 1.452677, 1.584319, 1.716057, 1.84789, 
    1.979819, 2.111841, 2.243958, 2.376168, 2.50847, 2.640864, 2.773349, 
    2.905925, 3.03859, 3.171345, 3.304188, 3.437119, 3.570138, 3.703243, 
    3.836434, 3.96971, 4.103071, 4.236516, 4.370043, 4.503654, 4.637345, 
    4.771119, 4.904972, 5.038906, 5.172917, 5.307008, 5.441176, 5.575421, 
    5.709742, 5.844138, 5.978609, 6.113154, 6.247772, 6.382462, 6.517224, 
    6.652057, 6.786961, 6.921933, 7.056974, 7.192084, 7.32726, 7.462503, 
    7.597812, 7.733185, 7.868622, 8.004123, 8.139686, 8.275311, 8.410996, 
    8.546742, 8.682548, 8.818412, 8.954333, 9.090312, 9.226347, 9.362437, 
    9.498582, 9.63478, 9.771031, 9.907334, 10.04369, 10.18009, 10.31655, 
    10.45305, 10.5896, 10.7262, 10.86285, 10.99954, 11.13627, 11.27305, 
    11.40987, 11.54674, 11.68364, 11.82059, 11.95757, 12.0946, 12.23166, 
    12.36876, 12.50589, 12.64306, 12.78027, 12.91751, 13.05478, 13.19208, 
    13.32941, 13.46678, 13.60417, 13.74159, 13.87904, 14.01652, 14.15402, 
    14.29154, 14.42909, 14.56667, 14.70426, 14.84188, 14.97952, 15.11717, 
    15.25485, 15.39254, 15.53025, 15.66798, 15.80572, 15.94347, 16.08124, 
    16.21902, 16.35682, 16.49462, 16.63243, 16.77025, 16.90808, 17.04592, 
    17.18376, 17.32161, 17.45947, 17.59732, 17.73518, 17.87304, 18.0109, 
    18.14877, 18.28663, 18.42448, 18.56234, 18.70019, 18.83804, 18.97588, 
    19.11372, 19.25155, 19.38937, 19.52718, 19.66498, 19.80277, 19.94055, 
    20.07832, 20.21607, 20.35381, 20.49153, 20.62924, 20.76693, 20.9046, 
    21.04226, 21.17989, 21.3175, 21.4551, 21.59266, 21.73021, 21.86773, 
    22.00523, 22.1427, 22.28015, 22.41756, 22.55495, 22.69231, 22.82964, 
    22.96694, 23.1042, 23.24144, 23.37864, 23.5158, 23.65293, 23.79002, 
    23.92708, 24.0641, 24.20108, 24.33801, 24.47491, 24.61177, 24.74859, 
    24.88536, 25.02209, 25.15877, 25.29541, 25.432, 25.56854, 25.70504, 
    25.84149, 25.97788, 26.11423, 26.25052, 26.38677, 26.52296, 26.65909, 
    26.79518, 26.9312, 27.06717, 27.20308, 27.33894, 27.47473, 27.61047, 
    27.74615, 27.88176, 28.01731, 28.15281, 28.28823, 28.4236, 28.5589, 
    28.69413, 28.82929, 28.96439, 29.09942, 29.23438, 29.36928, 29.5041, 
    29.63885, 29.77353, 29.90813, 30.04267, 30.17713, 30.31151, 30.44582, 
    30.58005, 30.71421, 30.84829, 30.98229, 31.11621, 31.25005, 31.38381, 
    31.51749, 31.65108, 31.7846, 31.91803, 32.05138, 32.18464, 32.31782, 
    32.45091, 32.58392, 32.71683, 32.84966, 32.9824, 33.11505, 33.24762, 
    33.38008, 33.51246, 33.64475, 33.77695, 33.90905, 34.04106, 34.17297, 
    34.30479, 34.43651, 34.56814, 34.69967, 34.8311, 34.96243, 35.09367, 
    35.2248, 35.35584, 35.48677, 35.61761, 35.74834, 35.87897, 36.0095, 
    36.13993, 36.27025, 36.40046, 36.53057, 36.66058, 36.79048, 36.92027, 
    37.04996, 37.17954, 37.30901, 37.43837, 37.56762, 37.69676, 37.82579, 
    37.95472, 38.08352, 38.21222, 38.34081, 38.46928, 38.59764, 38.72589, 
    38.85402, 38.98204, 39.10994, 39.23772, 39.36539, 39.49295, 39.62038, 
    39.7477, 39.8749, 40.00199, 40.12896, 40.2558, 40.38253, 40.50913, 
    40.63562, 40.76198, 40.88823,
  -16.09687, -15.98292, -15.86883, -15.7546, -15.64023, -15.52572, -15.41107, 
    -15.29627, -15.18133, -15.06625, -14.95104, -14.83568, -14.72018, 
    -14.60453, -14.48875, -14.37283, -14.25676, -14.14056, -14.02422, 
    -13.90773, -13.79111, -13.67434, -13.55743, -13.44039, -13.3232, 
    -13.20588, -13.08841, -12.97081, -12.85306, -12.73518, -12.61716, 
    -12.499, -12.3807, -12.26226, -12.14368, -12.02497, -11.90612, -11.78712, 
    -11.668, -11.54873, -11.42932, -11.30978, -11.1901, -11.07029, -10.95033, 
    -10.83024, -10.71002, -10.58966, -10.46916, -10.34852, -10.22775, 
    -10.10685, -9.985809, -9.864635, -9.743324, -9.621881, -9.500301, 
    -9.37859, -9.256742, -9.134763, -9.01265, -8.890404, -8.768025, 
    -8.645514, -8.52287, -8.400095, -8.277187, -8.154149, -8.030979, 
    -7.907679, -7.784248, -7.660686, -7.536995, -7.413175, -7.289225, 
    -7.165146, -7.040938, -6.916602, -6.792138, -6.667547, -6.542828, 
    -6.417982, -6.293009, -6.16791, -6.042685, -5.917334, -5.791859, 
    -5.666258, -5.540533, -5.414683, -5.288711, -5.162614, -5.036395, 
    -4.910053, -4.783589, -4.657003, -4.530296, -4.403468, -4.276519, 
    -4.14945, -4.022262, -3.894953, -3.767527, -3.639982, -3.512319, 
    -3.384538, -3.256641, -3.128626, -3.000496, -2.87225, -2.743889, 
    -2.615413, -2.486822, -2.358118, -2.229301, -2.10037, -1.971328, 
    -1.842173, -1.712908, -1.583531, -1.454044, -1.324448, -1.194742, 
    -1.064927, -0.9350042, -0.8049735, -0.6748358, -0.5445914, -0.414241, 
    -0.2837851, -0.1532242, -0.02255888, 0.1082103, 0.2390827, 0.3700578, 
    0.5011351, 0.6323138, 0.7635936, 0.8949738, 1.026454, 1.158033, 1.289711, 
    1.421486, 1.553359, 1.685329, 1.817395, 1.949556, 2.081813, 2.214164, 
    2.346608, 2.479145, 2.611775, 2.744496, 2.877309, 3.010211, 3.143204, 
    3.276286, 3.409456, 3.542714, 3.676059, 3.80949, 3.943007, 4.076609, 
    4.210296, 4.344066, 4.477919, 4.611855, 4.745872, 4.87997, 5.014148, 
    5.148405, 5.282742, 5.417156, 5.551647, 5.686215, 5.820859, 5.955578, 
    6.090372, 6.225239, 6.360178, 6.49519, 6.630274, 6.765428, 6.900651, 
    7.035944, 7.171306, 7.306735, 7.44223, 7.577792, 7.713418, 7.84911, 
    7.984865, 8.120683, 8.256562, 8.392504, 8.528505, 8.664567, 8.800688, 
    8.936866, 9.073102, 9.209394, 9.345742, 9.482145, 9.618603, 9.755113, 
    9.891675, 10.02829, 10.16496, 10.30167, 10.43843, 10.57525, 10.71211, 
    10.84901, 10.98596, 11.12296, 11.26, 11.39709, 11.53421, 11.67138, 
    11.80859, 11.94584, 12.08313, 12.22045, 12.35782, 12.49522, 12.63265, 
    12.77012, 12.90762, 13.04516, 13.18273, 13.32033, 13.45796, 13.59562, 
    13.7333, 13.87102, 14.00876, 14.14653, 14.28432, 14.42214, 14.55998, 
    14.69784, 14.83573, 14.97363, 15.11155, 15.2495, 15.38746, 15.52544, 
    15.66343, 15.80144, 15.93946, 16.0775, 16.21555, 16.35361, 16.49168, 
    16.62976, 16.76785, 16.90595, 17.04406, 17.18217, 17.32029, 17.45841, 
    17.59654, 17.73466, 17.8728, 18.01093, 18.14906, 18.28719, 18.42531, 
    18.56344, 18.70156, 18.83968, 18.97779, 19.11589, 19.25399, 19.39208, 
    19.53016, 19.66823, 19.80629, 19.94434, 20.08237, 20.22039, 20.3584, 
    20.49639, 20.63437, 20.77232, 20.91026, 21.04819, 21.18609, 21.32397, 
    21.46183, 21.59966, 21.73748, 21.87527, 22.01303, 22.15077, 22.28848, 
    22.42616, 22.56382, 22.70144, 22.83904, 22.9766, 23.11413, 23.25163, 
    23.38909, 23.52652, 23.66392, 23.80127, 23.93859, 24.07587, 24.21312, 
    24.35032, 24.48748, 24.6246, 24.76168, 24.89871, 25.0357, 25.17265, 
    25.30955, 25.4464, 25.5832, 25.71996, 25.85667, 25.99332, 26.12993, 
    26.26649, 26.40299, 26.53943, 26.67583, 26.81217, 26.94845, 27.08468, 
    27.22085, 27.35696, 27.49301, 27.629, 27.76494, 27.90081, 28.03661, 
    28.17236, 28.30804, 28.44366, 28.57921, 28.71469, 28.85011, 28.98546, 
    29.12074, 29.25596, 29.3911, 29.52617, 29.66117, 29.7961, 29.93096, 
    30.06574, 30.20045, 30.33508, 30.46963, 30.60411, 30.73851, 30.87284, 
    31.00708, 31.14125, 31.27533, 31.40934, 31.54326, 31.6771, 31.81086, 
    31.94453, 32.07812, 32.21162, 32.34504, 32.47837, 32.61161, 32.74477, 
    32.87784, 33.01082, 33.14371, 33.2765, 33.40921, 33.54183, 33.67435, 
    33.80678, 33.93911, 34.07135, 34.2035, 34.33555, 34.46751, 34.59937, 
    34.73112, 34.86279, 34.99435, 35.12582, 35.25718, 35.38844, 35.51961, 
    35.65067, 35.78163, 35.91248, 36.04324, 36.17389, 36.30443, 36.43487, 
    36.5652, 36.69543, 36.82555, 36.95556, 37.08547, 37.21527, 37.34496, 
    37.47453, 37.604, 37.73336, 37.86261, 37.99175, 38.12077, 38.24968, 
    38.37849, 38.50717, 38.63574, 38.7642, 38.89254, 39.02077, 39.14888, 
    39.27688, 39.40476, 39.53252, 39.66016, 39.78769, 39.9151, 40.04239, 
    40.16956, 40.29661, 40.42354, 40.55035, 40.67704, 40.8036, 40.93005,
  -16.15456, -16.04047, -15.92624, -15.81187, -15.69736, -15.5827, -15.46791, 
    -15.35297, -15.23789, -15.12267, -15.0073, -14.8918, -14.77615, 
    -14.66036, -14.54443, -14.42836, -14.31215, -14.19579, -14.0793, 
    -13.96266, -13.84589, -13.72897, -13.61191, -13.49471, -13.37737, 
    -13.25989, -13.14227, -13.02451, -12.90661, -12.78857, -12.67039, 
    -12.55207, -12.43361, -12.31501, -12.19627, -12.0774, -11.95838, 
    -11.83923, -11.71993, -11.6005, -11.48093, -11.36123, -11.24138, 
    -11.1214, -11.00128, -10.88102, -10.76062, -10.64009, -10.51942, 
    -10.39862, -10.27768, -10.1566, -10.03539, -9.914037, -9.792553, 
    -9.670934, -9.549179, -9.42729, -9.305267, -9.183109, -9.060818, 
    -8.938393, -8.815834, -8.693142, -8.570317, -8.44736, -8.32427, 
    -8.201048, -8.077695, -7.95421, -7.830594, -7.706846, -7.582969, 
    -7.458961, -7.334823, -7.210555, -7.086158, -6.961632, -6.836977, 
    -6.712194, -6.587283, -6.462245, -6.337078, -6.211785, -6.086366, 
    -5.96082, -5.835148, -5.709351, -5.583428, -5.457381, -5.331209, 
    -5.204913, -5.078494, -4.951951, -4.825285, -4.698498, -4.571588, 
    -4.444556, -4.317403, -4.19013, -4.062736, -3.935222, -3.807589, 
    -3.679837, -3.551965, -3.423976, -3.29587, -3.167645, -3.039304, 
    -2.910847, -2.782274, -2.653585, -2.524782, -2.395864, -2.266832, 
    -2.137687, -2.008429, -1.879058, -1.749576, -1.619982, -1.490277, 
    -1.360461, -1.230536, -1.100501, -0.9703576, -0.8401058, -0.7097462, 
    -0.5792794, -0.4487059, -0.3180263, -0.1872411, -0.05635094, 0.07464366, 
    0.2057421, 0.3369439, 0.4682484, 0.599655, 0.7311631, 0.8627723, 
    0.9944817, 1.126291, 1.258199, 1.390206, 1.522311, 1.654514, 1.786812, 
    1.919207, 2.051698, 2.184283, 2.316963, 2.449736, 2.582602, 2.71556, 
    2.84861, 2.98175, 3.114981, 3.248302, 3.381712, 3.51521, 3.648795, 
    3.782468, 3.916226, 4.05007, 4.184, 4.318013, 4.45211, 4.586289, 
    4.720551, 4.854894, 4.989317, 5.123821, 5.258403, 5.393064, 5.527803, 
    5.662619, 5.797512, 5.932479, 6.067522, 6.202639, 6.337828, 6.473091, 
    6.608425, 6.743831, 6.879306, 7.014851, 7.150465, 7.286147, 7.421896, 
    7.557712, 7.693593, 7.829539, 7.965549, 8.101622, 8.237758, 8.373956, 
    8.510214, 8.646532, 8.78291, 8.919346, 9.05584, 9.19239, 9.328998, 
    9.465659, 9.602376, 9.739146, 9.875969, 10.01284, 10.14977, 10.28675, 
    10.42377, 10.56084, 10.69797, 10.83513, 10.97235, 11.10961, 11.24691, 
    11.38426, 11.52165, 11.65908, 11.79656, 11.93407, 12.07162, 12.20921, 
    12.34684, 12.4845, 12.6222, 12.75994, 12.89771, 13.03551, 13.17335, 
    13.31121, 13.44911, 13.58703, 13.72499, 13.86297, 14.00098, 14.13902, 
    14.27708, 14.41516, 14.55327, 14.6914, 14.82955, 14.96773, 15.10592, 
    15.24413, 15.38236, 15.52061, 15.65887, 15.79715, 15.93544, 16.07375, 
    16.21206, 16.3504, 16.48874, 16.62709, 16.76545, 16.90382, 17.04219, 
    17.18057, 17.31896, 17.45735, 17.59575, 17.73415, 17.87255, 18.01095, 
    18.14935, 18.28775, 18.42614, 18.56454, 18.70293, 18.84132, 18.9797, 
    19.11807, 19.25644, 19.3948, 19.53315, 19.67149, 19.80981, 19.94813, 
    20.08644, 20.22473, 20.363, 20.50126, 20.63951, 20.77773, 20.91594, 
    21.05413, 21.1923, 21.33045, 21.46858, 21.60668, 21.74476, 21.88282, 
    22.02085, 22.15886, 22.29683, 22.43479, 22.57271, 22.7106, 22.84846, 
    22.98629, 23.12409, 23.26185, 23.39958, 23.53728, 23.67493, 23.81256, 
    23.95014, 24.08769, 24.22519, 24.36266, 24.50009, 24.63747, 24.77481, 
    24.91211, 25.04936, 25.18657, 25.32373, 25.46084, 25.59791, 25.73493, 
    25.87189, 26.00881, 26.14568, 26.28249, 26.41925, 26.55596, 26.69262, 
    26.82921, 26.96576, 27.10224, 27.23867, 27.37504, 27.51134, 27.64759, 
    27.78378, 27.91991, 28.05597, 28.19197, 28.32791, 28.46378, 28.59958, 
    28.73532, 28.87099, 29.00659, 29.14213, 29.27759, 29.41299, 29.54831, 
    29.68356, 29.81874, 29.95384, 30.08887, 30.22383, 30.35871, 30.49352, 
    30.62824, 30.76289, 30.89746, 31.03195, 31.16636, 31.30069, 31.43494, 
    31.56911, 31.70319, 31.83719, 31.97111, 32.10494, 32.23868, 32.37234, 
    32.50591, 32.6394, 32.77279, 32.9061, 33.03932, 33.17244, 33.30548, 
    33.43842, 33.57127, 33.70403, 33.8367, 33.96926, 34.10174, 34.23412, 
    34.36641, 34.49859, 34.63068, 34.76267, 34.89457, 35.02636, 35.15805, 
    35.28965, 35.42114, 35.55253, 35.68382, 35.815, 35.94608, 36.07706, 
    36.20794, 36.3387, 36.46937, 36.59993, 36.73037, 36.86072, 36.99095, 
    37.12108, 37.25109, 37.381, 37.5108, 37.64049, 37.77007, 37.89953, 
    38.02888, 38.15812, 38.28725, 38.41626, 38.54517, 38.67395, 38.80262, 
    38.93118, 39.05961, 39.18793, 39.31614, 39.44423, 39.5722, 39.70005, 
    39.82779, 39.9554, 40.0829, 40.21027, 40.33752, 40.46466, 40.59167, 
    40.71856, 40.84533, 40.97198,
  -16.21237, -16.09815, -15.98378, -15.86927, -15.75461, -15.63982, 
    -15.52488, -15.4098, -15.29457, -15.1792, -15.06369, -14.94804, 
    -14.83225, -14.71631, -14.60024, -14.48402, -14.36765, -14.25115, 
    -14.13451, -14.01772, -13.90079, -13.78372, -13.66651, -13.54916, 
    -13.43166, -13.31403, -13.19625, -13.07833, -12.96028, -12.84208, 
    -12.72374, -12.60526, -12.48664, -12.36788, -12.24898, -12.12995, 
    -12.01077, -11.89145, -11.77199, -11.6524, -11.53266, -11.41279, 
    -11.29278, -11.17263, -11.05234, -10.93191, -10.81135, -10.69065, 
    -10.56981, -10.44883, -10.32772, -10.20647, -10.08508, -9.963561, 
    -9.841903, -9.720108, -9.598178, -9.476112, -9.353911, -9.231576, 
    -9.109105, -8.986501, -8.863762, -8.74089, -8.617884, -8.494744, 
    -8.371471, -8.248066, -8.124529, -8.000858, -7.877057, -7.753124, 
    -7.629059, -7.504863, -7.380537, -7.256081, -7.131494, -7.006778, 
    -6.881932, -6.756958, -6.631854, -6.506622, -6.381263, -6.255775, 
    -6.130161, -6.004419, -5.878551, -5.752556, -5.626436, -5.50019, 
    -5.373819, -5.247324, -5.120704, -4.99396, -4.867094, -4.740103, 
    -4.61299, -4.485755, -4.358397, -4.230919, -4.10332, -3.975599, 
    -3.847759, -3.719799, -3.59172, -3.463521, -3.335205, -3.20677, 
    -3.078219, -2.94955, -2.820765, -2.691863, -2.562846, -2.433714, 
    -2.304467, -2.175107, -2.045632, -1.916045, -1.786345, -1.656533, 
    -1.526609, -1.396575, -1.26643, -1.136174, -1.00581, -0.8753363, 
    -0.7447544, -0.6140646, -0.4832676, -0.3523639, -0.2213539, -0.09023842, 
    0.04098215, 0.1723072, 0.3037361, 0.4352683, 0.5669033, 0.6986404, 
    0.830479, 0.9624186, 1.094459, 1.226598, 1.358837, 1.491174, 1.62361, 
    1.756142, 1.888771, 2.021496, 2.154317, 2.287232, 2.420241, 2.553344, 
    2.68654, 2.819828, 2.953207, 3.086677, 3.220237, 3.353887, 3.487625, 
    3.621452, 3.755366, 3.889367, 4.023454, 4.157626, 4.291883, 4.426224, 
    4.560648, 4.695155, 4.829743, 4.964413, 5.099163, 5.233993, 5.368902, 
    5.503889, 5.638953, 5.774094, 5.909311, 6.044604, 6.179971, 6.315412, 
    6.450925, 6.586511, 6.722168, 6.857897, 6.993695, 7.129562, 7.265498, 
    7.401501, 7.537571, 7.673707, 7.809908, 7.946174, 8.082504, 8.218896, 
    8.35535, 8.491866, 8.628443, 8.765079, 8.901772, 9.038526, 9.175335, 
    9.312201, 9.449123, 9.5861, 9.72313, 9.860214, 9.99735, 10.13454, 
    10.27177, 10.40906, 10.5464, 10.68378, 10.82121, 10.95869, 11.09622, 
    11.23378, 11.37139, 11.50905, 11.64675, 11.78448, 11.92226, 12.06008, 
    12.19794, 12.33583, 12.47376, 12.61173, 12.74973, 12.88776, 13.02583, 
    13.16393, 13.30207, 13.44023, 13.57843, 13.71665, 13.8549, 13.99318, 
    14.13148, 14.26981, 14.40816, 14.54654, 14.68494, 14.82336, 14.9618, 
    15.10026, 15.23875, 15.37724, 15.51576, 15.65429, 15.79284, 15.93141, 
    16.06998, 16.20857, 16.34717, 16.48578, 16.6244, 16.76303, 16.90167, 
    17.04032, 17.17897, 17.31763, 17.45629, 17.59496, 17.73363, 17.8723, 
    18.01097, 18.14964, 18.28831, 18.42698, 18.56564, 18.7043, 18.84296, 
    18.98161, 19.12026, 19.25889, 19.39752, 19.53614, 19.67475, 19.81335, 
    19.95194, 20.09051, 20.22907, 20.36762, 20.50615, 20.64466, 20.78316, 
    20.92164, 21.0601, 21.19854, 21.33696, 21.47535, 21.61373, 21.75208, 
    21.8904, 22.0287, 22.16697, 22.30522, 22.44344, 22.58162, 22.71978, 
    22.85791, 22.99601, 23.13407, 23.2721, 23.4101, 23.54806, 23.68599, 
    23.82387, 23.96172, 24.09953, 24.23731, 24.37504, 24.51273, 24.65038, 
    24.78798, 24.92554, 25.06306, 25.20053, 25.33795, 25.47533, 25.61266, 
    25.74994, 25.88717, 26.02435, 26.16147, 26.29855, 26.43557, 26.57254, 
    26.70945, 26.84631, 26.98311, 27.11985, 27.25654, 27.39317, 27.52973, 
    27.66624, 27.80268, 27.93907, 28.07538, 28.21164, 28.34783, 28.48396, 
    28.62002, 28.75601, 28.89194, 29.02779, 29.16358, 29.2993, 29.43494, 
    29.57052, 29.70602, 29.84145, 29.9768, 30.11208, 30.24729, 30.38242, 
    30.51747, 30.65244, 30.78734, 30.92216, 31.05689, 31.19155, 31.32613, 
    31.46062, 31.59503, 31.72936, 31.8636, 31.99776, 32.13184, 32.26582, 
    32.39972, 32.53354, 32.66726, 32.8009, 32.93444, 33.0679, 33.20126, 
    33.33454, 33.46772, 33.6008, 33.7338, 33.8667, 33.9995, 34.13221, 
    34.26483, 34.39735, 34.52977, 34.66209, 34.79431, 34.92643, 35.05846, 
    35.19038, 35.3222, 35.45393, 35.58554, 35.71706, 35.84847, 35.97978, 
    36.11098, 36.24208, 36.37308, 36.50396, 36.63475, 36.76542, 36.89598, 
    37.02644, 37.15679, 37.28703, 37.41715, 37.54717, 37.67707, 37.80687, 
    37.93655, 38.06612, 38.19558, 38.32492, 38.45415, 38.58326, 38.71226, 
    38.84114, 38.96991, 39.09856, 39.2271, 39.35551, 39.48381, 39.61199, 
    39.74005, 39.86799, 39.99581, 40.12351, 40.25109, 40.37855, 40.50589, 
    40.63311, 40.7602, 40.88717, 41.01402,
  -16.27031, -16.15595, -16.04144, -15.92679, -15.81199, -15.69705, 
    -15.58197, -15.46675, -15.35138, -15.23587, -15.12021, -15.00442, 
    -14.88848, -14.77239, -14.65617, -14.5398, -14.42329, -14.30663, 
    -14.18984, -14.0729, -13.95582, -13.8386, -13.72123, -13.60373, 
    -13.48608, -13.36829, -13.25036, -13.13228, -13.01407, -12.89571, 
    -12.77722, -12.65858, -12.5398, -12.42088, -12.30182, -12.18262, 
    -12.06328, -11.9438, -11.82418, -11.70442, -11.58452, -11.46448, 
    -11.3443, -11.22398, -11.10353, -10.98293, -10.8622, -10.74133, 
    -10.62032, -10.49917, -10.37789, -10.25646, -10.1349, -10.01321, 
    -9.891375, -9.769404, -9.647298, -9.525056, -9.402678, -9.280164, 
    -9.157515, -9.03473, -8.911811, -8.788757, -8.66557, -8.542248, 
    -8.418793, -8.295204, -8.171482, -8.047626, -7.923639, -7.79952, 
    -7.675268, -7.550884, -7.42637, -7.301724, -7.176948, -7.052041, 
    -6.927004, -6.801837, -6.676541, -6.551116, -6.425562, -6.299881, 
    -6.17407, -6.048133, -5.922068, -5.795877, -5.669558, -5.543114, 
    -5.416543, -5.289848, -5.163027, -5.036082, -4.909013, -4.78182, 
    -4.654503, -4.527064, -4.399502, -4.271818, -4.144012, -4.016086, 
    -3.888038, -3.75987, -3.631582, -3.503174, -3.374648, -3.246003, 
    -3.117239, -2.988358, -2.85936, -2.730246, -2.601015, -2.471668, 
    -2.342206, -2.21263, -2.082939, -1.953135, -1.823217, -1.693186, 
    -1.563044, -1.432789, -1.302424, -1.171948, -1.041362, -0.9106658, 
    -0.7798612, -0.648948, -0.5179269, -0.3867985, -0.2555633, -0.1242219, 
    0.007225093, 0.1387772, 0.2704338, 0.4021943, 0.5340581, 0.6660247, 
    0.7980934, 0.9302636, 1.062535, 1.194906, 1.327377, 1.459948, 1.592616, 
    1.725383, 1.858247, 1.991207, 2.124264, 2.257415, 2.390661, 2.524002, 
    2.657435, 2.790962, 2.92458, 3.05829, 3.19209, 3.32598, 3.45996, 
    3.594028, 3.728185, 3.862428, 3.996758, 4.131175, 4.265676, 4.400261, 
    4.534931, 4.669684, 4.804519, 4.939435, 5.074432, 5.20951, 5.344667, 
    5.479903, 5.615216, 5.750607, 5.886075, 6.021617, 6.157236, 6.292928, 
    6.428693, 6.564531, 6.700442, 6.836423, 6.972475, 7.108596, 7.244786, 
    7.381044, 7.51737, 7.653761, 7.790219, 7.926742, 8.063328, 8.199978, 
    8.33669, 8.473463, 8.610298, 8.747192, 8.884146, 9.021158, 9.158228, 
    9.295355, 9.432537, 9.569775, 9.707066, 9.844411, 9.981809, 10.11926, 
    10.25676, 10.39431, 10.53191, 10.66956, 10.80725, 10.94499, 11.08278, 
    11.22061, 11.35849, 11.49641, 11.63437, 11.77237, 11.91042, 12.0485, 
    12.18662, 12.32479, 12.46298, 12.60122, 12.73948, 12.87779, 13.01612, 
    13.15449, 13.2929, 13.43133, 13.56979, 13.70828, 13.8468, 13.98535, 
    14.12392, 14.26252, 14.40114, 14.53979, 14.67846, 14.81715, 14.95586, 
    15.09459, 15.23335, 15.37211, 15.5109, 15.6497, 15.78852, 15.92736, 
    16.0662, 16.20506, 16.34394, 16.48282, 16.62171, 16.76061, 16.89952, 
    17.03844, 17.17736, 17.31629, 17.45523, 17.59417, 17.7331, 17.87205, 
    18.01099, 18.14993, 18.28887, 18.42781, 18.56675, 18.70568, 18.84461, 
    18.98353, 19.12245, 19.26136, 19.40026, 19.53915, 19.67803, 19.8169, 
    19.95576, 20.0946, 20.23344, 20.37225, 20.51105, 20.64984, 20.7886, 
    20.92735, 21.06608, 21.20479, 21.34348, 21.48215, 21.62079, 21.75941, 
    21.898, 22.03657, 22.17511, 22.31363, 22.45211, 22.59057, 22.729, 
    22.8674, 23.00576, 23.14409, 23.28239, 23.42065, 23.55888, 23.69707, 
    23.83523, 23.97334, 24.11142, 24.24946, 24.38745, 24.52541, 24.66332, 
    24.80119, 24.93902, 25.0768, 25.21453, 25.35222, 25.48986, 25.62745, 
    25.765, 25.90249, 26.03993, 26.17732, 26.31466, 26.45194, 26.58917, 
    26.72634, 26.86346, 27.00052, 27.13752, 27.27447, 27.41135, 27.54818, 
    27.68494, 27.82164, 27.95828, 28.09486, 28.23137, 28.36782, 28.5042, 
    28.64051, 28.77676, 28.91294, 29.04905, 29.18509, 29.32106, 29.45696, 
    29.59279, 29.72854, 29.86422, 29.99983, 30.13536, 30.27081, 30.40619, 
    30.54149, 30.67672, 30.81186, 30.94693, 31.08191, 31.21682, 31.35164, 
    31.48638, 31.62103, 31.75561, 31.89009, 32.0245, 32.15881, 32.29304, 
    32.42719, 32.56124, 32.69521, 32.82908, 32.96287, 33.09656, 33.23017, 
    33.36368, 33.4971, 33.63042, 33.76365, 33.89679, 34.02983, 34.16278, 
    34.29562, 34.42838, 34.56103, 34.69358, 34.82604, 34.9584, 35.09065, 
    35.22281, 35.35486, 35.48681, 35.61866, 35.7504, 35.88204, 36.01358, 
    36.145, 36.27633, 36.40755, 36.53866, 36.66966, 36.80056, 36.93135, 
    37.06203, 37.19259, 37.32305, 37.4534, 37.58364, 37.71376, 37.84378, 
    37.97367, 38.10346, 38.23314, 38.36269, 38.49214, 38.62146, 38.75068, 
    38.87977, 39.00875, 39.13762, 39.26636, 39.39499, 39.52349, 39.65188, 
    39.78015, 39.9083, 40.03633, 40.16424, 40.29202, 40.41969, 40.54723, 
    40.67465, 40.80195, 40.92912, 41.05617,
  -16.32838, -16.21387, -16.09923, -15.98443, -15.8695, -15.75442, -15.63919, 
    -15.52382, -15.40831, -15.29266, -15.17686, -15.06091, -14.94483, 
    -14.8286, -14.71223, -14.59571, -14.47905, -14.36225, -14.2453, 
    -14.12821, -14.01098, -13.8936, -13.77608, -13.65843, -13.54062, 
    -13.42268, -13.30459, -13.18636, -13.06799, -12.94947, -12.83082, 
    -12.71202, -12.59308, -12.474, -12.35478, -12.23542, -12.11592, 
    -11.99627, -11.87649, -11.75657, -11.6365, -11.5163, -11.39595, 
    -11.27547, -11.15484, -11.03408, -10.91318, -10.79213, -10.67095, 
    -10.54963, -10.42818, -10.30658, -10.18485, -10.06298, -9.940969, 
    -9.818823, -9.696541, -9.574121, -9.451565, -9.328873, -9.206045, 
    -9.083081, -8.959981, -8.836747, -8.713377, -8.589872, -8.466234, 
    -8.342462, -8.218554, -8.094515, -7.970341, -7.846035, -7.721595, 
    -7.597024, -7.472321, -7.347486, -7.222519, -7.097421, -6.972193, 
    -6.846834, -6.721345, -6.595726, -6.469979, -6.344102, -6.218096, 
    -6.091962, -5.965701, -5.839311, -5.712794, -5.586151, -5.459381, 
    -5.332485, -5.205463, -5.078317, -4.951045, -4.823649, -4.696129, 
    -4.568485, -4.440718, -4.312828, -4.184816, -4.056682, -3.928427, 
    -3.80005, -3.671553, -3.542935, -3.414198, -3.285342, -3.156367, 
    -3.027274, -2.898063, -2.768734, -2.639289, -2.509728, -2.38005, 
    -2.250257, -2.120349, -1.990327, -1.860191, -1.729942, -1.59958, 
    -1.469105, -1.338519, -1.207822, -1.077013, -0.946095, -0.8150671, 
    -0.68393, -0.5526844, -0.4213308, -0.2898699, -0.1583021, -0.02662813, 
    0.1051516, 0.2370363, 0.3690256, 0.5011188, 0.6333154, 0.7656146, 
    0.898016, 1.030519, 1.163123, 1.295827, 1.428631, 1.561533, 1.694535, 
    1.827634, 1.96083, 2.094123, 2.227511, 2.360995, 2.494573, 2.628245, 
    2.762011, 2.895869, 3.029819, 3.16386, 3.297992, 3.432213, 3.566524, 
    3.700923, 3.83541, 3.969984, 4.104645, 4.239391, 4.374222, 4.509138, 
    4.644137, 4.779219, 4.914382, 5.049628, 5.184954, 5.32036, 5.455845, 
    5.591408, 5.72705, 5.862768, 5.998562, 6.134432, 6.270376, 6.406394, 
    6.542486, 6.678649, 6.814885, 6.95119, 7.087567, 7.224012, 7.360526, 
    7.497107, 7.633755, 7.77047, 7.907249, 8.044093, 8.181001, 8.317971, 
    8.455004, 8.592098, 8.729252, 8.866466, 9.003738, 9.141068, 9.278456, 
    9.415899, 9.553398, 9.690952, 9.82856, 9.96622, 10.10393, 10.2417, 
    10.37951, 10.51737, 10.65528, 10.79324, 10.93125, 11.0693, 11.2074, 
    11.34554, 11.48373, 11.62196, 11.76023, 11.89854, 12.03689, 12.17528, 
    12.31371, 12.45217, 12.59067, 12.72921, 12.86778, 13.00639, 13.14503, 
    13.2837, 13.4224, 13.56113, 13.69989, 13.83868, 13.97749, 14.11634, 
    14.25521, 14.3941, 14.53302, 14.67196, 14.81092, 14.9499, 15.0889, 
    15.22793, 15.36697, 15.50603, 15.6451, 15.78419, 15.9233, 16.06242, 
    16.20155, 16.34069, 16.47985, 16.61901, 16.75818, 16.89737, 17.03656, 
    17.17575, 17.31495, 17.45416, 17.59337, 17.73258, 17.8718, 18.01101, 
    18.15022, 18.28944, 18.42865, 18.56786, 18.70707, 18.84627, 18.98546, 
    19.12465, 19.26383, 19.403, 19.54217, 19.68132, 19.82046, 19.95959, 
    20.09871, 20.23781, 20.3769, 20.51597, 20.65503, 20.79407, 20.93308, 
    21.07208, 21.21107, 21.35002, 21.48896, 21.62787, 21.76676, 21.90563, 
    22.04447, 22.18328, 22.32206, 22.46082, 22.59955, 22.73824, 22.87691, 
    23.01554, 23.15414, 23.29271, 23.43124, 23.56973, 23.70819, 23.84661, 
    23.985, 24.12334, 24.26165, 24.39991, 24.53813, 24.67631, 24.81445, 
    24.95254, 25.09058, 25.22858, 25.36653, 25.50444, 25.64229, 25.7801, 
    25.91786, 26.05556, 26.19321, 26.33081, 26.46836, 26.60585, 26.74328, 
    26.88066, 27.01798, 27.15524, 27.29245, 27.42959, 27.56668, 27.7037, 
    27.84066, 27.97756, 28.11439, 28.25116, 28.38787, 28.5245, 28.66107, 
    28.79758, 28.93401, 29.07038, 29.20667, 29.34289, 29.47905, 29.61513, 
    29.75113, 29.88707, 30.02292, 30.15871, 30.29441, 30.43004, 30.56559, 
    30.70107, 30.83646, 30.97177, 31.107, 31.24216, 31.37722, 31.51221, 
    31.64711, 31.78193, 31.91666, 32.05131, 32.18587, 32.32034, 32.45473, 
    32.58902, 32.72323, 32.85735, 32.99137, 33.12531, 33.25916, 33.39291, 
    33.52656, 33.66013, 33.79359, 33.92697, 34.06025, 34.19343, 34.32651, 
    34.4595, 34.59238, 34.72517, 34.85786, 34.99045, 35.12294, 35.25532, 
    35.3876, 35.51978, 35.65186, 35.78383, 35.9157, 36.04746, 36.17912, 
    36.31067, 36.44212, 36.57345, 36.70468, 36.8358, 36.96681, 37.09771, 
    37.2285, 37.35918, 37.48975, 37.62021, 37.75055, 37.88078, 38.0109, 
    38.14091, 38.2708, 38.40057, 38.53023, 38.65977, 38.7892, 38.91851, 
    39.0477, 39.17678, 39.30573, 39.43457, 39.56329, 39.69189, 39.82037, 
    39.94872, 40.07696, 40.20507, 40.33307, 40.46094, 40.58868, 40.71631, 
    40.84381, 40.97119, 41.09844,
  -16.38657, -16.27193, -16.15714, -16.04221, -15.92713, -15.81191, 
    -15.69654, -15.58103, -15.46537, -15.34958, -15.23363, -15.11754, 
    -15.00131, -14.88493, -14.76841, -14.65175, -14.53494, -14.41798, 
    -14.30089, -14.18365, -14.06626, -13.94874, -13.83106, -13.71325, 
    -13.59529, -13.47719, -13.35895, -13.24056, -13.12203, -13.00336, 
    -12.88455, -12.76559, -12.64649, -12.52725, -12.40787, -12.28835, 
    -12.16868, -12.04887, -11.92893, -11.80884, -11.68861, -11.56824, 
    -11.44772, -11.32707, -11.20628, -11.08535, -10.96427, -10.84306, 
    -10.72171, -10.60022, -10.47859, -10.35682, -10.23492, -10.11287, 
    -9.990686, -9.868365, -9.745906, -9.623309, -9.500576, -9.377705, 
    -9.254698, -9.131554, -9.008273, -8.884857, -8.761306, -8.637619, 
    -8.513797, -8.38984, -8.265748, -8.141522, -8.017163, -7.89267, 
    -7.768043, -7.643283, -7.518391, -7.393366, -7.268209, -7.14292, -7.0175, 
    -6.891949, -6.766267, -6.640454, -6.514512, -6.38844, -6.262238, 
    -6.135908, -6.009449, -5.882861, -5.756146, -5.629303, -5.502333, 
    -5.375237, -5.248013, -5.120665, -4.99319, -4.865591, -4.737866, 
    -4.610018, -4.482045, -4.35395, -4.22573, -4.097389, -3.968925, -3.84034, 
    -3.711633, -3.582806, -3.453858, -3.32479, -3.195603, -3.066297, 
    -2.936872, -2.80733, -2.67767, -2.547893, -2.417999, -2.28799, -2.157864, 
    -2.027624, -1.897269, -1.766801, -1.636219, -1.505524, -1.374716, 
    -1.243797, -1.112766, -0.9816245, -0.8503727, -0.7190113, -0.5875407, 
    -0.4559615, -0.3242743, -0.1924797, -0.06057817, 0.07142962, 0.2035431, 
    0.3357617, 0.4680848, 0.6005119, 0.7330423, 0.8656754, 0.9984106, 
    1.131247, 1.264185, 1.397223, 1.53036, 1.663597, 1.796932, 1.930364, 
    2.063894, 2.19752, 2.331242, 2.465059, 2.59897, 2.732975, 2.867074, 
    3.001264, 3.135547, 3.26992, 3.404384, 3.538938, 3.673581, 3.808312, 
    3.943131, 4.078036, 4.213028, 4.348105, 4.483268, 4.618514, 4.753843, 
    4.889256, 5.024749, 5.160325, 5.29598, 5.431715, 5.567529, 5.703421, 
    5.839391, 5.975437, 6.111559, 6.247756, 6.384028, 6.520373, 6.656791, 
    6.793281, 6.929842, 7.066473, 7.203175, 7.339945, 7.476783, 7.613688, 
    7.75066, 7.887698, 8.0248, 8.161966, 8.299196, 8.436488, 8.573842, 
    8.711256, 8.848731, 8.986264, 9.123856, 9.261505, 9.399211, 9.536972, 
    9.674788, 9.812659, 9.950583, 10.08856, 10.22659, 10.36467, 10.50279, 
    10.64097, 10.77919, 10.91747, 11.05579, 11.19415, 11.33256, 11.47101, 
    11.60951, 11.74804, 11.88662, 12.02524, 12.1639, 12.30259, 12.44133, 
    12.5801, 12.7189, 12.85774, 12.99662, 13.13553, 13.27447, 13.41344, 
    13.55244, 13.69147, 13.83053, 13.96962, 14.10873, 14.24787, 14.38703, 
    14.52622, 14.66543, 14.80467, 14.94392, 15.0832, 15.22249, 15.36181, 
    15.50114, 15.64048, 15.77985, 15.91922, 16.05861, 16.19802, 16.33744, 
    16.47686, 16.6163, 16.75575, 16.8952, 17.03467, 17.17414, 17.31361, 
    17.45309, 17.59257, 17.73206, 17.87154, 18.01103, 18.15052, 18.29001, 
    18.42949, 18.56898, 18.70845, 18.84793, 18.98739, 19.12686, 19.26631, 
    19.40576, 19.54519, 19.68462, 19.82403, 19.96343, 20.10283, 20.2422, 
    20.38156, 20.5209, 20.66023, 20.79954, 20.93884, 21.07811, 21.21736, 
    21.35659, 21.4958, 21.63498, 21.77414, 21.91328, 22.05239, 22.19147, 
    22.33052, 22.46955, 22.60855, 22.74751, 22.88645, 23.02535, 23.16422, 
    23.30306, 23.44186, 23.58062, 23.71935, 23.85804, 23.99669, 24.1353, 
    24.27387, 24.41241, 24.55089, 24.68934, 24.82774, 24.9661, 25.10441, 
    25.24267, 25.38089, 25.51906, 25.65718, 25.79525, 25.93327, 26.07124, 
    26.20915, 26.34702, 26.48482, 26.62258, 26.76027, 26.89791, 27.0355, 
    27.17302, 27.31048, 27.44789, 27.58523, 27.72252, 27.85974, 27.99689, 
    28.13398, 28.27101, 28.40797, 28.54487, 28.68169, 28.81845, 28.95514, 
    29.09176, 29.22832, 29.36479, 29.5012, 29.63753, 29.77379, 29.90998, 
    30.04609, 30.18212, 30.31808, 30.45396, 30.58976, 30.72548, 30.86113, 
    30.99669, 31.13217, 31.26757, 31.40289, 31.53812, 31.67327, 31.80833, 
    31.94331, 32.0782, 32.21301, 32.34772, 32.48235, 32.61689, 32.75134, 
    32.8857, 33.01997, 33.15414, 33.28823, 33.42222, 33.55611, 33.68992, 
    33.82362, 33.95723, 34.09075, 34.22417, 34.35749, 34.49071, 34.62383, 
    34.75685, 34.88977, 35.02259, 35.15531, 35.28793, 35.42044, 35.55285, 
    35.68516, 35.81736, 35.94946, 36.08145, 36.21333, 36.34511, 36.47678, 
    36.60835, 36.7398, 36.87114, 37.00238, 37.1335, 37.26451, 37.39542, 
    37.52621, 37.65688, 37.78745, 37.9179, 38.04823, 38.17846, 38.30856, 
    38.43855, 38.56843, 38.69819, 38.82783, 38.95735, 39.08676, 39.21605, 
    39.34521, 39.47426, 39.60319, 39.732, 39.86069, 39.98925, 40.1177, 
    40.24602, 40.37422, 40.5023, 40.63025, 40.75808, 40.88578, 41.01336, 
    41.14082,
  -16.44489, -16.33011, -16.21519, -16.10011, -15.98489, -15.86953, 
    -15.75402, -15.63836, -15.52256, -15.40662, -15.29053, -15.1743, 
    -15.05792, -14.94139, -14.82472, -14.70791, -14.59095, -14.47385, 
    -14.3566, -14.23921, -14.12167, -14.00399, -13.88617, -13.7682, 
    -13.65009, -13.53184, -13.41344, -13.29489, -13.17621, -13.05738, 
    -12.93841, -12.81929, -12.70003, -12.58063, -12.46109, -12.3414, 
    -12.22157, -12.1016, -11.98149, -11.86123, -11.74084, -11.6203, 
    -11.49962, -11.3788, -11.25784, -11.13674, -11.0155, -10.89412, 
    -10.77259, -10.65093, -10.52913, -10.40719, -10.28511, -10.16289, 
    -10.04053, -9.918032, -9.795396, -9.672622, -9.54971, -9.426661, 
    -9.303473, -9.180149, -9.056688, -8.933091, -8.809357, -8.685487, 
    -8.561481, -8.43734, -8.313064, -8.188652, -8.064106, -7.939425, 
    -7.81461, -7.689662, -7.56458, -7.439366, -7.314018, -7.188538, 
    -7.062926, -6.937182, -6.811306, -6.6853, -6.559163, -6.432895, 
    -6.306498, -6.17997, -6.053313, -5.926528, -5.799613, -5.672571, 
    -5.545401, -5.418103, -5.290678, -5.163127, -5.035449, -4.907646, 
    -4.779717, -4.651663, -4.523485, -4.395183, -4.266757, -4.138207, 
    -4.009535, -3.88074, -3.751824, -3.622786, -3.493627, -3.364347, 
    -3.234947, -3.105428, -2.97579, -2.846033, -2.716157, -2.586164, 
    -2.456054, -2.325827, -2.195484, -2.065026, -1.934452, -1.803764, 
    -1.672961, -1.542045, -1.411016, -1.279874, -1.14862, -1.017255, 
    -0.885779, -0.7541926, -0.6224965, -0.4906912, -0.3587772, -0.2267552, 
    -0.09462567, 0.03761074, 0.1699535, 0.3024019, 0.4349555, 0.5676136, 
    0.7003757, 0.833241, 0.9662091, 1.099279, 1.232451, 1.365723, 1.499096, 
    1.632568, 1.76614, 1.899809, 2.033576, 2.16744, 2.301401, 2.435457, 
    2.569608, 2.703854, 2.838193, 2.972625, 3.10715, 3.241766, 3.376473, 
    3.51127, 3.646157, 3.781133, 3.916197, 4.051348, 4.186586, 4.32191, 
    4.45732, 4.592814, 4.728392, 4.864052, 4.999796, 5.135621, 5.271526, 
    5.407512, 5.543578, 5.679721, 5.815943, 5.952242, 6.088617, 6.225068, 
    6.361593, 6.498193, 6.634866, 6.771611, 6.908428, 7.045316, 7.182274, 
    7.319301, 7.456397, 7.59356, 7.73079, 7.868086, 8.005447, 8.142874, 
    8.280363, 8.417915, 8.55553, 8.693206, 8.830941, 8.968737, 9.10659, 
    9.244502, 9.382471, 9.520495, 9.658575, 9.79671, 9.934897, 10.07314, 
    10.21143, 10.34977, 10.48817, 10.62661, 10.7651, 10.90364, 11.04222, 
    11.18086, 11.31953, 11.45825, 11.59701, 11.73582, 11.87467, 12.01355, 
    12.15248, 12.29144, 12.43045, 12.56949, 12.70856, 12.84767, 12.98682, 
    13.126, 13.26521, 13.40445, 13.54372, 13.68302, 13.82236, 13.96171, 
    14.1011, 14.24051, 14.37995, 14.51941, 14.65889, 14.7984, 14.93793, 
    15.07747, 15.21704, 15.35663, 15.49623, 15.63585, 15.77549, 15.91514, 
    16.0548, 16.19448, 16.33417, 16.47387, 16.61358, 16.7533, 16.89303, 
    17.03277, 17.17251, 17.31226, 17.45201, 17.59177, 17.73153, 17.87129, 
    18.01105, 18.15082, 18.29058, 18.43034, 18.57009, 18.70984, 18.84959, 
    18.98933, 19.12907, 19.2688, 19.40852, 19.54823, 19.68793, 19.82761, 
    19.96729, 20.10695, 20.2466, 20.38624, 20.52585, 20.66545, 20.80504, 
    20.9446, 21.08415, 21.22367, 21.36317, 21.50266, 21.64211, 21.78154, 
    21.92095, 22.06033, 22.19969, 22.33901, 22.47831, 22.61758, 22.75681, 
    22.89602, 23.03519, 23.17433, 23.31344, 23.45251, 23.59154, 23.73054, 
    23.8695, 24.00842, 24.1473, 24.28614, 24.42494, 24.56369, 24.70241, 
    24.84108, 24.9797, 25.11828, 25.25681, 25.39529, 25.53373, 25.67211, 
    25.81045, 25.94873, 26.08697, 26.22515, 26.36327, 26.50134, 26.63936, 
    26.77732, 26.91522, 27.05306, 27.19085, 27.32858, 27.46624, 27.60385, 
    27.74139, 27.87887, 28.01628, 28.15364, 28.29092, 28.42814, 28.56529, 
    28.70238, 28.8394, 28.97634, 29.11322, 29.25002, 29.38676, 29.52342, 
    29.66001, 29.79652, 29.93296, 30.06932, 30.20561, 30.34182, 30.47795, 
    30.614, 30.74998, 30.88587, 31.02168, 31.15741, 31.29306, 31.42863, 
    31.56411, 31.6995, 31.83481, 31.97004, 32.10518, 32.24022, 32.37519, 
    32.51006, 32.64484, 32.77953, 32.91413, 33.04865, 33.18306, 33.31739, 
    33.45162, 33.58575, 33.7198, 33.85374, 33.98759, 34.12134, 34.255, 
    34.38855, 34.52201, 34.65536, 34.78862, 34.92178, 35.05483, 35.18778, 
    35.32063, 35.45338, 35.58602, 35.71856, 35.85099, 35.98331, 36.11553, 
    36.24765, 36.37965, 36.51155, 36.64334, 36.77501, 36.90659, 37.03804, 
    37.16939, 37.30062, 37.43175, 37.56276, 37.69366, 37.82444, 37.95512, 
    38.08567, 38.21611, 38.34644, 38.47664, 38.60674, 38.73671, 38.86657, 
    38.9963, 39.12592, 39.25542, 39.3848, 39.51406, 39.6432, 39.77222, 
    39.90112, 40.0299, 40.15855, 40.28708, 40.41549, 40.54377, 40.67193, 
    40.79996, 40.92787, 41.05565, 41.18331,
  -16.50335, -16.38842, -16.27336, -16.15814, -16.04278, -15.92728, 
    -15.81163, -15.69583, -15.57988, -15.46379, -15.34756, -15.23118, 
    -15.11465, -14.99798, -14.88117, -14.7642, -14.6471, -14.52984, 
    -14.41245, -14.2949, -14.17722, -14.05938, -13.94141, -13.82328, 
    -13.70502, -13.58661, -13.46805, -13.34935, -13.23051, -13.11152, 
    -12.99239, -12.87312, -12.7537, -12.63414, -12.51443, -12.39458, 
    -12.27459, -12.15446, -12.03418, -11.91376, -11.7932, -11.67249, 
    -11.55165, -11.43066, -11.30953, -11.18826, -11.06685, -10.9453, 
    -10.8236, -10.70177, -10.57979, -10.45768, -10.33543, -10.21303, 
    -10.0905, -9.967823, -9.84501, -9.722058, -9.598969, -9.47574, -9.352373, 
    -9.228869, -9.105227, -8.981447, -8.857532, -8.733478, -8.609288, 
    -8.484962, -8.3605, -8.235903, -8.11117, -7.986302, -7.8613, -7.736163, 
    -7.610891, -7.485487, -7.359948, -7.234276, -7.108472, -6.982535, 
    -6.856465, -6.730265, -6.603932, -6.477468, -6.350874, -6.22415, 
    -6.097295, -5.970311, -5.843197, -5.715955, -5.588584, -5.461085, 
    -5.333458, -5.205704, -5.077823, -4.949815, -4.821682, -4.693423, 
    -4.565038, -4.436529, -4.307895, -4.179137, -4.050256, -3.921252, 
    -3.792125, -3.662876, -3.533506, -3.404014, -3.274401, -3.144668, 
    -3.014815, -2.884843, -2.754752, -2.624543, -2.494216, -2.363772, 
    -2.23321, -2.102533, -1.971739, -1.840831, -1.709807, -1.578669, 
    -1.447418, -1.316054, -1.184576, -1.052987, -0.9212863, -0.7894745, 
    -0.6575524, -0.5255204, -0.3933792, -0.2611293, -0.1287713, 0.00369428, 
    0.1362668, 0.2689456, 0.4017302, 0.5346199, 0.6676142, 0.8007123, 
    0.9339138, 1.067218, 1.200624, 1.334132, 1.46774, 1.601449, 1.735257, 
    1.869164, 2.00317, 2.137272, 2.271472, 2.405768, 2.54016, 2.674646, 
    2.809227, 2.943901, 3.078668, 3.213528, 3.348479, 3.48352, 3.618652, 
    3.753873, 3.889183, 4.02458, 4.160065, 4.295637, 4.431294, 4.567037, 
    4.702863, 4.838774, 4.974767, 5.110842, 5.246999, 5.383236, 5.519553, 
    5.65595, 5.792424, 5.928977, 6.065606, 6.202311, 6.339091, 6.475945, 
    6.612874, 6.749875, 6.886949, 7.024094, 7.161309, 7.298594, 7.435947, 
    7.57337, 7.710859, 7.848414, 7.986036, 8.123722, 8.261473, 8.399285, 
    8.537162, 8.675098, 8.813097, 8.951155, 9.089272, 9.227447, 9.365679, 
    9.503967, 9.642311, 9.78071, 9.919164, 10.05767, 10.19623, 10.33484, 
    10.4735, 10.61221, 10.75096, 10.88977, 11.02862, 11.16752, 11.30647, 
    11.44545, 11.58449, 11.72356, 11.86267, 12.00183, 12.14103, 12.28026, 
    12.41953, 12.55885, 12.69819, 12.83757, 12.97699, 13.11644, 13.25592, 
    13.39543, 13.53498, 13.67455, 13.81416, 13.95379, 14.09344, 14.23313, 
    14.37284, 14.51257, 14.65233, 14.79211, 14.93191, 15.07173, 15.21157, 
    15.35143, 15.49131, 15.6312, 15.77111, 15.91104, 16.05098, 16.19093, 
    16.33089, 16.47087, 16.61086, 16.75085, 16.89086, 17.03087, 17.17089, 
    17.31091, 17.45094, 17.59097, 17.731, 17.87104, 18.01108, 18.15111, 
    18.29115, 18.43118, 18.57121, 18.71124, 18.85126, 18.99128, 19.13129, 
    19.27129, 19.41129, 19.55127, 19.69125, 19.83121, 19.97116, 20.1111, 
    20.25102, 20.39093, 20.53082, 20.67069, 20.81055, 20.95039, 21.09021, 
    21.23, 21.36978, 21.50953, 21.64926, 21.78897, 21.92865, 22.0683, 
    22.20793, 22.34753, 22.4871, 22.62664, 22.76615, 22.90562, 23.04507, 
    23.18448, 23.32385, 23.46319, 23.6025, 23.74177, 23.88099, 24.02018, 
    24.15933, 24.29844, 24.43751, 24.57654, 24.71552, 24.85445, 24.99335, 
    25.13219, 25.27099, 25.40974, 25.54844, 25.68709, 25.82569, 25.96424, 
    26.10274, 26.24119, 26.37958, 26.51791, 26.65619, 26.79441, 26.93258, 
    27.07069, 27.20874, 27.34673, 27.48465, 27.62252, 27.76032, 27.89806, 
    28.03574, 28.17335, 28.31089, 28.44837, 28.58578, 28.72313, 28.8604, 
    28.99761, 29.13474, 29.2718, 29.40879, 29.54571, 29.68255, 29.81932, 
    29.95601, 30.09263, 30.22917, 30.36563, 30.50202, 30.63832, 30.77454, 
    30.91069, 31.04675, 31.18273, 31.31863, 31.45444, 31.59017, 31.72581, 
    31.86137, 31.99684, 32.13223, 32.26752, 32.40273, 32.53785, 32.67287, 
    32.80781, 32.94266, 33.07741, 33.21207, 33.34663, 33.48111, 33.61548, 
    33.74976, 33.88395, 34.01804, 34.15202, 34.28592, 34.41971, 34.5534, 
    34.68699, 34.82048, 34.95388, 35.08716, 35.22035, 35.35343, 35.48641, 
    35.61928, 35.75205, 35.88471, 36.01727, 36.14972, 36.28205, 36.41429, 
    36.54641, 36.67843, 36.81033, 36.94213, 37.07381, 37.20538, 37.33684, 
    37.46819, 37.59942, 37.73054, 37.86155, 37.99244, 38.12321, 38.25387, 
    38.38441, 38.51484, 38.64515, 38.77534, 38.90541, 39.03536, 39.1652, 
    39.29491, 39.42451, 39.55398, 39.68333, 39.81256, 39.94167, 40.07065, 
    40.19951, 40.32825, 40.45686, 40.58535, 40.71372, 40.84196, 40.97007, 
    41.09806, 41.22592,
  -16.56193, -16.44687, -16.33166, -16.2163, -16.1008, -15.98516, -15.86936, 
    -15.75342, -15.63733, -15.5211, -15.40472, -15.28819, -15.17152, 
    -15.0547, -14.93774, -14.82063, -14.70337, -14.58597, -14.46842, 
    -14.35073, -14.23289, -14.1149, -13.99677, -13.87849, -13.76007, 
    -13.64151, -13.5228, -13.40394, -13.28494, -13.16579, -13.0465, 
    -12.92707, -12.80749, -12.68777, -12.5679, -12.44789, -12.32774, 
    -12.20744, -12.087, -11.96641, -11.84569, -11.72482, -11.6038, -11.48265, 
    -11.36135, -11.23991, -11.11833, -10.9966, -10.87474, -10.75273, 
    -10.63059, -10.5083, -10.38587, -10.2633, -10.14059, -10.01774, -9.89475, 
    -9.771621, -9.648352, -9.524944, -9.401398, -9.277713, -9.15389, 
    -9.029928, -8.905829, -8.781592, -8.657219, -8.532708, -8.408061, 
    -8.283278, -8.158358, -8.033301, -7.908111, -7.782784, -7.657323, 
    -7.531728, -7.405998, -7.280135, -7.154138, -7.028008, -6.901744, 
    -6.775349, -6.648821, -6.522161, -6.39537, -6.268448, -6.141395, 
    -6.014212, -5.886899, -5.759456, -5.631884, -5.504183, -5.376354, 
    -5.248397, -5.120312, -4.9921, -4.863761, -4.735296, -4.606705, 
    -4.477988, -4.349147, -4.220181, -4.09109, -3.961876, -3.832538, 
    -3.703078, -3.573495, -3.443791, -3.313965, -3.184018, -3.05395, 
    -2.923763, -2.793456, -2.66303, -2.532485, -2.401823, -2.271043, 
    -2.140146, -2.009132, -1.878003, -1.746758, -1.615398, -1.483924, 
    -1.352336, -1.220635, -1.088821, -0.9568955, -0.8248578, -0.6927092, 
    -0.5604501, -0.428081, -0.2956027, -0.1630156, -0.03032041, 0.1024824, 
    0.2353921, 0.3684082, 0.5015301, 0.634757, 0.7680886, 0.9015241, 
    1.035063, 1.168704, 1.302448, 1.436292, 1.570238, 1.704284, 1.838429, 
    1.972673, 2.107015, 2.241455, 2.375991, 2.510624, 2.645352, 2.780174, 
    2.915092, 3.050102, 3.185205, 3.3204, 3.455687, 3.591064, 3.726531, 
    3.862087, 3.997732, 4.133464, 4.269284, 4.40519, 4.541182, 4.677258, 
    4.813418, 4.949662, 5.085989, 5.222397, 5.358886, 5.495456, 5.632105, 
    5.768834, 5.90564, 6.042523, 6.179483, 6.316519, 6.45363, 6.590815, 
    6.728073, 6.865403, 7.002806, 7.140279, 7.277822, 7.415436, 7.553117, 
    7.690866, 7.828682, 7.966564, 8.104511, 8.242523, 8.380598, 8.518736, 
    8.656936, 8.795197, 8.933518, 9.071898, 9.210338, 9.348834, 9.487388, 
    9.625997, 9.764662, 9.90338, 10.04215, 10.18098, 10.31985, 10.45878, 
    10.59776, 10.73678, 10.87586, 11.01498, 11.15414, 11.29336, 11.43261, 
    11.57192, 11.71126, 11.85065, 11.99007, 12.12954, 12.26904, 12.40859, 
    12.54817, 12.68779, 12.82744, 12.96713, 13.10685, 13.2466, 13.38639, 
    13.52621, 13.66605, 13.80593, 13.94583, 14.08577, 14.22572, 14.36571, 
    14.50571, 14.64575, 14.7858, 14.92587, 15.06597, 15.20609, 15.34622, 
    15.48637, 15.62654, 15.76673, 15.90693, 16.04714, 16.18737, 16.32761, 
    16.46786, 16.60812, 16.74839, 16.88867, 17.02896, 17.16925, 17.30955, 
    17.44986, 17.59016, 17.73047, 17.87078, 18.0111, 18.15141, 18.29172, 
    18.43203, 18.57234, 18.71264, 18.85294, 18.99323, 19.13352, 19.2738, 
    19.41407, 19.55433, 19.69458, 19.83481, 19.97504, 20.11525, 20.25545, 
    20.39563, 20.5358, 20.67595, 20.81608, 20.95619, 21.09628, 21.23636, 
    21.37641, 21.51644, 21.65644, 21.79642, 21.93637, 22.0763, 22.2162, 
    22.35607, 22.49591, 22.63573, 22.77551, 22.91525, 23.05497, 23.19465, 
    23.3343, 23.47391, 23.61349, 23.75303, 23.89253, 24.03199, 24.17141, 
    24.31079, 24.45012, 24.58942, 24.72867, 24.86787, 25.00703, 25.14615, 
    25.28521, 25.42423, 25.5632, 25.70212, 25.84099, 25.9798, 26.11857, 
    26.25728, 26.39593, 26.53453, 26.67308, 26.81157, 26.95, 27.08837, 
    27.22668, 27.36493, 27.50312, 27.64125, 27.77931, 27.91731, 28.05525, 
    28.19312, 28.33093, 28.46867, 28.60634, 28.74394, 28.88147, 29.01893, 
    29.15632, 29.29364, 29.43089, 29.56806, 29.70516, 29.84219, 29.97913, 
    30.116, 30.2528, 30.38951, 30.52615, 30.66271, 30.79919, 30.93558, 
    31.0719, 31.20813, 31.34427, 31.48034, 31.61631, 31.75221, 31.88801, 
    32.02373, 32.15936, 32.2949, 32.43036, 32.56572, 32.70099, 32.83617, 
    32.97126, 33.10625, 33.24116, 33.37597, 33.51068, 33.6453, 33.77982, 
    33.91424, 34.04857, 34.1828, 34.31693, 34.45096, 34.58488, 34.71872, 
    34.85244, 34.98607, 35.11959, 35.25301, 35.38633, 35.51954, 35.65264, 
    35.78564, 35.91853, 36.05132, 36.18399, 36.31657, 36.44903, 36.58138, 
    36.71362, 36.84575, 36.97777, 37.10968, 37.24147, 37.37316, 37.50473, 
    37.63618, 37.76753, 37.89875, 38.02987, 38.16086, 38.29174, 38.4225, 
    38.55314, 38.68367, 38.81408, 38.94436, 39.07453, 39.20458, 39.33451, 
    39.46432, 39.594, 39.72356, 39.853, 39.98232, 40.11152, 40.24059, 
    40.36954, 40.49836, 40.62706, 40.75563, 40.88407, 41.01239, 41.14058, 
    41.26865,
  -16.62064, -16.50544, -16.39009, -16.2746, -16.15895, -16.04316, -15.92723, 
    -15.81114, -15.69491, -15.57853, -15.46201, -15.34534, -15.22852, 
    -15.11155, -14.99444, -14.87718, -14.75977, -14.64222, -14.52452, 
    -14.40668, -14.28869, -14.17055, -14.05227, -13.93384, -13.81526, 
    -13.69654, -13.57767, -13.45866, -13.3395, -13.2202, -13.10075, 
    -12.98115, -12.86141, -12.74153, -12.6215, -12.50133, -12.38101, 
    -12.26055, -12.13995, -12.0192, -11.8983, -11.77727, -11.65609, 
    -11.53476, -11.4133, -11.29169, -11.16993, -11.04804, -10.926, -10.80383, 
    -10.68151, -10.55904, -10.43644, -10.31369, -10.19081, -10.06778, 
    -9.944615, -9.821308, -9.697862, -9.574274, -9.450548, -9.326682, 
    -9.202678, -9.078534, -8.954252, -8.829832, -8.705274, -8.580578, 
    -8.455745, -8.330774, -8.205667, -8.080424, -7.955044, -7.829529, 
    -7.703878, -7.578092, -7.45217, -7.326115, -7.199925, -7.073601, 
    -6.947144, -6.820553, -6.69383, -6.566973, -6.439985, -6.312865, 
    -6.185614, -6.058231, -5.930718, -5.803075, -5.675302, -5.547399, 
    -5.419367, -5.291206, -5.162917, -5.0345, -4.905956, -4.777285, 
    -4.648487, -4.519562, -4.390512, -4.261337, -4.132037, -4.002613, 
    -3.873064, -3.743392, -3.613597, -3.483679, -3.353639, -3.223478, 
    -3.093195, -2.962792, -2.832268, -2.701625, -2.570863, -2.439982, 
    -2.308983, -2.177866, -2.046632, -1.915281, -1.783814, -1.652232, 
    -1.520535, -1.388723, -1.256798, -1.124759, -0.9926071, -0.8603431, 
    -0.7279674, -0.5954806, -0.4628833, -0.3301761, -0.1973594, -0.06443399, 
    0.0685996, 0.2017408, 0.334989, 0.4683435, 0.6018038, 0.7353693, 
    0.8690392, 1.002813, 1.13669, 1.27067, 1.404752, 1.538935, 1.673219, 
    1.807603, 1.942086, 2.076668, 2.211348, 2.346125, 2.481, 2.61597, 
    2.751035, 2.886196, 3.02145, 3.156798, 3.292238, 3.42777, 3.563393, 
    3.699107, 3.83491, 3.970803, 4.106783, 4.242852, 4.379007, 4.515248, 
    4.651575, 4.787986, 4.924481, 5.061059, 5.19772, 5.334462, 5.471285, 
    5.608189, 5.745171, 5.882232, 6.019371, 6.156587, 6.293878, 6.431245, 
    6.568687, 6.706203, 6.843792, 6.981452, 7.119185, 7.256988, 7.39486, 
    7.532802, 7.670811, 7.808888, 7.947031, 8.08524, 8.223515, 8.361853, 
    8.500254, 8.638717, 8.777241, 8.915827, 9.054471, 9.193175, 9.331937, 
    9.470757, 9.609632, 9.748562, 9.887547, 10.02659, 10.16568, 10.30482, 
    10.44402, 10.58326, 10.72256, 10.8619, 11.00129, 11.14073, 11.28021, 
    11.41974, 11.55931, 11.69892, 11.83858, 11.97828, 12.11801, 12.25779, 
    12.39761, 12.53746, 12.67735, 12.81728, 12.95724, 13.09723, 13.23726, 
    13.37732, 13.51741, 13.65753, 13.79768, 13.93786, 14.07806, 14.21829, 
    14.35855, 14.49883, 14.63914, 14.77947, 14.91982, 15.06019, 15.20058, 
    15.34099, 15.48142, 15.62186, 15.76233, 15.9028, 16.04329, 16.1838, 
    16.32431, 16.46484, 16.60538, 16.74593, 16.88648, 17.02704, 17.16761, 
    17.30819, 17.44877, 17.58935, 17.72994, 17.87053, 18.01112, 18.15171, 
    18.2923, 18.43288, 18.57347, 18.71405, 18.85462, 18.99519, 19.13575, 
    19.27631, 19.41685, 19.55739, 19.69792, 19.83843, 19.97893, 20.11942, 
    20.25989, 20.40035, 20.54079, 20.68122, 20.82163, 20.96202, 21.10238, 
    21.24273, 21.38306, 21.52336, 21.66364, 21.80389, 21.94412, 22.08432, 
    22.22449, 22.36464, 22.50476, 22.64484, 22.78489, 22.92492, 23.06491, 
    23.20486, 23.34478, 23.48466, 23.62451, 23.76432, 23.90409, 24.04383, 
    24.18352, 24.32317, 24.46277, 24.60234, 24.74186, 24.88133, 25.02076, 
    25.16015, 25.29948, 25.43877, 25.578, 25.71719, 25.85633, 25.99541, 
    26.13444, 26.27342, 26.41234, 26.55121, 26.69002, 26.82877, 26.96746, 
    27.1061, 27.24467, 27.38319, 27.52164, 27.66003, 27.79836, 27.93663, 
    28.07483, 28.21296, 28.35102, 28.48902, 28.62695, 28.76481, 28.90261, 
    29.04033, 29.17798, 29.31556, 29.45306, 29.59049, 29.72784, 29.86512, 
    30.00233, 30.13945, 30.2765, 30.41347, 30.55036, 30.68717, 30.8239, 
    30.96055, 31.09712, 31.2336, 31.37, 31.50631, 31.64254, 31.77868, 
    31.91473, 32.0507, 32.18658, 32.32237, 32.45807, 32.59367, 32.72919, 
    32.86462, 32.99995, 33.13519, 33.27034, 33.40539, 33.54034, 33.6752, 
    33.80996, 33.94463, 34.07919, 34.21366, 34.34803, 34.4823, 34.61647, 
    34.75053, 34.88449, 35.01836, 35.15211, 35.28577, 35.41932, 35.55276, 
    35.6861, 35.81933, 35.95245, 36.08547, 36.21838, 36.35118, 36.48386, 
    36.61644, 36.74891, 36.88127, 37.01352, 37.14565, 37.27768, 37.40958, 
    37.54137, 37.67305, 37.80462, 37.93607, 38.0674, 38.19862, 38.32971, 
    38.46069, 38.59156, 38.7223, 38.85292, 38.98343, 39.11381, 39.24408, 
    39.37422, 39.50424, 39.63414, 39.76391, 39.89357, 40.02309, 40.1525, 
    40.28178, 40.41093, 40.53996, 40.66887, 40.79765, 40.9263, 41.05482, 
    41.18322, 41.31149,
  -16.67948, -16.56414, -16.44865, -16.33302, -16.21723, -16.1013, -15.98522, 
    -15.869, -15.75262, -15.6361, -15.51943, -15.40261, -15.28565, -15.16853, 
    -15.05127, -14.93386, -14.81631, -14.69861, -14.58076, -14.46276, 
    -14.34462, -14.22633, -14.10789, -13.98931, -13.87058, -13.7517, 
    -13.63268, -13.51351, -13.39419, -13.27473, -13.15512, -13.03537, 
    -12.91547, -12.79542, -12.67523, -12.5549, -12.43442, -12.31379, 
    -12.19302, -12.07211, -11.95105, -11.82984, -11.7085, -11.587, -11.46537, 
    -11.34359, -11.22167, -11.0996, -10.9774, -10.85504, -10.73255, 
    -10.60992, -10.48714, -10.36422, -10.24116, -10.11795, -9.994609, 
    -9.871123, -9.747498, -9.623731, -9.499825, -9.375777, -9.251591, 
    -9.127265, -9.0028, -8.878196, -8.753453, -8.628572, -8.503553, 
    -8.378396, -8.253101, -8.12767, -8.002102, -7.876397, -7.750556, 
    -7.624578, -7.498465, -7.372217, -7.245834, -7.119316, -6.992664, 
    -6.865878, -6.738959, -6.611906, -6.48472, -6.357402, -6.229952, 
    -6.10237, -5.974657, -5.846812, -5.718837, -5.590732, -5.462497, 
    -5.334133, -5.205639, -5.077017, -4.948267, -4.819389, -4.690383, 
    -4.561251, -4.431993, -4.302608, -4.173098, -4.043462, -3.913702, 
    -3.783818, -3.65381, -3.523679, -3.393425, -3.263049, -3.13255, 
    -3.001931, -2.87119, -2.74033, -2.609349, -2.478249, -2.34703, -2.215693, 
    -2.084238, -1.952666, -1.820977, -1.689172, -1.557251, -1.425215, 
    -1.293064, -1.1608, -1.028422, -0.895931, -0.7633278, -0.6306129, 
    -0.4977867, -0.36485, -0.2318033, -0.09864712, 0.03461784, 0.167991, 
    0.3014718, 0.4350595, 0.5687537, 0.7025536, 0.8364587, 0.9704683, 
    1.104582, 1.238798, 1.373118, 1.507539, 1.642061, 1.776685, 1.911408, 
    2.04623, 2.181151, 2.31617, 2.451287, 2.5865, 2.721809, 2.857213, 
    2.992712, 3.128305, 3.26399, 3.399769, 3.535639, 3.671599, 3.807651, 
    3.943791, 4.080021, 4.216339, 4.352744, 4.489236, 4.625813, 4.762476, 
    4.899223, 5.036054, 5.172968, 5.309964, 5.447041, 5.584198, 5.721436, 
    5.858752, 5.996147, 6.133619, 6.271168, 6.408792, 6.546492, 6.684266, 
    6.822113, 6.960033, 7.098025, 7.236088, 7.374221, 7.512424, 7.650694, 
    7.789033, 7.927438, 8.06591, 8.204447, 8.343048, 8.481712, 8.62044, 
    8.75923, 8.89808, 9.03699, 9.17596, 9.314987, 9.454073, 9.593215, 
    9.732412, 9.871665, 10.01097, 10.15033, 10.28974, 10.42921, 10.56872, 
    10.70829, 10.8479, 10.98756, 11.12726, 11.26702, 11.40682, 11.54666, 
    11.68654, 11.82647, 11.96644, 12.10645, 12.2465, 12.38659, 12.52672, 
    12.66688, 12.80708, 12.94731, 13.08758, 13.22788, 13.36821, 13.50858, 
    13.64898, 13.7894, 13.92985, 14.07033, 14.21084, 14.35137, 14.49193, 
    14.63251, 14.77312, 14.91374, 15.05439, 15.19506, 15.33575, 15.47645, 
    15.61717, 15.75791, 15.89866, 16.03943, 16.18021, 16.321, 16.46181, 
    16.60262, 16.74345, 16.88428, 17.02512, 17.16597, 17.30682, 17.44768, 
    17.58854, 17.72941, 17.87027, 18.01114, 18.15201, 18.29288, 18.43374, 
    18.5746, 18.71546, 18.85631, 18.99716, 19.13799, 19.27883, 19.41965, 
    19.56046, 19.70127, 19.84206, 19.98284, 20.1236, 20.26435, 20.40509, 
    20.54581, 20.68651, 20.82719, 20.96786, 21.1085, 21.24912, 21.38972, 
    21.5303, 21.67086, 21.81139, 21.95189, 22.09237, 22.23281, 22.37324, 
    22.51363, 22.65399, 22.79431, 22.93461, 23.07487, 23.2151, 23.3553, 
    23.49545, 23.63557, 23.77566, 23.9157, 24.0557, 24.19567, 24.33559, 
    24.47547, 24.6153, 24.75509, 24.89484, 25.03454, 25.17419, 25.3138, 
    25.45335, 25.59286, 25.73231, 25.87172, 26.01107, 26.15037, 26.28961, 
    26.4288, 26.56793, 26.70701, 26.84603, 26.98499, 27.12389, 27.26273, 
    27.40151, 27.54023, 27.67888, 27.81747, 27.956, 28.09446, 28.23285, 
    28.37118, 28.50944, 28.64763, 28.78576, 28.92381, 29.06179, 29.1997, 
    29.33753, 29.47529, 29.61298, 29.7506, 29.88813, 30.02559, 30.16298, 
    30.30028, 30.4375, 30.57465, 30.71171, 30.8487, 30.9856, 31.12241, 
    31.25915, 31.3958, 31.53236, 31.66884, 31.80523, 31.94153, 32.07775, 
    32.21387, 32.34991, 32.48586, 32.62172, 32.75748, 32.89315, 33.02873, 
    33.16421, 33.2996, 33.43489, 33.57009, 33.70519, 33.8402, 33.9751, 
    34.10991, 34.24462, 34.37922, 34.51373, 34.64814, 34.78244, 34.91664, 
    35.05074, 35.18473, 35.31862, 35.4524, 35.58608, 35.71965, 35.85312, 
    35.98647, 36.11972, 36.25286, 36.38589, 36.51881, 36.65162, 36.78431, 
    36.9169, 37.04937, 37.18173, 37.31398, 37.44611, 37.57812, 37.71003, 
    37.84182, 37.97349, 38.10504, 38.23648, 38.36779, 38.499, 38.63008, 
    38.76104, 38.89188, 39.0226, 39.1532, 39.28368, 39.41404, 39.54427, 
    39.67439, 39.80437, 39.93424, 40.06398, 40.19359, 40.32308, 40.45245, 
    40.58169, 40.7108, 40.83978, 40.96864, 41.09737, 41.22598, 41.35445,
  -16.73845, -16.62298, -16.50735, -16.39157, -16.27565, -16.15957, 
    -16.04335, -15.92698, -15.81046, -15.6938, -15.57698, -15.46002, 
    -15.34291, -15.22565, -15.10824, -14.99068, -14.87298, -14.75513, 
    -14.63712, -14.51898, -14.40068, -14.28224, -14.16365, -14.04491, 
    -13.92602, -13.80699, -13.68781, -13.56849, -13.44901, -13.32939, 
    -13.20962, -13.08971, -12.96965, -12.84945, -12.72909, -12.6086, 
    -12.48795, -12.36716, -12.24623, -12.12515, -12.00392, -11.88255, 
    -11.76104, -11.63938, -11.51757, -11.39563, -11.27353, -11.1513, 
    -11.02892, -10.90639, -10.78373, -10.66092, -10.53796, -10.41487, 
    -10.29163, -10.16825, -10.04473, -9.921065, -9.79726, -9.673314, 
    -9.549228, -9.424999, -9.300632, -9.176123, -9.051474, -8.926686, 
    -8.801759, -8.676692, -8.551487, -8.426143, -8.300661, -8.175041, 
    -8.049283, -7.923388, -7.797357, -7.671188, -7.544883, -7.418442, 
    -7.291866, -7.165154, -7.038307, -6.911325, -6.78421, -6.65696, 
    -6.529576, -6.40206, -6.27441, -6.146628, -6.018714, -5.890669, 
    -5.762492, -5.634184, -5.505745, -5.377177, -5.248478, -5.119651, 
    -4.990695, -4.861609, -4.732397, -4.603056, -4.473588, -4.343994, 
    -4.214273, -4.084427, -3.954455, -3.824358, -3.694137, -3.563792, 
    -3.433323, -3.302731, -3.172017, -3.041181, -2.910223, -2.779144, 
    -2.647945, -2.516625, -2.385186, -2.253628, -2.121952, -1.990158, 
    -1.858246, -1.726218, -1.594073, -1.461812, -1.329436, -1.196945, 
    -1.064341, -0.9316223, -0.7987911, -0.6658474, -0.5327919, -0.3996252, 
    -0.2663479, -0.1329605, 0.0005363904, 0.1341421, 0.267856, 0.4016776, 
    0.5356061, 0.6696411, 0.8037818, 0.9380276, 1.072378, 1.206832, 1.34139, 
    1.476049, 1.610811, 1.745674, 1.880638, 2.015702, 2.150864, 2.286126, 
    2.421485, 2.556942, 2.692495, 2.828143, 2.963887, 3.099725, 3.235658, 
    3.371683, 3.5078, 3.644009, 3.780308, 3.916698, 4.053177, 4.189745, 
    4.326401, 4.463144, 4.599973, 4.736888, 4.873888, 5.010972, 5.148139, 
    5.285389, 5.422721, 5.560134, 5.697627, 5.8352, 5.972851, 6.11058, 
    6.248387, 6.38627, 6.524228, 6.662261, 6.800367, 6.938547, 7.076799, 
    7.215123, 7.353518, 7.491982, 7.630515, 7.769115, 7.907784, 8.046519, 
    8.18532, 8.324184, 8.463114, 8.602106, 8.74116, 8.880277, 9.019453, 
    9.158689, 9.297984, 9.437336, 9.576746, 9.716211, 9.855733, 9.995308, 
    10.13494, 10.27462, 10.41435, 10.55414, 10.69397, 10.83385, 10.97378, 
    11.11376, 11.25379, 11.39386, 11.53397, 11.67413, 11.81433, 11.95457, 
    12.09485, 12.23518, 12.37554, 12.51594, 12.65637, 12.79685, 12.93736, 
    13.0779, 13.21848, 13.35908, 13.49972, 13.6404, 13.7811, 13.92182, 
    14.06258, 14.20336, 14.34417, 14.48501, 14.62587, 14.76675, 14.90765, 
    15.04858, 15.18952, 15.33048, 15.47147, 15.61247, 15.75348, 15.89451, 
    16.03556, 16.17662, 16.31769, 16.45877, 16.59986, 16.74097, 16.88208, 
    17.0232, 17.16432, 17.30545, 17.44659, 17.58773, 17.72887, 17.87002, 
    18.01116, 18.15231, 18.29345, 18.4346, 18.57574, 18.71687, 18.858, 
    18.99913, 19.14025, 19.28135, 19.42246, 19.56355, 19.70463, 19.8457, 
    19.98676, 20.1278, 20.26883, 20.40984, 20.55084, 20.69181, 20.83278, 
    20.97372, 21.11464, 21.25554, 21.39642, 21.53727, 21.6781, 21.81891, 
    21.95969, 22.10044, 22.24116, 22.38186, 22.52253, 22.66316, 22.80376, 
    22.94433, 23.08487, 23.22538, 23.36584, 23.50627, 23.64667, 23.78702, 
    23.92734, 24.06762, 24.20785, 24.34805, 24.4882, 24.62831, 24.76837, 
    24.90838, 25.04836, 25.18828, 25.32815, 25.46798, 25.60776, 25.74748, 
    25.88715, 26.02678, 26.16634, 26.30585, 26.44531, 26.58471, 26.72405, 
    26.86334, 27.00257, 27.14173, 27.28084, 27.41988, 27.55887, 27.69779, 
    27.83664, 27.97543, 28.11415, 28.25281, 28.3914, 28.52993, 28.66838, 
    28.80676, 28.94507, 29.08331, 29.22148, 29.35958, 29.4976, 29.63555, 
    29.77342, 29.91121, 30.04893, 30.18657, 30.32413, 30.46161, 30.59901, 
    30.73633, 30.87356, 31.01072, 31.14779, 31.28477, 31.42168, 31.55849, 
    31.69522, 31.83186, 31.96842, 32.10488, 32.24126, 32.37754, 32.51374, 
    32.64984, 32.78585, 32.92177, 33.05759, 33.19332, 33.32895, 33.46449, 
    33.59993, 33.73528, 33.87052, 34.00567, 34.14072, 34.27567, 34.41051, 
    34.54526, 34.6799, 34.81444, 34.94888, 35.08321, 35.21745, 35.35157, 
    35.48559, 35.6195, 35.7533, 35.887, 36.02059, 36.15407, 36.28744, 
    36.4207, 36.55385, 36.68689, 36.81981, 36.95263, 37.08532, 37.21791, 
    37.35038, 37.48274, 37.61498, 37.74711, 37.87912, 38.01101, 38.14279, 
    38.27445, 38.40599, 38.53741, 38.6687, 38.79989, 38.93095, 39.06189, 
    39.1927, 39.3234, 39.45397, 39.58442, 39.71474, 39.84494, 39.97502, 
    40.10498, 40.2348, 40.3645, 40.49408, 40.62352, 40.75285, 40.88204, 
    41.0111, 41.14004, 41.26884, 41.39752,
  -16.79756, -16.68194, -16.56618, -16.45026, -16.33419, -16.21798, 
    -16.10161, -15.9851, -15.86844, -15.75163, -15.63467, -15.51756, 
    -15.4003, -15.28289, -15.16534, -15.04763, -14.92978, -14.81177, 
    -14.69362, -14.57532, -14.45688, -14.33828, -14.21954, -14.10064, 
    -13.9816, -13.86242, -13.74308, -13.6236, -13.50397, -13.38419, 
    -13.26426, -13.14419, -13.02397, -12.9036, -12.78309, -12.66243, 
    -12.54162, -12.42067, -12.29957, -12.17832, -12.05693, -11.93539, 
    -11.81371, -11.69188, -11.56991, -11.44779, -11.32553, -11.20312, 
    -11.08057, -10.95787, -10.83503, -10.71205, -10.58892, -10.46565, 
    -10.34223, -10.21868, -10.09498, -9.971136, -9.847153, -9.723026, 
    -9.598759, -9.474349, -9.349798, -9.225107, -9.100275, -8.975303, 
    -8.85019, -8.724938, -8.599546, -8.474015, -8.348345, -8.222537, 
    -8.09659, -7.970505, -7.844282, -7.717922, -7.591425, -7.464791, 
    -7.338021, -7.211114, -7.084073, -6.956895, -6.829583, -6.702136, 
    -6.574554, -6.446839, -6.31899, -6.191008, -6.062893, -5.934646, 
    -5.806266, -5.677755, -5.549113, -5.42034, -5.291437, -5.162403, 
    -5.03324, -4.903948, -4.774527, -4.644977, -4.5153, -4.385496, -4.255564, 
    -4.125506, -3.995322, -3.865012, -3.734577, -3.604017, -3.473334, 
    -3.342526, -3.211596, -3.080542, -2.949367, -2.818069, -2.686651, 
    -2.555112, -2.423452, -2.291673, -2.159775, -2.027758, -1.895623, 
    -1.76337, -1.631001, -1.498515, -1.365913, -1.233196, -1.100364, 
    -0.9674176, -0.8343578, -0.7011849, -0.5678996, -0.4345024, -0.3009939, 
    -0.1673747, -0.0336454, 0.1001934, 0.234141, 0.3681969, 0.5023605, 
    0.636631, 0.7710079, 0.9054906, 1.040078, 1.174771, 1.309567, 1.444466, 
    1.579468, 1.714571, 1.849776, 1.985081, 2.120486, 2.255991, 2.391593, 
    2.527294, 2.663091, 2.798985, 2.934975, 3.07106, 3.207239, 3.343511, 
    3.479877, 3.616334, 3.752883, 3.889522, 4.026252, 4.16307, 4.299977, 
    4.436972, 4.574054, 4.711222, 4.848475, 4.985813, 5.123234, 5.260739, 
    5.398326, 5.535995, 5.673745, 5.811574, 5.949483, 6.087471, 6.225535, 
    6.363677, 6.501894, 6.640187, 6.778554, 6.916994, 7.055508, 7.194093, 
    7.332749, 7.471476, 7.610271, 7.749136, 7.888068, 8.027067, 8.166132, 
    8.305263, 8.444457, 8.583714, 8.723036, 8.862418, 9.001861, 9.141364, 
    9.280927, 9.420547, 9.560225, 9.69996, 9.839749, 9.979594, 10.11949, 
    10.25944, 10.39945, 10.5395, 10.67961, 10.81976, 10.95996, 11.10021, 
    11.24051, 11.38085, 11.52124, 11.66167, 11.80214, 11.94266, 12.08322, 
    12.22381, 12.36445, 12.50513, 12.64584, 12.78658, 12.92737, 13.06819, 
    13.20904, 13.34992, 13.49084, 13.63179, 13.77276, 13.91377, 14.0548, 
    14.19586, 14.33695, 14.47806, 14.6192, 14.76036, 14.90154, 15.04274, 
    15.18396, 15.32521, 15.46647, 15.60774, 15.74904, 15.89035, 16.03167, 
    16.17301, 16.31436, 16.45572, 16.59709, 16.73847, 16.87987, 17.02126, 
    17.16267, 17.30408, 17.4455, 17.58691, 17.72834, 17.86976, 18.01118, 
    18.15261, 18.29403, 18.43546, 18.57688, 18.71829, 18.8597, 19.0011, 
    19.1425, 19.28389, 19.42527, 19.56664, 19.708, 19.84935, 19.99068, 
    20.13201, 20.27331, 20.41461, 20.55588, 20.69714, 20.83838, 20.9796, 
    21.1208, 21.26197, 21.40313, 21.54426, 21.68537, 21.82645, 21.96751, 
    22.10854, 22.24954, 22.39051, 22.53145, 22.67236, 22.81324, 22.95409, 
    23.0949, 23.23568, 23.37642, 23.51713, 23.6578, 23.79843, 23.93902, 
    24.07957, 24.22008, 24.36055, 24.50097, 24.64135, 24.78168, 24.92197, 
    25.06222, 25.20241, 25.34256, 25.48266, 25.6227, 25.7627, 25.90264, 
    26.04253, 26.18237, 26.32215, 26.46187, 26.60154, 26.74115, 26.88071, 
    27.0202, 27.15963, 27.29901, 27.43832, 27.57757, 27.71675, 27.85587, 
    27.99492, 28.13391, 28.27283, 28.41169, 28.55047, 28.68919, 28.82783, 
    28.96641, 29.10491, 29.24334, 29.38169, 29.51998, 29.65818, 29.79631, 
    29.93436, 30.07234, 30.21023, 30.34805, 30.48579, 30.62344, 30.76102, 
    30.89851, 31.03592, 31.17324, 31.31048, 31.44764, 31.5847, 31.72169, 
    31.85858, 31.99538, 32.1321, 32.26872, 32.40526, 32.5417, 32.67805, 
    32.81431, 32.95047, 33.08654, 33.22252, 33.35839, 33.49418, 33.62986, 
    33.76545, 33.90094, 34.03633, 34.17162, 34.30681, 34.44189, 34.57688, 
    34.71176, 34.84654, 34.98122, 35.11579, 35.25026, 35.38462, 35.51887, 
    35.65302, 35.78706, 35.92099, 36.05481, 36.18852, 36.32212, 36.45561, 
    36.58899, 36.72226, 36.85541, 36.98846, 37.12138, 37.2542, 37.3869, 
    37.51948, 37.65195, 37.7843, 37.91653, 38.04865, 38.18065, 38.31253, 
    38.44429, 38.57593, 38.70745, 38.83885, 38.97012, 39.10128, 39.23232, 
    39.36323, 39.49401, 39.62468, 39.75522, 39.88563, 40.01592, 40.14609, 
    40.27613, 40.40604, 40.53582, 40.66548, 40.79501, 40.92441, 41.05368, 
    41.18282, 41.31184, 41.44072,
  -16.8568, -16.74104, -16.62514, -16.50908, -16.39287, -16.27652, -16.16001, 
    -16.04335, -15.92655, -15.80959, -15.69249, -15.57523, -15.45782, 
    -15.34027, -15.22257, -15.10471, -14.98671, -14.86856, -14.75026, 
    -14.63181, -14.51321, -14.39446, -14.27556, -14.15651, -14.03732, 
    -13.91797, -13.79848, -13.67884, -13.55905, -13.43912, -13.31903, 
    -13.1988, -13.07842, -12.95789, -12.83721, -12.71639, -12.59542, 
    -12.4743, -12.35304, -12.23163, -12.11007, -11.98836, -11.86651, 
    -11.74452, -11.62237, -11.50009, -11.37765, -11.25507, -11.13235, 
    -11.00948, -10.88647, -10.76331, -10.64001, -10.51656, -10.39297, 
    -10.26923, -10.14536, -10.02134, -9.897173, -9.772866, -9.648417, 
    -9.523827, -9.399095, -9.27422, -9.149204, -9.024047, -8.898749, 
    -8.773312, -8.647733, -8.522015, -8.396156, -8.270159, -8.144022, 
    -8.017747, -7.891333, -7.764781, -7.638092, -7.511264, -7.3843, 
    -7.257199, -7.129961, -7.002588, -6.875079, -6.747434, -6.619654, 
    -6.49174, -6.363691, -6.235508, -6.107193, -5.978743, -5.850161, 
    -5.721447, -5.5926, -5.463623, -5.334514, -5.205274, -5.075903, 
    -4.946404, -4.816774, -4.687016, -4.557129, -4.427114, -4.296971, 
    -4.166701, -4.036304, -3.905781, -3.775132, -3.644357, -3.513458, 
    -3.382435, -3.251287, -3.120016, -2.988622, -2.857106, -2.725468, 
    -2.593708, -2.461828, -2.329827, -2.197706, -2.065466, -1.933108, 
    -1.800631, -1.668036, -1.535324, -1.402496, -1.269552, -1.136492, 
    -1.003318, -0.8700287, -0.7366261, -0.6031104, -0.4694822, -0.335742, 
    -0.2018905, -0.0679282, 0.06614419, 0.2003261, 0.3346169, 0.469016, 
    0.6035227, 0.7381364, 0.8728565, 1.007682, 1.142613, 1.277649, 1.412788, 
    1.54803, 1.683375, 1.818821, 1.954369, 2.090017, 2.225765, 2.361611, 
    2.497556, 2.633599, 2.769739, 2.905975, 3.042307, 3.178733, 3.315254, 
    3.451868, 3.588575, 3.725373, 3.862263, 3.999243, 4.136313, 4.273472, 
    4.41072, 4.548054, 4.685476, 4.822983, 4.960576, 5.098253, 5.236013, 
    5.373857, 5.511782, 5.649788, 5.787876, 5.926043, 6.064288, 6.202612, 
    6.341013, 6.479491, 6.618044, 6.756672, 6.895374, 7.034149, 7.172997, 
    7.311915, 7.450905, 7.589965, 7.729093, 7.86829, 8.007554, 8.146884, 
    8.28628, 8.42574, 8.565265, 8.704853, 8.844502, 8.984213, 9.123984, 
    9.263815, 9.403705, 9.543652, 9.683656, 9.823715, 9.96383, 10.104, 
    10.24422, 10.3845, 10.52482, 10.6652, 10.80562, 10.9461, 11.08662, 
    11.22719, 11.36781, 11.50847, 11.64917, 11.78992, 11.93071, 12.07154, 
    12.21242, 12.35333, 12.49428, 12.63527, 12.77629, 12.91735, 13.05844, 
    13.19957, 13.34073, 13.48193, 13.62315, 13.76441, 13.90569, 14.047, 
    14.18834, 14.3297, 14.47109, 14.61251, 14.75395, 14.89541, 15.03689, 
    15.17839, 15.31991, 15.46145, 15.60301, 15.74458, 15.88617, 16.02777, 
    16.16939, 16.31102, 16.45266, 16.59431, 16.73598, 16.87765, 17.01932, 
    17.16101, 17.3027, 17.4444, 17.5861, 17.7278, 17.8695, 18.01121, 
    18.15291, 18.29462, 18.43632, 18.57802, 18.71971, 18.8614, 19.00309, 
    19.14476, 19.28643, 19.42809, 19.56975, 19.71139, 19.85301, 19.99463, 
    20.13623, 20.27782, 20.41939, 20.56094, 20.70248, 20.844, 20.98549, 
    21.12697, 21.26843, 21.40986, 21.55127, 21.69266, 21.83402, 21.97536, 
    22.11666, 22.25794, 22.39919, 22.54041, 22.6816, 22.82275, 22.96388, 
    23.10497, 23.24602, 23.38704, 23.52802, 23.66896, 23.80987, 23.95074, 
    24.09156, 24.23235, 24.37309, 24.51378, 24.65444, 24.79505, 24.93561, 
    25.07612, 25.21659, 25.35701, 25.49738, 25.6377, 25.77796, 25.91818, 
    26.05834, 26.19844, 26.3385, 26.47849, 26.61843, 26.75831, 26.89813, 
    27.03789, 27.17759, 27.31723, 27.45681, 27.59632, 27.73577, 27.87516, 
    28.01448, 28.15373, 28.29292, 28.43204, 28.57108, 28.71006, 28.84897, 
    28.98781, 29.12657, 29.26526, 29.40388, 29.54242, 29.68089, 29.81927, 
    29.95758, 30.09582, 30.23397, 30.37205, 30.51004, 30.64795, 30.78578, 
    30.92353, 31.0612, 31.19877, 31.33627, 31.47367, 31.611, 31.74823, 
    31.88537, 32.02243, 32.1594, 32.29627, 32.43306, 32.56975, 32.70635, 
    32.84285, 32.97926, 33.11558, 33.2518, 33.38793, 33.52396, 33.65989, 
    33.79572, 33.93145, 34.06708, 34.20261, 34.33804, 34.47337, 34.6086, 
    34.74372, 34.87874, 35.01365, 35.14846, 35.28316, 35.41776, 35.55225, 
    35.68663, 35.82091, 35.95507, 36.08913, 36.22307, 36.35691, 36.49063, 
    36.62424, 36.75774, 36.89112, 37.02439, 37.15755, 37.29059, 37.42352, 
    37.55632, 37.68902, 37.82159, 37.95405, 38.08639, 38.21861, 38.35072, 
    38.4827, 38.61456, 38.7463, 38.87792, 39.00941, 39.14079, 39.27204, 
    39.40317, 39.53417, 39.66505, 39.79581, 39.92644, 40.05694, 40.18732, 
    40.31757, 40.44769, 40.57768, 40.70755, 40.83729, 40.9669, 41.09638, 
    41.22573, 41.35495, 41.48403,
  -16.91617, -16.80028, -16.68423, -16.56804, -16.45169, -16.33519, 
    -16.21854, -16.10174, -15.98479, -15.86769, -15.75044, -15.63304, 
    -15.51549, -15.39778, -15.27993, -15.16193, -15.04378, -14.92548, 
    -14.80702, -14.68842, -14.56967, -14.45077, -14.33172, -14.21251, 
    -14.09317, -13.97367, -13.85402, -13.73422, -13.61427, -13.49418, 
    -13.37393, -13.25354, -13.133, -13.01231, -12.89147, -12.77048, 
    -12.64935, -12.52807, -12.40664, -12.28506, -12.16334, -12.04147, 
    -11.91945, -11.79728, -11.67497, -11.55251, -11.42991, -11.30716, 
    -11.18426, -11.06122, -10.93803, -10.8147, -10.69122, -10.5676, 
    -10.44383, -10.31992, -10.19587, -10.07167, -9.947323, -9.822837, 
    -9.698207, -9.573434, -9.448519, -9.323462, -9.198261, -9.07292, 
    -8.947436, -8.821813, -8.696047, -8.570141, -8.444094, -8.317907, 
    -8.191581, -8.065115, -7.93851, -7.811766, -7.684884, -7.557863, 
    -7.430705, -7.303409, -7.175975, -7.048405, -6.920699, -6.792856, 
    -6.664878, -6.536764, -6.408515, -6.280132, -6.151614, -6.022963, 
    -5.894177, -5.765259, -5.636209, -5.507025, -5.37771, -5.248264, 
    -5.118687, -4.988978, -4.85914, -4.729172, -4.599075, -4.468849, 
    -4.338494, -4.208012, -4.077402, -3.946665, -3.815802, -3.684812, 
    -3.553697, -3.422457, -3.291092, -3.159603, -3.027991, -2.896255, 
    -2.764397, -2.632416, -2.500314, -2.368092, -2.235748, -2.103285, 
    -1.970702, -1.838, -1.70518, -1.572242, -1.439186, -1.306015, -1.172727, 
    -1.039323, -0.9058046, -0.7721717, -0.6384251, -0.5045653, -0.3705929, 
    -0.2365085, -0.1023127, 0.03199387, 0.1664106, 0.3009368, 0.435572, 
    0.5703154, 0.7051665, 0.8401246, 0.9751891, 1.110359, 1.245634, 1.381014, 
    1.516497, 1.652084, 1.787773, 1.923563, 2.059455, 2.195446, 2.331538, 
    2.467729, 2.604017, 2.740404, 2.876887, 3.013466, 3.150141, 3.28691, 
    3.423774, 3.56073, 3.697779, 3.83492, 3.972152, 4.109474, 4.246886, 
    4.384386, 4.521975, 4.65965, 4.797412, 4.93526, 5.073193, 5.21121, 
    5.34931, 5.487493, 5.625758, 5.764103, 5.902529, 6.041034, 6.179617, 
    6.318279, 6.457017, 6.595831, 6.734721, 6.873685, 7.012723, 7.151834, 
    7.291016, 7.43027, 7.569594, 7.708987, 7.848449, 7.987978, 8.127575, 
    8.267238, 8.406965, 8.546757, 8.686612, 8.82653, 8.966509, 9.106549, 
    9.24665, 9.386808, 9.527025, 9.667299, 9.80763, 9.948016, 10.08846, 
    10.22895, 10.3695, 10.5101, 10.65075, 10.79144, 10.93219, 11.07299, 
    11.21383, 11.35472, 11.49566, 11.63664, 11.77766, 11.91873, 12.05983, 
    12.20098, 12.34217, 12.48339, 12.62466, 12.76596, 12.9073, 13.04867, 
    13.19007, 13.33151, 13.47299, 13.61449, 13.75602, 13.89758, 14.03917, 
    14.18079, 14.32243, 14.4641, 14.6058, 14.74751, 14.88925, 15.03101, 
    15.1728, 15.3146, 15.45642, 15.59825, 15.74011, 15.88198, 16.02386, 
    16.16576, 16.30767, 16.44959, 16.59152, 16.73347, 16.87542, 17.01738, 
    17.15935, 17.30132, 17.44329, 17.58527, 17.72726, 17.86924, 18.01123, 
    18.15322, 18.2952, 18.43719, 18.57916, 18.72114, 18.86311, 19.00508, 
    19.14704, 19.28899, 19.43093, 19.57286, 19.71478, 19.85669, 19.99858, 
    20.14047, 20.28233, 20.42418, 20.56602, 20.70784, 20.84963, 20.99141, 
    21.13317, 21.27491, 21.41662, 21.55831, 21.69997, 21.84161, 21.98323, 
    22.12481, 22.26637, 22.4079, 22.54939, 22.69086, 22.83229, 22.9737, 
    23.11506, 23.25639, 23.39769, 23.53895, 23.68017, 23.82135, 23.96249, 
    24.10359, 24.24465, 24.38567, 24.52664, 24.66757, 24.80845, 24.94929, 
    25.09007, 25.23082, 25.37151, 25.51215, 25.65274, 25.79328, 25.93376, 
    26.07419, 26.21457, 26.35489, 26.49516, 26.63537, 26.77552, 26.91561, 
    27.05564, 27.19561, 27.33551, 27.47536, 27.61514, 27.75486, 27.89451, 
    28.0341, 28.17362, 28.31307, 28.45245, 28.59176, 28.731, 28.87018, 
    29.00928, 29.1483, 29.28725, 29.42613, 29.56493, 29.70366, 29.84231, 
    29.98088, 30.11937, 30.25779, 30.39612, 30.53437, 30.67254, 30.81063, 
    30.94863, 31.08655, 31.22438, 31.36213, 31.4998, 31.63737, 31.77486, 
    31.91225, 32.04956, 32.18678, 32.32391, 32.46094, 32.59788, 32.73473, 
    32.87149, 33.00814, 33.14471, 33.28118, 33.41755, 33.55382, 33.68999, 
    33.82607, 33.96205, 34.09792, 34.2337, 34.36937, 34.50494, 34.64041, 
    34.77577, 34.91103, 35.04618, 35.18123, 35.31617, 35.45101, 35.58573, 
    35.72035, 35.85486, 35.98926, 36.12355, 36.25772, 36.39179, 36.52575, 
    36.65959, 36.79332, 36.92693, 37.06043, 37.19382, 37.32709, 37.46024, 
    37.59328, 37.7262, 37.859, 37.99168, 38.12424, 38.25669, 38.38902, 
    38.52122, 38.6533, 38.78526, 38.9171, 39.04882, 39.18041, 39.31188, 
    39.44323, 39.57445, 39.70554, 39.83651, 39.96735, 40.09807, 40.22866, 
    40.35912, 40.48946, 40.61966, 40.74974, 40.87969, 41.00951, 41.13919, 
    41.26875, 41.39817, 41.52747,
  -16.97568, -16.85965, -16.74346, -16.62712, -16.51064, -16.394, -16.2772, 
    -16.16026, -16.04317, -15.92592, -15.80853, -15.69098, -15.57328, 
    -15.45543, -15.33743, -15.21928, -15.10098, -14.98253, -14.86392, 
    -14.74517, -14.62627, -14.50721, -14.38801, -14.26865, -14.14915, 
    -14.02949, -13.90969, -13.78973, -13.66963, -13.54937, -13.42897, 
    -13.30842, -13.18771, -13.06686, -12.94586, -12.82471, -12.70342, 
    -12.58197, -12.46038, -12.33863, -12.21674, -12.0947, -11.97252, 
    -11.85018, -11.7277, -11.60507, -11.4823, -11.35938, -11.23631, 
    -11.11309, -10.98973, -10.86622, -10.74257, -10.61877, -10.49483, 
    -10.37074, -10.2465, -10.12213, -9.997603, -9.872936, -9.748126, 
    -9.623171, -9.498074, -9.372832, -9.247448, -9.121922, -8.996253, 
    -8.870441, -8.74449, -8.618395, -8.49216, -8.365784, -8.239267, 
    -8.112611, -7.985814, -7.858878, -7.731802, -7.604588, -7.477235, 
    -7.349743, -7.222114, -7.094347, -6.966444, -6.838402, -6.710225, 
    -6.581912, -6.453463, -6.324878, -6.196158, -6.067304, -5.938315, 
    -5.809193, -5.679938, -5.550549, -5.421028, -5.291374, -5.161589, 
    -5.031673, -4.901625, -4.771448, -4.64114, -4.510702, -4.380136, 
    -4.249441, -4.118617, -3.987666, -3.856588, -3.725383, -3.594051, 
    -3.462594, -3.331012, -3.199304, -3.067472, -2.935517, -2.803438, 
    -2.671237, -2.538913, -2.406467, -2.2739, -2.141213, -2.008405, 
    -1.875478, -1.742432, -1.609267, -1.475984, -1.342584, -1.209068, 
    -1.075435, -0.941686, -0.8078224, -0.6738443, -0.5397524, -0.4055473, 
    -0.2712294, -0.1367996, -0.002258277, 0.1323938, 0.2671561, 0.4020279, 
    0.5370086, 0.6720977, 0.8072944, 0.942598, 1.078008, 1.213524, 1.349144, 
    1.484869, 1.620698, 1.75663, 1.892664, 2.0288, 2.165036, 2.301373, 
    2.437809, 2.574345, 2.710978, 2.847709, 2.984537, 3.12146, 3.258479, 
    3.395593, 3.5328, 3.6701, 3.807492, 3.944977, 4.082551, 4.220217, 
    4.357971, 4.495814, 4.633745, 4.771762, 4.909866, 5.048055, 5.186329, 
    5.324687, 5.463128, 5.601651, 5.740256, 5.878941, 6.017706, 6.15655, 
    6.295473, 6.434473, 6.573549, 6.712701, 6.851928, 6.99123, 7.130604, 
    7.270051, 7.409569, 7.549158, 7.688818, 7.828545, 7.968341, 8.108205, 
    8.248135, 8.388129, 8.52819, 8.668313, 8.8085, 8.948749, 9.089059, 
    9.229428, 9.369858, 9.510345, 9.650891, 9.791493, 9.932151, 10.07286, 
    10.21363, 10.35445, 10.49532, 10.63624, 10.77722, 10.91824, 11.05931, 
    11.20043, 11.34159, 11.48281, 11.62406, 11.76536, 11.9067, 12.04808, 
    12.18951, 12.33097, 12.47248, 12.61402, 12.7556, 12.89721, 13.03886, 
    13.18055, 13.32226, 13.46402, 13.6058, 13.74761, 13.88945, 14.03132, 
    14.17322, 14.31514, 14.45709, 14.59906, 14.74106, 14.88308, 15.02512, 
    15.16718, 15.30927, 15.45137, 15.59348, 15.73562, 15.87777, 16.01994, 
    16.16212, 16.30431, 16.44651, 16.58873, 16.73095, 16.87318, 17.01543, 
    17.15767, 17.29993, 17.44219, 17.58445, 17.72672, 17.86898, 18.01125, 
    18.15352, 18.29579, 18.43805, 18.58032, 18.72257, 18.86483, 19.00707, 
    19.14931, 19.29155, 19.43377, 19.57598, 19.71819, 19.86038, 20.00255, 
    20.14472, 20.28687, 20.429, 20.57111, 20.71321, 20.85529, 20.99735, 
    21.13939, 21.2814, 21.4234, 21.56537, 21.70731, 21.84923, 21.99113, 
    22.13299, 22.27483, 22.41663, 22.55841, 22.70016, 22.84187, 22.98355, 
    23.12519, 23.2668, 23.40837, 23.54991, 23.69141, 23.83286, 23.97428, 
    24.11566, 24.25699, 24.39829, 24.53954, 24.68074, 24.8219, 24.96301, 
    25.10407, 25.24508, 25.38605, 25.52697, 25.66783, 25.80864, 25.9494, 
    26.0901, 26.23075, 26.37135, 26.51188, 26.65236, 26.79278, 26.93314, 
    27.07344, 27.21368, 27.35386, 27.49397, 27.63402, 27.774, 27.91392, 
    28.05378, 28.19356, 28.33328, 28.47293, 28.6125, 28.75201, 28.89145, 
    29.03081, 29.1701, 29.30931, 29.44846, 29.58752, 29.72651, 29.86542, 
    30.00425, 30.143, 30.28168, 30.42027, 30.55878, 30.6972, 30.83555, 
    30.97381, 31.11199, 31.25008, 31.38808, 31.526, 31.66383, 31.80157, 
    31.93922, 32.07678, 32.21425, 32.35162, 32.48891, 32.6261, 32.7632, 
    32.9002, 33.03711, 33.17393, 33.31064, 33.44726, 33.58378, 33.7202, 
    33.85652, 33.99274, 34.12886, 34.26488, 34.40079, 34.53661, 34.67232, 
    34.80792, 34.94342, 35.07881, 35.2141, 35.34928, 35.48435, 35.61931, 
    35.75417, 35.88891, 36.02355, 36.15807, 36.29248, 36.42678, 36.56097, 
    36.69505, 36.82901, 36.96285, 37.09658, 37.23019, 37.36369, 37.49707, 
    37.63034, 37.76348, 37.89651, 38.02942, 38.16221, 38.29488, 38.42743, 
    38.55985, 38.69216, 38.82434, 38.9564, 39.08833, 39.22015, 39.35183, 
    39.4834, 39.61483, 39.74615, 39.87733, 40.00839, 40.13932, 40.27012, 
    40.4008, 40.53135, 40.66176, 40.79205, 40.92221, 41.05223, 41.18213, 
    41.31189, 41.44152, 41.57103,
  -17.03533, -16.91915, -16.80283, -16.68635, -16.56972, -16.45294, -16.336, 
    -16.21892, -16.10168, -15.98429, -15.86675, -15.74906, -15.63121, 
    -15.51322, -15.39507, -15.27677, -15.15832, -15.03971, -14.92096, 
    -14.80206, -14.683, -14.56379, -14.44443, -14.32492, -14.20526, 
    -14.08545, -13.96549, -13.84538, -13.72512, -13.6047, -13.48414, 
    -13.36343, -13.24257, -13.12155, -13.00039, -12.87908, -12.75762, 
    -12.63601, -12.51425, -12.39234, -12.27028, -12.14807, -12.02572, 
    -11.90322, -11.78057, -11.65777, -11.53482, -11.41173, -11.28849, 
    -11.1651, -11.04156, -10.91788, -10.79405, -10.67008, -10.54596, 
    -10.42169, -10.29728, -10.17272, -10.04802, -9.923168, -9.798176, 
    -9.673038, -9.547758, -9.422333, -9.296764, -9.171053, -9.045198, 
    -8.919201, -8.793061, -8.666779, -8.540355, -8.413789, -8.287082, 
    -8.160234, -8.033246, -7.906117, -7.778848, -7.651439, -7.523891, 
    -7.396204, -7.268379, -7.140415, -7.012313, -6.884074, -6.755697, 
    -6.627184, -6.498534, -6.369748, -6.240826, -6.111769, -5.982576, 
    -5.85325, -5.723789, -5.594194, -5.464467, -5.334606, -5.204613, 
    -5.074487, -4.944231, -4.813842, -4.683323, -4.552674, -4.421896, 
    -4.290987, -4.15995, -4.028784, -3.897491, -3.766069, -3.634521, 
    -3.502846, -3.371046, -3.23912, -3.107068, -2.974892, -2.842592, 
    -2.710169, -2.577623, -2.444954, -2.312164, -2.179252, -2.046219, 
    -1.913066, -1.779793, -1.646401, -1.512891, -1.379262, -1.245516, 
    -1.111653, -0.9776738, -0.8435789, -0.7093688, -0.5750443, -0.4406058, 
    -0.306054, -0.1713895, -0.03661293, 0.09827511, 0.233274, 0.368383, 
    0.5036017, 0.6389292, 0.7743651, 0.9099085, 1.045559, 1.181316, 1.317178, 
    1.453145, 1.589217, 1.725392, 1.861671, 1.998051, 2.134533, 2.271116, 
    2.407799, 2.544581, 2.681463, 2.818442, 2.955518, 3.092692, 3.22996, 
    3.367325, 3.504783, 3.642335, 3.77998, 3.917717, 4.055546, 4.193465, 
    4.331474, 4.469572, 4.607758, 4.746032, 4.884392, 5.022839, 5.161371, 
    5.299987, 5.438687, 5.577469, 5.716333, 5.855279, 5.994305, 6.133411, 
    6.272595, 6.411857, 6.551196, 6.690612, 6.830102, 6.969668, 7.109307, 
    7.249019, 7.388803, 7.528658, 7.668583, 7.808578, 7.948641, 8.088773, 
    8.228971, 8.369234, 8.509563, 8.649956, 8.790413, 8.930931, 9.071511, 
    9.212152, 9.352853, 9.493612, 9.63443, 9.775305, 9.916235, 10.05722, 
    10.19826, 10.33935, 10.4805, 10.6217, 10.76295, 10.90424, 11.04559, 
    11.18698, 11.32842, 11.46991, 11.61144, 11.75302, 11.89464, 12.0363, 
    12.178, 12.31974, 12.46152, 12.60334, 12.7452, 12.8871, 13.02902, 
    13.17099, 13.31299, 13.45502, 13.59708, 13.73917, 13.88129, 14.02344, 
    14.16562, 14.30782, 14.45005, 14.59231, 14.73459, 14.87689, 15.01921, 
    15.16155, 15.30392, 15.4463, 15.5887, 15.73112, 15.87355, 16.016, 
    16.15846, 16.30094, 16.44342, 16.58592, 16.72843, 16.87094, 17.01347, 
    17.156, 17.29854, 17.44108, 17.58362, 17.72617, 17.86872, 18.01127, 
    18.15383, 18.29638, 18.43892, 18.58147, 18.72401, 18.86655, 19.00908, 
    19.1516, 19.29412, 19.43662, 19.57912, 19.7216, 19.86407, 20.00653, 
    20.14898, 20.29141, 20.43383, 20.57622, 20.7186, 20.86096, 21.00331, 
    21.14562, 21.28792, 21.4302, 21.57245, 21.71467, 21.85687, 21.99905, 
    22.14119, 22.28331, 22.4254, 22.56745, 22.70948, 22.85147, 22.99343, 
    23.13535, 23.27724, 23.41909, 23.56091, 23.70268, 23.84442, 23.98611, 
    24.12777, 24.26938, 24.41095, 24.55247, 24.69395, 24.83539, 24.97677, 
    25.11811, 25.2594, 25.40064, 25.54183, 25.68297, 25.82405, 25.96508, 
    26.10606, 26.24698, 26.38785, 26.52866, 26.66941, 26.8101, 26.95073, 
    27.0913, 27.23181, 27.37226, 27.51264, 27.65296, 27.79321, 27.9334, 
    28.07352, 28.21357, 28.35356, 28.49347, 28.63331, 28.77309, 28.91279, 
    29.05241, 29.19197, 29.33145, 29.47085, 29.61018, 29.74943, 29.8886, 
    30.02769, 30.16671, 30.30564, 30.44449, 30.58326, 30.72194, 30.86055, 
    30.99907, 31.1375, 31.27585, 31.41411, 31.55228, 31.69036, 31.82836, 
    31.96626, 32.10408, 32.2418, 32.37943, 32.51697, 32.65441, 32.79176, 
    32.92901, 33.06617, 33.20323, 33.34019, 33.47706, 33.61383, 33.7505, 
    33.88706, 34.02353, 34.15989, 34.29615, 34.43232, 34.56837, 34.70432, 
    34.84016, 34.97591, 35.11154, 35.24707, 35.38248, 35.5178, 35.653, 
    35.78809, 35.92307, 36.05794, 36.1927, 36.32735, 36.46188, 36.5963, 
    36.73061, 36.8648, 36.99887, 37.13284, 37.26668, 37.40041, 37.53402, 
    37.66751, 37.80088, 37.93414, 38.06727, 38.20028, 38.33318, 38.46595, 
    38.5986, 38.73112, 38.86353, 38.99581, 39.12796, 39.26, 39.3919, 
    39.52369, 39.65534, 39.78687, 39.91827, 40.04954, 40.18069, 40.3117, 
    40.44259, 40.57335, 40.70398, 40.83448, 40.96484, 41.09508, 41.22519, 
    41.35516, 41.485, 41.6147,
  -17.09511, -16.97879, -16.86233, -16.74571, -16.62894, -16.51202, 
    -16.39494, -16.27771, -16.16033, -16.0428, -15.92511, -15.80727, 
    -15.68928, -15.57114, -15.45284, -15.33439, -15.21579, -15.09704, 
    -14.97813, -14.85908, -14.73987, -14.62051, -14.501, -14.38133, 
    -14.26152, -14.14155, -14.02143, -13.90116, -13.78074, -13.66017, 
    -13.53945, -13.41858, -13.29755, -13.17638, -13.05505, -12.93358, 
    -12.81195, -12.69018, -12.56825, -12.44618, -12.32395, -12.20158, 
    -12.07906, -11.95639, -11.83356, -11.7106, -11.58748, -11.46421, 
    -11.3408, -11.21724, -11.09353, -10.96967, -10.84567, -10.72151, 
    -10.59722, -10.47277, -10.34818, -10.22344, -10.09856, -9.973532, 
    -9.848357, -9.723039, -9.597574, -9.471966, -9.346212, -9.220315, 
    -9.094275, -8.96809, -8.841763, -8.715292, -8.588678, -8.461924, 
    -8.335026, -8.207987, -8.080806, -7.953484, -7.826022, -7.698419, 
    -7.570676, -7.442793, -7.314771, -7.186609, -7.05831, -6.929872, 
    -6.801295, -6.672581, -6.54373, -6.414742, -6.285618, -6.156357, 
    -6.026961, -5.89743, -5.767764, -5.637963, -5.508028, -5.377959, 
    -5.247757, -5.117423, -4.986956, -4.856358, -4.725627, -4.594766, 
    -4.463774, -4.332652, -4.201401, -4.07002, -3.938511, -3.806873, 
    -3.675108, -3.543215, -3.411196, -3.27905, -3.146779, -3.014382, 
    -2.881861, -2.749216, -2.616446, -2.483554, -2.350539, -2.217402, 
    -2.084144, -1.950765, -1.817265, -1.683645, -1.549906, -1.416048, 
    -1.282072, -1.147979, -1.013769, -0.8794419, -0.7449993, -0.6104415, 
    -0.4757692, -0.3409829, -0.2060832, -0.07107077, 0.06405377, 0.1992898, 
    0.3346367, 0.4700938, 0.6056604, 0.741336, 0.8771198, 1.013011, 1.14901, 
    1.285114, 1.421325, 1.55764, 1.694059, 1.830582, 1.967208, 2.103936, 
    2.240766, 2.377696, 2.514726, 2.651856, 2.789084, 2.92641, 3.063834, 
    3.201354, 3.338969, 3.476679, 3.614484, 3.752382, 3.890373, 4.028455, 
    4.166629, 4.304893, 4.443247, 4.58169, 4.720221, 4.858839, 4.997543, 
    5.136334, 5.275209, 5.414168, 5.553211, 5.692336, 5.831542, 5.97083, 
    6.110198, 6.249645, 6.38917, 6.528772, 6.668452, 6.808208, 6.948038, 
    7.087942, 7.22792, 7.36797, 7.508092, 7.648284, 7.788547, 7.928878, 
    8.069278, 8.209744, 8.350278, 8.490876, 8.631539, 8.772266, 8.913056, 
    9.053908, 9.19482, 9.335793, 9.476826, 9.617916, 9.759064, 9.900268, 
    10.04153, 10.18284, 10.32421, 10.46563, 10.6071, 10.74863, 10.8902, 
    11.03182, 11.17349, 11.31521, 11.45697, 11.59878, 11.74064, 11.88253, 
    12.02447, 12.16645, 12.30847, 12.45053, 12.59263, 12.73477, 12.87694, 
    13.01915, 13.1614, 13.30367, 13.44599, 13.58833, 13.7307, 13.8731, 
    14.01553, 14.15799, 14.30048, 14.44299, 14.58553, 14.72809, 14.87067, 
    15.01328, 15.15591, 15.29855, 15.44122, 15.5839, 15.7266, 15.86932, 
    16.01205, 16.15479, 16.29755, 16.44032, 16.5831, 16.72589, 16.86869, 
    17.0115, 17.15432, 17.29714, 17.43996, 17.58279, 17.72563, 17.86846, 
    18.0113, 18.15413, 18.29697, 18.4398, 18.58263, 18.72545, 18.86827, 
    19.01109, 19.15389, 19.29669, 19.43948, 19.58226, 19.72503, 19.86779, 
    20.01053, 20.15326, 20.29597, 20.43867, 20.58135, 20.72401, 20.86666, 
    21.00928, 21.15188, 21.29446, 21.43702, 21.57955, 21.72206, 21.86454, 
    22.007, 22.14943, 22.29182, 22.43419, 22.57653, 22.71883, 22.8611, 
    23.00334, 23.14555, 23.28772, 23.42985, 23.57194, 23.71399, 23.85601, 
    23.99798, 24.13992, 24.28181, 24.42365, 24.56545, 24.70721, 24.84892, 
    24.99058, 25.1322, 25.27376, 25.41528, 25.55674, 25.69816, 25.83952, 
    25.98082, 26.12207, 26.26327, 26.40441, 26.54549, 26.68651, 26.82747, 
    26.96838, 27.10922, 27.25, 27.39071, 27.53137, 27.67196, 27.81248, 
    27.95294, 28.09332, 28.23364, 28.3739, 28.51408, 28.65419, 28.79423, 
    28.93419, 29.07409, 29.21391, 29.35365, 29.49331, 29.63291, 29.77242, 
    29.91185, 30.05121, 30.19048, 30.32968, 30.46879, 30.60782, 30.74677, 
    30.88563, 31.0244, 31.16309, 31.3017, 31.44022, 31.57864, 31.71698, 
    31.85523, 31.99339, 32.13146, 32.26944, 32.40732, 32.54511, 32.68281, 
    32.82041, 32.95791, 33.09532, 33.23263, 33.36984, 33.50696, 33.64397, 
    33.78088, 33.9177, 34.05441, 34.19102, 34.32753, 34.46393, 34.60023, 
    34.73642, 34.87251, 35.00849, 35.14437, 35.28013, 35.41579, 35.55134, 
    35.68678, 35.82211, 35.95733, 36.09243, 36.22743, 36.36231, 36.49708, 
    36.63173, 36.76627, 36.9007, 37.03501, 37.1692, 37.30327, 37.43723, 
    37.57107, 37.70479, 37.83839, 37.97187, 38.10523, 38.23847, 38.37159, 
    38.50459, 38.63745, 38.77021, 38.90283, 39.03534, 39.16771, 39.29996, 
    39.43209, 39.56409, 39.69596, 39.82771, 39.95932, 40.09081, 40.22217, 
    40.3534, 40.4845, 40.61547, 40.74632, 40.87703, 41.0076, 41.13805, 
    41.26836, 41.39854, 41.52859, 41.6585,
  -17.15502, -17.03857, -16.92197, -16.80521, -16.6883, -16.57123, -16.45401, 
    -16.33664, -16.21912, -16.10144, -15.98361, -15.86562, -15.74749, 
    -15.62919, -15.51075, -15.39215, -15.2734, -15.1545, -15.03545, 
    -14.91624, -14.79688, -14.67736, -14.5577, -14.43788, -14.31791, 
    -14.19779, -14.07751, -13.95708, -13.83651, -13.71578, -13.59489, 
    -13.47386, -13.35268, -13.23134, -13.10985, -12.98821, -12.86642, 
    -12.74448, -12.62239, -12.50015, -12.37776, -12.25522, -12.13253, 
    -12.00969, -11.8867, -11.76356, -11.64027, -11.51683, -11.39324, 
    -11.26951, -11.14563, -11.02159, -10.89741, -10.77309, -10.64861, 
    -10.52399, -10.39922, -10.2743, -10.14924, -10.02403, -9.898672, 
    -9.77317, -9.647523, -9.521729, -9.395792, -9.26971, -9.143482, 
    -9.017111, -8.890595, -8.763936, -8.637134, -8.510187, -8.3831, 
    -8.255868, -8.128495, -8.00098, -7.873324, -7.745526, -7.617588, 
    -7.489509, -7.36129, -7.232931, -7.104433, -6.975795, -6.847019, 
    -6.718105, -6.589052, -6.459862, -6.330535, -6.201071, -6.07147, 
    -5.941734, -5.811862, -5.681854, -5.551712, -5.421435, -5.291025, 
    -5.16048, -5.029804, -4.898993, -4.768052, -4.636978, -4.505773, 
    -4.374437, -4.242971, -4.111375, -3.979649, -3.847795, -3.715812, 
    -3.583701, -3.451462, -3.319097, -3.186605, -3.053988, -2.921244, 
    -2.788376, -2.655384, -2.522267, -2.389028, -2.255665, -2.122181, 
    -1.988574, -1.854847, -1.720999, -1.587031, -1.452944, -1.318738, 
    -1.184413, -1.049971, -0.915412, -0.7807364, -0.6459449, -0.5110382, 
    -0.3760168, -0.2408813, -0.1056325, 0.0297291, 0.1652029, 0.3007881, 
    0.4364843, 0.5722907, 0.7082066, 0.8442314, 0.9803645, 1.116605, 
    1.252953, 1.389407, 1.525966, 1.66263, 1.799399, 1.936271, 2.073245, 
    2.210322, 2.3475, 2.484779, 2.622158, 2.759636, 2.897212, 3.034886, 
    3.172657, 3.310525, 3.448488, 3.586546, 3.724698, 3.862943, 4.00128, 
    4.139709, 4.27823, 4.41684, 4.55554, 4.694329, 4.833205, 4.972168, 
    5.111217, 5.250353, 5.389572, 5.528876, 5.668262, 5.807731, 5.94728, 
    6.086911, 6.226621, 6.36641, 6.506277, 6.646222, 6.786242, 6.926338, 
    7.066509, 7.206753, 7.347071, 7.48746, 7.627921, 7.768452, 7.909052, 
    8.049721, 8.190457, 8.331261, 8.47213, 8.613064, 8.754063, 8.895123, 
    9.036247, 9.177433, 9.318679, 9.459984, 9.601348, 9.742769, 9.884248, 
    10.02578, 10.16737, 10.30902, 10.45071, 10.59246, 10.73426, 10.87611, 
    11.01801, 11.15996, 11.30195, 11.444, 11.58608, 11.72821, 11.87039, 
    12.01261, 12.15487, 12.29717, 12.43951, 12.58189, 12.72431, 12.86676, 
    13.00925, 13.15178, 13.29433, 13.43693, 13.57955, 13.72221, 13.86489, 
    14.0076, 14.15034, 14.29311, 14.43591, 14.57873, 14.72157, 14.86444, 
    15.00733, 15.15024, 15.29317, 15.43612, 15.57909, 15.72207, 15.86507, 
    16.00809, 16.15112, 16.29416, 16.43721, 16.58028, 16.72335, 16.86644, 
    17.00953, 17.15263, 17.29574, 17.43885, 17.58196, 17.72508, 17.8682, 
    18.01132, 18.15444, 18.29756, 18.44068, 18.58379, 18.7269, 18.87, 
    19.0131, 19.15619, 19.29928, 19.44235, 19.58542, 19.72847, 19.87151, 
    20.01454, 20.15755, 20.30055, 20.44353, 20.58649, 20.72944, 20.87237, 
    21.01528, 21.15816, 21.30103, 21.44386, 21.58668, 21.72947, 21.87224, 
    22.01497, 22.15768, 22.30036, 22.44301, 22.58563, 22.72822, 22.87077, 
    23.01329, 23.15578, 23.29822, 23.44064, 23.58301, 23.72534, 23.86764, 
    24.00989, 24.1521, 24.29427, 24.4364, 24.57848, 24.72051, 24.8625, 
    25.00444, 25.14633, 25.28817, 25.42997, 25.57171, 25.71339, 25.85503, 
    25.99661, 26.13814, 26.27961, 26.42102, 26.56237, 26.70367, 26.8449, 
    26.98608, 27.12719, 27.26825, 27.40923, 27.55016, 27.69102, 27.83181, 
    27.97254, 28.11319, 28.25378, 28.3943, 28.53475, 28.67513, 28.81544, 
    28.95567, 29.09583, 29.23591, 29.37592, 29.51585, 29.65571, 29.79548, 
    29.93518, 30.0748, 30.21434, 30.35379, 30.49317, 30.63246, 30.77166, 
    30.91078, 31.04982, 31.18877, 31.32763, 31.46641, 31.60509, 31.74369, 
    31.88219, 32.02061, 32.15893, 32.29716, 32.4353, 32.57334, 32.71129, 
    32.84914, 32.9869, 33.12456, 33.26212, 33.39958, 33.53694, 33.67421, 
    33.81137, 33.94843, 34.08539, 34.22224, 34.35899, 34.49564, 34.63219, 
    34.76862, 34.90495, 35.04118, 35.17729, 35.3133, 35.4492, 35.58499, 
    35.72066, 35.85624, 35.99169, 36.12703, 36.26226, 36.39738, 36.53239, 
    36.66727, 36.80205, 36.93671, 37.07125, 37.20567, 37.33997, 37.47416, 
    37.60823, 37.74218, 37.87601, 38.00972, 38.1433, 38.27677, 38.41011, 
    38.54333, 38.67643, 38.8094, 38.94225, 39.07497, 39.20757, 39.34004, 
    39.47239, 39.60461, 39.7367, 39.86866, 40.0005, 40.1322, 40.26377, 
    40.39522, 40.52654, 40.65772, 40.78877, 40.91969, 41.05048, 41.18114, 
    41.31166, 41.44205, 41.57231, 41.70243,
  -17.21508, -17.09849, -16.98174, -16.86485, -16.74779, -16.63059, 
    -16.51323, -16.39571, -16.27804, -16.16022, -16.04224, -15.92411, 
    -15.80583, -15.68739, -15.5688, -15.45005, -15.33115, -15.2121, 
    -15.09289, -14.97353, -14.85402, -14.73435, -14.61454, -14.49456, 
    -14.37444, -14.25416, -14.13373, -14.01314, -13.89241, -13.77152, 
    -13.65048, -13.52928, -13.40794, -13.28644, -13.16479, -13.04299, 
    -12.92103, -12.79893, -12.67667, -12.55427, -12.43171, -12.309, 
    -12.18614, -12.06313, -11.93997, -11.81666, -11.6932, -11.56959, 
    -11.44583, -11.32192, -11.19786, -11.07365, -10.9493, -10.82479, 
    -10.70014, -10.57534, -10.45039, -10.32529, -10.20005, -10.07466, 
    -9.94912, -9.823435, -9.697604, -9.571627, -9.445504, -9.319236, 
    -9.192822, -9.066262, -8.939559, -8.812711, -8.685719, -8.558583, 
    -8.431303, -8.303881, -8.176314, -8.048607, -7.920756, -7.792763, 
    -7.664629, -7.536354, -7.407938, -7.279381, -7.150684, -7.021847, 
    -6.89287, -6.763755, -6.634501, -6.505108, -6.375578, -6.24591, 
    -6.116105, -5.986163, -5.856084, -5.72587, -5.59552, -5.465034, 
    -5.334415, -5.203661, -5.072773, -4.941752, -4.810598, -4.679311, 
    -4.547892, -4.416342, -4.284661, -4.152849, -4.020906, -3.888835, 
    -3.756634, -3.624304, -3.491846, -3.359261, -3.226548, -3.093709, 
    -2.960743, -2.827652, -2.694435, -2.561095, -2.42763, -2.294041, 
    -2.16033, -2.026496, -1.892541, -1.758464, -1.624267, -1.489949, 
    -1.355512, -1.220956, -1.086282, -0.9514901, -0.8165809, -0.6815551, 
    -0.5464134, -0.4111564, -0.2757846, -0.1402988, -0.00469958, 0.1310125, 
    0.2668367, 0.4027725, 0.5388191, 0.6749761, 0.8112425, 0.9476178, 
    1.084101, 1.220693, 1.35739, 1.494195, 1.631104, 1.768119, 1.905237, 
    2.042459, 2.179784, 2.317211, 2.454739, 2.592367, 2.730095, 2.867923, 
    3.005849, 3.143872, 3.281992, 3.420208, 3.55852, 3.696927, 3.835427, 
    3.97402, 4.112705, 4.251482, 4.39035, 4.529308, 4.668355, 4.80749, 
    4.946712, 5.086022, 5.225418, 5.364898, 5.504463, 5.644112, 5.783843, 
    5.923656, 6.06355, 6.203524, 6.343578, 6.48371, 6.62392, 6.764206, 
    6.904569, 7.045007, 7.185519, 7.326104, 7.466762, 7.607491, 7.748291, 
    7.889162, 8.030101, 8.171107, 8.312181, 8.453322, 8.594528, 8.735799, 
    8.877133, 9.01853, 9.159988, 9.301508, 9.443088, 9.584726, 9.726422, 
    9.868176, 10.00999, 10.15185, 10.29377, 10.43574, 10.57777, 10.71985, 
    10.86198, 11.00415, 11.14638, 11.28865, 11.43097, 11.57334, 11.71575, 
    11.85821, 12.00071, 12.14325, 12.28583, 12.42845, 12.57111, 12.71381, 
    12.85654, 12.99932, 13.14212, 13.28496, 13.42784, 13.57074, 13.71368, 
    13.85665, 13.99965, 14.14267, 14.28572, 14.4288, 14.57191, 14.71503, 
    14.85818, 15.00136, 15.14455, 15.28777, 15.431, 15.57425, 15.71752, 
    15.86081, 16.00411, 16.14742, 16.29075, 16.43409, 16.57744, 16.7208, 
    16.86418, 17.00755, 17.15094, 17.29433, 17.43773, 17.58113, 17.72453, 
    17.86794, 18.01134, 18.15475, 18.29815, 18.44156, 18.58496, 18.72835, 
    18.87174, 19.01513, 19.1585, 19.30187, 19.44523, 19.58858, 19.73192, 
    19.87525, 20.01856, 20.16186, 20.30514, 20.44841, 20.59166, 20.73489, 
    20.8781, 21.02129, 21.16446, 21.30761, 21.45073, 21.59383, 21.73691, 
    21.87996, 22.02298, 22.16597, 22.30893, 22.45186, 22.59476, 22.73763, 
    22.88047, 23.02327, 23.16604, 23.30877, 23.45146, 23.59411, 23.73673, 
    23.8793, 24.02184, 24.16433, 24.30678, 24.44918, 24.59154, 24.73386, 
    24.87612, 25.01834, 25.16051, 25.30263, 25.4447, 25.58672, 25.72868, 
    25.87059, 26.01245, 26.15425, 26.296, 26.43768, 26.57931, 26.72088, 
    26.86239, 27.00384, 27.14523, 27.28655, 27.42781, 27.56901, 27.71014, 
    27.8512, 27.9922, 28.13313, 28.27398, 28.41477, 28.55549, 28.69614, 
    28.83671, 28.97721, 29.11764, 29.25799, 29.39826, 29.53846, 29.67858, 
    29.81862, 29.95858, 30.09846, 30.23827, 30.37798, 30.51762, 30.65717, 
    30.79664, 30.93602, 31.07532, 31.21453, 31.35365, 31.49268, 31.63162, 
    31.77048, 31.90924, 32.04791, 32.18649, 32.32497, 32.46336, 32.60166, 
    32.73986, 32.87797, 33.01598, 33.15388, 33.2917, 33.42941, 33.56702, 
    33.70454, 33.84195, 33.97926, 34.11646, 34.25356, 34.39056, 34.52745, 
    34.66424, 34.80092, 34.9375, 35.07396, 35.21032, 35.34657, 35.48271, 
    35.61874, 35.75466, 35.89046, 36.02616, 36.16174, 36.29721, 36.43256, 
    36.5678, 36.70292, 36.83793, 36.97282, 37.10759, 37.24225, 37.37679, 
    37.5112, 37.6455, 37.77968, 37.91374, 38.04768, 38.18149, 38.31518, 
    38.44875, 38.5822, 38.71552, 38.84871, 38.98178, 39.11473, 39.24755, 
    39.38024, 39.51281, 39.64524, 39.77755, 39.90974, 40.04179, 40.17371, 
    40.3055, 40.43716, 40.56869, 40.70009, 40.83135, 40.96249, 41.09349, 
    41.22435, 41.35509, 41.48568, 41.61615, 41.74648,
  -17.27527, -17.15854, -17.04166, -16.92462, -16.80743, -16.69008, 
    -16.57258, -16.45492, -16.33711, -16.21914, -16.10102, -15.98274, 
    -15.86431, -15.74572, -15.62698, -15.50809, -15.38904, -15.26984, 
    -15.15048, -15.03097, -14.91131, -14.79149, -14.67151, -14.55138, 
    -14.4311, -14.31067, -14.19008, -14.06934, -13.94845, -13.8274, -13.7062, 
    -13.58484, -13.46334, -13.34167, -13.21986, -13.0979, -12.97578, 
    -12.85351, -12.73109, -12.60852, -12.48579, -12.36291, -12.23989, 
    -12.11671, -11.99338, -11.86989, -11.74626, -11.62248, -11.49855, 
    -11.37446, -11.25023, -11.12585, -11.00132, -10.87663, -10.7518, 
    -10.62682, -10.5017, -10.37642, -10.25099, -10.12542, -9.999701, 
    -9.873834, -9.747819, -9.621657, -9.495349, -9.368895, -9.242294, 
    -9.115547, -8.988656, -8.861618, -8.734436, -8.60711, -8.479639, 
    -8.352024, -8.224265, -8.096363, -7.968318, -7.84013, -7.711801, 
    -7.583328, -7.454715, -7.32596, -7.197063, -7.068027, -6.93885, 
    -6.809533, -6.680077, -6.550482, -6.420748, -6.290875, -6.160865, 
    -6.030717, -5.900432, -5.77001, -5.639452, -5.508759, -5.377929, 
    -5.246964, -5.115866, -4.984632, -4.853266, -4.721766, -4.590133, 
    -4.458368, -4.326471, -4.194443, -4.062284, -3.929994, -3.797575, 
    -3.665026, -3.532348, -3.399542, -3.266608, -3.133546, -3.000358, 
    -2.867043, -2.733603, -2.600037, -2.466346, -2.332531, -2.198593, 
    -2.064531, -1.930347, -1.796041, -1.661614, -1.527066, -1.392397, 
    -1.257609, -1.122702, -0.9876768, -0.8525335, -0.7172729, -0.5818956, 
    -0.4464024, -0.3107938, -0.1750705, -0.03923299, 0.09671797, 0.2327818, 
    0.3689578, 0.5052453, 0.6416437, 0.7781523, 0.9147705, 1.051498, 
    1.188333, 1.325276, 1.462325, 1.599481, 1.736742, 1.874108, 2.011578, 
    2.149151, 2.286827, 2.424605, 2.562484, 2.700463, 2.838542, 2.97672, 
    3.114996, 3.25337, 3.39184, 3.530406, 3.669068, 3.807824, 3.946673, 
    4.085616, 4.22465, 4.363776, 4.502992, 4.642298, 4.781693, 4.921176, 
    5.060746, 5.200403, 5.340146, 5.479973, 5.619884, 5.759879, 5.899956, 
    6.040114, 6.180353, 6.320673, 6.461071, 6.601547, 6.7421, 6.88273, 
    7.023436, 7.164216, 7.305069, 7.445997, 7.586996, 7.728066, 7.869206, 
    8.010416, 8.151695, 8.293041, 8.434454, 8.575933, 8.717476, 8.859084, 
    9.000754, 9.142488, 9.284282, 9.426136, 9.568049, 9.710022, 9.852052, 
    9.994139, 10.13628, 10.27848, 10.42073, 10.56303, 10.70539, 10.84779, 
    10.99025, 11.13276, 11.27531, 11.41791, 11.56056, 11.70325, 11.84598, 
    11.98876, 12.13159, 12.27445, 12.41735, 12.56029, 12.70327, 12.84629, 
    12.98935, 13.13244, 13.27556, 13.41872, 13.56191, 13.70513, 13.84838, 
    13.99166, 14.13497, 14.27831, 14.42167, 14.56506, 14.70847, 14.85191, 
    14.99537, 15.13885, 15.28235, 15.42587, 15.56941, 15.71296, 15.85653, 
    16.00012, 16.14372, 16.28734, 16.43096, 16.5746, 16.71825, 16.8619, 
    17.00557, 17.14924, 17.29292, 17.4366, 17.58029, 17.72398, 17.86767, 
    18.01137, 18.15506, 18.29875, 18.44244, 18.58613, 18.72981, 18.87349, 
    19.01716, 19.16082, 19.30448, 19.44812, 19.59176, 19.73538, 19.879, 
    20.02259, 20.16618, 20.30975, 20.4533, 20.59683, 20.74035, 20.88385, 
    21.02733, 21.17078, 21.31421, 21.45762, 21.60101, 21.74437, 21.8877, 
    22.031, 22.17428, 22.31753, 22.46074, 22.60393, 22.74708, 22.8902, 
    23.03329, 23.17633, 23.31935, 23.46232, 23.60526, 23.74815, 23.89101, 
    24.03382, 24.1766, 24.31933, 24.46201, 24.60465, 24.74724, 24.88979, 
    25.03229, 25.17474, 25.31713, 25.45948, 25.60178, 25.74402, 25.88621, 
    26.02834, 26.17042, 26.31244, 26.4544, 26.59631, 26.73815, 26.87994, 
    27.02166, 27.16332, 27.30492, 27.44645, 27.58792, 27.72932, 27.87066, 
    28.01192, 28.15312, 28.29425, 28.43531, 28.5763, 28.71722, 28.85806, 
    28.99883, 29.13952, 29.28014, 29.42068, 29.56114, 29.70153, 29.84184, 
    29.98206, 30.12221, 30.26227, 30.40225, 30.54215, 30.68196, 30.82169, 
    30.96134, 31.10089, 31.24036, 31.37974, 31.51904, 31.65824, 31.79735, 
    31.93637, 32.0753, 32.21413, 32.35287, 32.49152, 32.63007, 32.76852, 
    32.90688, 33.04514, 33.18331, 33.32137, 33.45933, 33.59719, 33.73496, 
    33.87262, 34.01017, 34.14763, 34.28498, 34.42222, 34.55936, 34.69639, 
    34.83332, 34.97014, 35.10685, 35.24345, 35.37994, 35.51632, 35.65259, 
    35.78875, 35.92479, 36.06073, 36.19655, 36.33225, 36.46784, 36.60332, 
    36.73868, 36.87392, 37.00904, 37.14405, 37.27894, 37.41371, 37.54836, 
    37.68289, 37.8173, 37.95158, 38.08575, 38.21979, 38.35371, 38.4875, 
    38.62117, 38.75472, 38.88814, 39.02143, 39.1546, 39.28764, 39.42056, 
    39.55334, 39.686, 39.81853, 39.95093, 40.0832, 40.21534, 40.34734, 
    40.47922, 40.61097, 40.74258, 40.87405, 41.0054, 41.13661, 41.26769, 
    41.39863, 41.52944, 41.66011, 41.79065,
  -17.33561, -17.21874, -17.10172, -16.98454, -16.8672, -16.74971, -16.63207, 
    -16.51427, -16.39631, -16.2782, -16.15993, -16.04151, -15.92293, 
    -15.8042, -15.68531, -15.56627, -15.44707, -15.32772, -15.20821, 
    -15.08855, -14.96873, -14.84876, -14.72863, -14.60835, -14.48791, 
    -14.36732, -14.24658, -14.12568, -14.00462, -13.88342, -13.76206, 
    -13.64054, -13.51887, -13.39705, -13.27507, -13.15295, -13.03067, 
    -12.90823, -12.78564, -12.6629, -12.54001, -12.41697, -12.29377, 
    -12.17042, -12.04692, -11.92327, -11.79946, -11.67551, -11.5514, 
    -11.42715, -11.30274, -11.17818, -11.05347, -10.92861, -10.8036, 
    -10.67844, -10.55314, -10.42768, -10.30208, -10.17632, -10.05042, 
    -9.924368, -9.798169, -9.671823, -9.545329, -9.418688, -9.291901, 
    -9.164966, -9.037886, -8.910659, -8.783287, -8.655769, -8.528107, 
    -8.400299, -8.272347, -8.144252, -8.016012, -7.887629, -7.759102, 
    -7.630433, -7.501622, -7.372668, -7.243573, -7.114336, -6.984958, 
    -6.85544, -6.725781, -6.595983, -6.466045, -6.335968, -6.205752, 
    -6.075398, -5.944906, -5.814277, -5.68351, -5.552607, -5.421567, 
    -5.290392, -5.159082, -5.027637, -4.896057, -4.764344, -4.632496, 
    -4.500516, -4.368403, -4.236158, -4.103782, -3.971274, -3.838636, 
    -3.705867, -3.572969, -3.439941, -3.306785, -3.173501, -3.04009, 
    -2.906551, -2.772886, -2.639094, -2.505177, -2.371136, -2.23697, 
    -2.10268, -1.968267, -1.833731, -1.699073, -1.564294, -1.429393, 
    -1.294373, -1.159232, -1.023973, -0.8885949, -0.7530989, -0.6174856, 
    -0.4817556, -0.3459096, -0.2099481, -0.07387184, 0.0623186, 0.1986226, 
    0.3350393, 0.4715684, 0.608209, 0.7449604, 0.881822, 1.018793, 1.155873, 
    1.293061, 1.430357, 1.56776, 1.705268, 1.842882, 1.9806, 2.118423, 
    2.256349, 2.394377, 2.532507, 2.670738, 2.809069, 2.9475, 3.08603, 
    3.224658, 3.363383, 3.502204, 3.641121, 3.780134, 3.91924, 4.05844, 
    4.197733, 4.337117, 4.476593, 4.616159, 4.755814, 4.895558, 5.03539, 
    5.175309, 5.315314, 5.455404, 5.595579, 5.735838, 5.876179, 6.016603, 
    6.157108, 6.297693, 6.438358, 6.579101, 6.719922, 6.86082, 7.001794, 
    7.142844, 7.283967, 7.425164, 7.566433, 7.707775, 7.849186, 7.990668, 
    8.132219, 8.273838, 8.415524, 8.557276, 8.699094, 8.840976, 8.982921, 
    9.124928, 9.266998, 9.409129, 9.551319, 9.693568, 9.835875, 9.978239, 
    10.12066, 10.26313, 10.40566, 10.54825, 10.69088, 10.83357, 10.9763, 
    11.11909, 11.26192, 11.4048, 11.54773, 11.6907, 11.83372, 11.97678, 
    12.11989, 12.26303, 12.40622, 12.54944, 12.69271, 12.83601, 12.97935, 
    13.12272, 13.26613, 13.40957, 13.55304, 13.69655, 13.84009, 13.98365, 
    14.12725, 14.27087, 14.41452, 14.55819, 14.70189, 14.84561, 14.98936, 
    15.13313, 15.27691, 15.42072, 15.56454, 15.70839, 15.85224, 15.99612, 
    16.14001, 16.28391, 16.42782, 16.57174, 16.71568, 16.85962, 17.00358, 
    17.14754, 17.2915, 17.43547, 17.57945, 17.72343, 17.86741, 18.01139, 
    18.15537, 18.29935, 18.44333, 18.5873, 18.73127, 18.87523, 19.01919, 
    19.16315, 19.30709, 19.45102, 19.59494, 19.73886, 19.88276, 20.02664, 
    20.17051, 20.31437, 20.45821, 20.60203, 20.74583, 20.88962, 21.03338, 
    21.17712, 21.32084, 21.46454, 21.60821, 21.75185, 21.89547, 22.03906, 
    22.18262, 22.32615, 22.46965, 22.61312, 22.75656, 22.89996, 23.04333, 
    23.18666, 23.32996, 23.47322, 23.61644, 23.75961, 23.90275, 24.04585, 
    24.18891, 24.33192, 24.47488, 24.6178, 24.76068, 24.9035, 25.04628, 
    25.18901, 25.33169, 25.47431, 25.61689, 25.75941, 25.90187, 26.04428, 
    26.18664, 26.32894, 26.47118, 26.61336, 26.75548, 26.89754, 27.03954, 
    27.18147, 27.32334, 27.46515, 27.60689, 27.74857, 27.89018, 28.03172, 
    28.17319, 28.31459, 28.45592, 28.59718, 28.73836, 28.87947, 29.02051, 
    29.16147, 29.30236, 29.44317, 29.5839, 29.72455, 29.86512, 30.00562, 
    30.14603, 30.28635, 30.4266, 30.56676, 30.70684, 30.84683, 30.98673, 
    31.12655, 31.26628, 31.40592, 31.54548, 31.68494, 31.82431, 31.96358, 
    32.10277, 32.24186, 32.38086, 32.51976, 32.65857, 32.79728, 32.93589, 
    33.07441, 33.21282, 33.35114, 33.48935, 33.62746, 33.76548, 33.90339, 
    34.04119, 34.17889, 34.31649, 34.45398, 34.59137, 34.72865, 34.86582, 
    35.00288, 35.13984, 35.27668, 35.41341, 35.55004, 35.68655, 35.82294, 
    35.95923, 36.09541, 36.23146, 36.3674, 36.50323, 36.63895, 36.77454, 
    36.91002, 37.04538, 37.18062, 37.31574, 37.45074, 37.58562, 37.72038, 
    37.85502, 37.98954, 38.12393, 38.2582, 38.39235, 38.52637, 38.66027, 
    38.79404, 38.92768, 39.0612, 39.19459, 39.32786, 39.46099, 39.594, 
    39.72688, 39.85963, 39.99224, 40.12473, 40.25709, 40.38931, 40.5214, 
    40.65336, 40.78519, 40.91688, 41.04844, 41.17986, 41.31115, 41.44231, 
    41.57332, 41.7042, 41.83495,
  -17.39608, -17.27908, -17.16191, -17.04459, -16.92712, -16.80949, -16.6917, 
    -16.57376, -16.45566, -16.3374, -16.21899, -16.10042, -15.9817, 
    -15.86281, -15.74378, -15.62459, -15.50524, -15.38574, -15.26608, 
    -15.14626, -15.02629, -14.90617, -14.78589, -14.66545, -14.54486, 
    -14.42411, -14.30321, -14.18215, -14.06094, -13.93958, -13.81806, 
    -13.69638, -13.57455, -13.45257, -13.33043, -13.20814, -13.08569, 
    -12.96309, -12.84034, -12.71743, -12.59437, -12.47116, -12.34779, 
    -12.22427, -12.1006, -11.97678, -11.8528, -11.72868, -11.6044, -11.47997, 
    -11.35538, -11.23065, -11.10576, -10.98073, -10.85554, -10.7302, 
    -10.60472, -10.47908, -10.35329, -10.22736, -10.10127, -9.975038, 
    -9.848655, -9.722123, -9.595444, -9.468616, -9.341641, -9.214519, 
    -9.08725, -8.959833, -8.832271, -8.704562, -8.576708, -8.448708, 
    -8.320562, -8.192272, -8.063837, -7.935258, -7.806536, -7.677669, 
    -7.548659, -7.419507, -7.290212, -7.160775, -7.031196, -6.901475, 
    -6.771615, -6.641613, -6.51147, -6.381188, -6.250767, -6.120206, 
    -5.989507, -5.858669, -5.727694, -5.596581, -5.465332, -5.333946, 
    -5.202424, -5.070765, -4.938972, -4.807045, -4.674983, -4.542787, 
    -4.410458, -4.277996, -4.145401, -4.012675, -3.879817, -3.746828, 
    -3.613709, -3.48046, -3.347082, -3.213575, -3.079939, -2.946176, 
    -2.812285, -2.678268, -2.544125, -2.409855, -2.275461, -2.140943, 
    -2.0063, -1.871534, -1.736645, -1.601634, -1.466501, -1.331247, 
    -1.195873, -1.060379, -0.9247658, -0.7890339, -0.653184, -0.5172167, 
    -0.3811327, -0.2449325, -0.1086168, 0.02781367, 0.1643583, 0.3010166, 
    0.4377877, 0.574671, 0.7116658, 0.8487716, 0.9859875, 1.123313, 1.260747, 
    1.398289, 1.535939, 1.673696, 1.811558, 1.949526, 2.087598, 2.225775, 
    2.364054, 2.502436, 2.640919, 2.779504, 2.918188, 3.056972, 3.195854, 
    3.334835, 3.473912, 3.613086, 3.752356, 3.89172, 4.031178, 4.17073, 
    4.310374, 4.450109, 4.589936, 4.729852, 4.869858, 5.009952, 5.150134, 
    5.290402, 5.430756, 5.571196, 5.71172, 5.852326, 5.993016, 6.133787, 
    6.27464, 6.415572, 6.556583, 6.697672, 6.83884, 6.980083, 7.121402, 
    7.262796, 7.404263, 7.545805, 7.687418, 7.829102, 7.970856, 8.112679, 
    8.254572, 8.396532, 8.538558, 8.680651, 8.822807, 8.965029, 9.107313, 
    9.249659, 9.392066, 9.534534, 9.67706, 9.819645, 9.962287, 10.10499, 
    10.24774, 10.39055, 10.53341, 10.67632, 10.81929, 10.96231, 11.10537, 
    11.24849, 11.39165, 11.53486, 11.67812, 11.82142, 11.96476, 12.10815, 
    12.25158, 12.39504, 12.53855, 12.6821, 12.82569, 12.96931, 13.11297, 
    13.25666, 13.40039, 13.54415, 13.68794, 13.83176, 13.97561, 14.1195, 
    14.2634, 14.40734, 14.5513, 14.69529, 14.8393, 14.98333, 15.12738, 
    15.27146, 15.41555, 15.55966, 15.70379, 15.84794, 15.9921, 16.13628, 
    16.28047, 16.42467, 16.56888, 16.71311, 16.85734, 17.00158, 17.14583, 
    17.29008, 17.43434, 17.57861, 17.72287, 17.86714, 18.01141, 18.15568, 
    18.29995, 18.44421, 18.58848, 18.73274, 18.87699, 19.02124, 19.16548, 
    19.30971, 19.45393, 19.59814, 19.74234, 19.88653, 20.0307, 20.17486, 
    20.31901, 20.46313, 20.60724, 20.75134, 20.89541, 21.03946, 21.18349, 
    21.32749, 21.47147, 21.61543, 21.75936, 21.90326, 22.04714, 22.19099, 
    22.33481, 22.47859, 22.62235, 22.76607, 22.90976, 23.05341, 23.19703, 
    23.34061, 23.48415, 23.62765, 23.77112, 23.91454, 24.05792, 24.20125, 
    24.34455, 24.48779, 24.631, 24.77415, 24.91726, 25.06032, 25.20333, 
    25.34629, 25.48919, 25.63205, 25.77485, 25.91759, 26.06028, 26.20291, 
    26.34549, 26.48801, 26.63046, 26.77286, 26.9152, 27.05747, 27.19968, 
    27.34183, 27.48391, 27.62593, 27.76788, 27.90976, 28.05157, 28.19332, 
    28.33499, 28.47659, 28.61812, 28.75957, 28.90096, 29.04226, 29.1835, 
    29.32465, 29.46573, 29.60673, 29.74765, 29.88849, 30.02925, 30.16992, 
    30.31051, 30.45103, 30.59145, 30.73179, 30.87205, 31.01221, 31.15229, 
    31.29229, 31.43219, 31.572, 31.71172, 31.85135, 31.99089, 32.13033, 
    32.26968, 32.40894, 32.5481, 32.68716, 32.82612, 32.96499, 33.10376, 
    33.24242, 33.38099, 33.51946, 33.65783, 33.79609, 33.93425, 34.0723, 
    34.21025, 34.3481, 34.48584, 34.62347, 34.761, 34.89842, 35.03572, 
    35.17292, 35.31001, 35.44699, 35.58385, 35.72061, 35.85725, 35.99377, 
    36.13019, 36.26648, 36.40267, 36.53873, 36.67468, 36.81051, 36.94622, 
    37.08182, 37.2173, 37.35265, 37.48788, 37.623, 37.75799, 37.89286, 
    38.02761, 38.16223, 38.29673, 38.4311, 38.56535, 38.69947, 38.83347, 
    38.96734, 39.10109, 39.2347, 39.36819, 39.50154, 39.63478, 39.76787, 
    39.90084, 40.03368, 40.16639, 40.29896, 40.4314, 40.56371, 40.69588, 
    40.82792, 40.95983, 41.0916, 41.22324, 41.35474, 41.4861, 41.61733, 
    41.74842, 41.87938,
  -17.4567, -17.33955, -17.22225, -17.10479, -16.98717, -16.8694, -16.75147, 
    -16.63338, -16.51514, -16.39674, -16.27818, -16.15947, -16.0406, 
    -15.92157, -15.80239, -15.68305, -15.56355, -15.4439, -15.32409, 
    -15.20412, -15.084, -14.96372, -14.84328, -14.72269, -14.60195, 
    -14.48104, -14.35998, -14.23877, -14.1174, -13.99588, -13.8742, 
    -13.75236, -13.63037, -13.50822, -13.38592, -13.26347, -13.14086, 
    -13.01809, -12.89517, -12.7721, -12.64887, -12.52549, -12.40196, 
    -12.27827, -12.15443, -12.03043, -11.90628, -11.78198, -11.65753, 
    -11.53292, -11.40816, -11.28326, -11.15819, -11.03298, -10.90762, 
    -10.7821, -10.65643, -10.53062, -10.40465, -10.27853, -10.15226, 
    -10.02584, -9.899276, -9.772559, -9.645694, -9.51868, -9.391518, 
    -9.264207, -9.136748, -9.009143, -8.88139, -8.753489, -8.625443, 
    -8.49725, -8.368911, -8.240426, -8.111795, -7.983021, -7.854101, 
    -7.725037, -7.595829, -7.466477, -7.336982, -7.207345, -7.077564, 
    -6.947642, -6.817577, -6.687372, -6.557025, -6.426538, -6.29591, 
    -6.165143, -6.034235, -5.90319, -5.772005, -5.640683, -5.509222, 
    -5.377625, -5.24589, -5.114019, -4.982012, -4.84987, -4.717593, 
    -4.585181, -4.452635, -4.319955, -4.187142, -4.054197, -3.921119, 
    -3.78791, -3.65457, -3.521099, -3.387498, -3.253767, -3.119907, 
    -2.985919, -2.851803, -2.717559, -2.583189, -2.448691, -2.314069, 
    -2.17932, -2.044448, -1.909451, -1.77433, -1.639087, -1.503721, 
    -1.368234, -1.232625, -1.096896, -0.9610471, -0.8250787, -0.6889916, 
    -0.5527864, -0.4164638, -0.2800243, -0.1434687, -0.006797541, 0.1299885, 
    0.2668887, 0.4039025, 0.5410292, 0.678268, 0.8156185, 0.9530797, 
    1.090651, 1.228332, 1.366122, 1.504019, 1.642025, 1.780136, 1.918354, 
    2.056677, 2.195104, 2.333636, 2.47227, 2.611006, 2.749844, 2.888783, 
    3.027822, 3.16696, 3.306196, 3.445531, 3.584962, 3.724489, 3.864112, 
    4.003829, 4.143641, 4.283545, 4.423541, 4.563629, 4.703807, 4.844075, 
    4.984432, 5.124877, 5.26541, 5.406029, 5.546733, 5.687523, 5.828396, 
    5.969352, 6.110391, 6.251511, 6.392711, 6.533991, 6.67535, 6.816787, 
    6.958301, 7.099891, 7.241556, 7.383295, 7.525108, 7.666994, 7.80895, 
    7.950978, 8.093076, 8.235243, 8.377478, 8.519779, 8.662147, 8.80458, 
    8.947078, 9.089639, 9.232262, 9.374947, 9.517692, 9.660497, 9.80336, 
    9.946281, 10.08926, 10.23229, 10.37538, 10.51853, 10.66172, 10.80497, 
    10.94827, 11.09161, 11.23501, 11.37846, 11.52195, 11.66549, 11.80907, 
    11.9527, 12.09637, 12.24008, 12.38384, 12.52763, 12.67146, 12.81533, 
    12.95924, 13.10319, 13.24716, 13.39118, 13.53522, 13.6793, 13.82341, 
    13.96755, 14.11172, 14.25591, 14.40014, 14.54439, 14.68866, 14.83296, 
    14.97728, 15.12162, 15.26598, 15.41037, 15.55477, 15.69919, 15.84362, 
    15.98807, 16.13254, 16.27702, 16.42151, 16.56601, 16.71052, 16.85505, 
    16.99957, 17.14411, 17.28866, 17.43321, 17.57776, 17.72232, 17.86687, 
    18.01143, 18.15599, 18.30055, 18.44511, 18.58966, 18.73421, 18.87875, 
    19.02329, 19.16782, 19.31234, 19.45685, 19.60135, 19.74584, 19.89032, 
    20.03478, 20.17923, 20.32366, 20.46808, 20.61247, 20.75686, 20.90121, 
    21.04555, 21.18987, 21.33416, 21.47843, 21.62268, 21.7669, 21.91109, 
    22.05525, 22.19939, 22.34349, 22.48756, 22.63161, 22.77561, 22.91959, 
    23.06352, 23.20743, 23.35129, 23.49512, 23.63891, 23.78265, 23.92636, 
    24.07002, 24.21364, 24.35722, 24.50075, 24.64424, 24.78768, 24.93106, 
    25.07441, 25.2177, 25.36094, 25.50412, 25.64725, 25.79034, 25.93336, 
    26.07633, 26.21924, 26.3621, 26.50489, 26.64763, 26.7903, 26.93292, 
    27.07547, 27.21795, 27.36038, 27.50274, 27.64503, 27.78725, 27.92941, 
    28.07149, 28.21351, 28.35546, 28.49733, 28.63913, 28.78086, 28.92251, 
    29.06409, 29.20559, 29.34702, 29.48836, 29.62963, 29.77082, 29.91192, 
    30.05295, 30.19389, 30.33475, 30.47553, 30.61622, 30.75683, 30.89734, 
    31.03778, 31.17812, 31.31837, 31.45854, 31.59861, 31.73859, 31.87848, 
    32.01828, 32.15798, 32.29759, 32.4371, 32.57652, 32.71584, 32.85506, 
    32.99418, 33.1332, 33.27213, 33.41095, 33.54967, 33.68829, 33.8268, 
    33.96521, 34.10352, 34.24172, 34.37981, 34.5178, 34.65568, 34.79345, 
    34.93112, 35.06867, 35.20612, 35.34345, 35.48067, 35.61778, 35.75478, 
    35.89165, 36.02842, 36.16508, 36.30161, 36.43803, 36.57434, 36.71053, 
    36.8466, 36.98254, 37.11837, 37.25409, 37.38968, 37.52514, 37.66049, 
    37.79571, 37.93081, 38.06579, 38.20065, 38.33537, 38.46997, 38.60445, 
    38.7388, 38.87303, 39.00712, 39.14109, 39.27493, 39.40864, 39.54222, 
    39.67567, 39.80899, 39.94218, 40.07524, 40.20816, 40.34095, 40.47361, 
    40.60614, 40.73853, 40.87078, 41.0029, 41.13489, 41.26674, 41.39845, 
    41.53003, 41.66146, 41.79277, 41.92393,
  -17.51745, -17.40017, -17.28273, -17.16513, -17.04737, -16.92946, 
    -16.81139, -16.69316, -16.57477, -16.45622, -16.33752, -16.21866, 
    -16.09965, -15.98047, -15.86114, -15.74165, -15.622, -15.5022, -15.38224, 
    -15.26212, -15.14184, -15.02141, -14.90082, -14.78008, -14.65918, 
    -14.53812, -14.4169, -14.29553, -14.174, -14.05232, -13.93048, -13.80848, 
    -13.68633, -13.56402, -13.44156, -13.31894, -13.19616, -13.07323, 
    -12.95015, -12.82691, -12.70351, -12.57996, -12.45626, -12.3324, 
    -12.20839, -12.08422, -11.9599, -11.83543, -11.7108, -11.58602, 
    -11.46109, -11.336, -11.21076, -11.08537, -10.95983, -10.83413, 
    -10.70829, -10.58229, -10.45614, -10.32984, -10.20339, -10.07679, 
    -9.950035, -9.823133, -9.696081, -9.56888, -9.44153, -9.314031, 
    -9.186383, -9.058587, -8.930643, -8.802551, -8.674313, -8.545926, 
    -8.417393, -8.288713, -8.159888, -8.030916, -7.9018, -7.772538, 
    -7.643131, -7.51358, -7.383885, -7.254046, -7.124064, -6.993939, 
    -6.863671, -6.733261, -6.602709, -6.472016, -6.341182, -6.210207, 
    -6.079093, -5.947838, -5.816444, -5.684911, -5.55324, -5.42143, 
    -5.289483, -5.157399, -5.025178, -4.89282, -4.760327, -4.627699, 
    -4.494936, -4.362038, -4.229007, -4.095842, -3.962544, -3.829114, 
    -3.695552, -3.561858, -3.428034, -3.29408, -3.159995, -3.025781, 
    -2.891439, -2.756968, -2.62237, -2.487644, -2.352792, -2.217814, 
    -2.082711, -1.947483, -1.81213, -1.676654, -1.541055, -1.405333, 
    -1.26949, -1.133525, -0.9974394, -0.8612339, -0.7249091, -0.5884655, 
    -0.4519036, -0.3152243, -0.1784281, -0.04151575, 0.09551219, 0.232655, 
    0.3699121, 0.5072827, 0.6447663, 0.782362, 0.9200693, 1.057887, 1.195816, 
    1.333853, 1.472, 1.610254, 1.748616, 1.887084, 2.025658, 2.164337, 
    2.303121, 2.442008, 2.580999, 2.720091, 2.859285, 2.998579, 3.137973, 
    3.277467, 3.417058, 3.556748, 3.696534, 3.836416, 3.976393, 4.116465, 
    4.256629, 4.396887, 4.537237, 4.677678, 4.81821, 4.95883, 5.09954, 
    5.240337, 5.381222, 5.522192, 5.663248, 5.804388, 5.945612, 6.086919, 
    6.228307, 6.369777, 6.511326, 6.652955, 6.794662, 6.936447, 7.078309, 
    7.220246, 7.362257, 7.504344, 7.646502, 7.788733, 7.931036, 8.073408, 
    8.21585, 8.35836, 8.500937, 8.643582, 8.786292, 8.929067, 9.071905, 
    9.214807, 9.35777, 9.500794, 9.643879, 9.787022, 9.930223, 10.07348, 
    10.2168, 10.36017, 10.50359, 10.64707, 10.7906, 10.93418, 11.07781, 
    11.22149, 11.36522, 11.50899, 11.65282, 11.79668, 11.9406, 12.08455, 
    12.22855, 12.37259, 12.51667, 12.66079, 12.80494, 12.94914, 13.09337, 
    13.23764, 13.38194, 13.52627, 13.67064, 13.81503, 13.95946, 14.10392, 
    14.2484, 14.39291, 14.53745, 14.68201, 14.8266, 14.97121, 15.11584, 
    15.26049, 15.40516, 15.54985, 15.69456, 15.83929, 15.98403, 16.12878, 
    16.27355, 16.41833, 16.56313, 16.70793, 16.85274, 16.99756, 17.14239, 
    17.28723, 17.43207, 17.57691, 17.72176, 17.86661, 18.01146, 18.15631, 
    18.30116, 18.446, 18.59085, 18.73568, 18.88052, 19.02534, 19.17016, 
    19.31498, 19.45978, 19.60457, 19.74935, 19.89412, 20.03887, 20.18361, 
    20.32833, 20.47304, 20.61772, 20.76239, 20.90704, 21.05167, 21.19628, 
    21.34086, 21.48542, 21.62995, 21.77446, 21.91894, 22.06339, 22.20781, 
    22.3522, 22.49656, 22.64089, 22.78519, 22.92945, 23.07367, 23.21786, 
    23.36201, 23.50612, 23.6502, 23.79423, 23.93822, 24.08217, 24.22608, 
    24.36994, 24.51375, 24.65752, 24.80124, 24.94491, 25.08854, 25.23211, 
    25.37563, 25.5191, 25.66252, 25.80588, 25.94918, 26.09243, 26.23562, 
    26.37876, 26.52183, 26.66485, 26.8078, 26.95069, 27.09352, 27.23629, 
    27.37899, 27.52162, 27.66419, 27.80669, 27.94912, 28.09148, 28.23377, 
    28.37599, 28.51814, 28.66021, 28.80221, 28.94414, 29.08599, 29.22776, 
    29.36945, 29.51107, 29.65261, 29.79406, 29.93544, 30.07673, 30.21794, 
    30.35907, 30.50011, 30.64107, 30.78194, 30.92272, 31.06342, 31.20403, 
    31.34454, 31.48497, 31.62531, 31.76555, 31.9057, 32.04576, 32.18572, 
    32.32558, 32.46535, 32.60503, 32.74461, 32.88408, 33.02346, 33.16274, 
    33.30192, 33.44099, 33.57997, 33.71884, 33.8576, 33.99627, 34.13483, 
    34.27328, 34.41162, 34.54986, 34.68799, 34.82601, 34.96392, 35.10172, 
    35.23941, 35.37699, 35.51445, 35.65181, 35.78905, 35.92617, 36.06318, 
    36.20007, 36.33685, 36.47351, 36.61006, 36.74648, 36.88279, 37.01897, 
    37.15504, 37.29099, 37.42681, 37.56251, 37.69809, 37.83355, 37.96888, 
    38.10409, 38.23917, 38.37413, 38.50896, 38.64367, 38.77825, 38.9127, 
    39.04702, 39.18121, 39.31528, 39.44921, 39.58302, 39.71669, 39.85023, 
    39.98364, 40.11692, 40.25006, 40.38307, 40.51595, 40.64869, 40.7813, 
    40.91376, 41.0461, 41.1783, 41.31036, 41.44229, 41.57408, 41.70573, 
    41.83724, 41.96861,
  -17.57835, -17.46093, -17.34335, -17.22561, -17.10771, -16.98966, 
    -16.87144, -16.75307, -16.63454, -16.51585, -16.397, -16.278, -16.15883, 
    -16.03951, -15.92003, -15.8004, -15.6806, -15.56064, -15.44053, 
    -15.32026, -15.19984, -15.07925, -14.95851, -14.83761, -14.71655, 
    -14.59533, -14.47396, -14.35243, -14.23075, -14.1089, -13.9869, 
    -13.86474, -13.74243, -13.61996, -13.49733, -13.37455, -13.25161, 
    -13.12851, -13.00526, -12.88186, -12.75829, -12.63458, -12.5107, 
    -12.38667, -12.26249, -12.13815, -12.01366, -11.88902, -11.76421, 
    -11.63926, -11.51415, -11.38889, -11.26347, -11.13791, -11.01218, 
    -10.88631, -10.76028, -10.6341, -10.50777, -10.38129, -10.25465, 
    -10.12787, -10.00093, -9.873844, -9.746606, -9.619218, -9.49168, 
    -9.363992, -9.236155, -9.108169, -8.980033, -8.851749, -8.723318, 
    -8.594738, -8.466011, -8.337136, -8.208115, -8.078947, -7.949633, 
    -7.820172, -7.690567, -7.560816, -7.43092, -7.30088, -7.170696, 
    -7.040368, -6.909896, -6.779282, -6.648525, -6.517626, -6.386585, 
    -6.255403, -6.124079, -5.992616, -5.861012, -5.729268, -5.597385, 
    -5.465364, -5.333203, -5.200905, -5.06847, -4.935897, -4.803188, 
    -4.670342, -4.537362, -4.404246, -4.270995, -4.13761, -4.004092, 
    -3.87044, -3.736656, -3.60274, -3.468692, -3.334512, -3.200203, 
    -3.065763, -2.931194, -2.796496, -2.661669, -2.526715, -2.391633, 
    -2.256425, -2.12109, -1.98563, -1.850045, -1.714336, -1.578502, 
    -1.442546, -1.306467, -1.170266, -1.033944, -0.8975005, -0.7609373, 
    -0.6242545, -0.487453, -0.3505332, -0.2134959, -0.0763417, 0.06092878, 
    0.1983148, 0.3358158, 0.4734311, 0.6111599, 0.7490016, 0.8869554, 
    1.025021, 1.163197, 1.301483, 1.439879, 1.578383, 1.716996, 1.855715, 
    1.994541, 2.133473, 2.27251, 2.411651, 2.550895, 2.690243, 2.829692, 
    2.969243, 3.108894, 3.248645, 3.388495, 3.528443, 3.668488, 3.80863, 
    3.948868, 4.0892, 4.229628, 4.370148, 4.51076, 4.651465, 4.79226, 
    4.933146, 5.07412, 5.215183, 5.356334, 5.497571, 5.638894, 5.780302, 
    5.921794, 6.06337, 6.205028, 6.346767, 6.488587, 6.630486, 6.772465, 
    6.914522, 7.056656, 7.198865, 7.341151, 7.48351, 7.625944, 7.768449, 
    7.911026, 8.053675, 8.196393, 8.339179, 8.482034, 8.624956, 8.767943, 
    8.910996, 9.054113, 9.197294, 9.340537, 9.483841, 9.627205, 9.770629, 
    9.914111, 10.05765, 10.20125, 10.3449, 10.48861, 10.63237, 10.77618, 
    10.92004, 11.06396, 11.20792, 11.35193, 11.496, 11.6401, 11.78426, 
    11.92845, 12.07269, 12.21698, 12.3613, 12.50567, 12.65008, 12.79452, 
    12.939, 13.08352, 13.22808, 13.37266, 13.51728, 13.66194, 13.80662, 
    13.95134, 14.09609, 14.24086, 14.38566, 14.53049, 14.67534, 14.82022, 
    14.96512, 15.11004, 15.25498, 15.39994, 15.54492, 15.68992, 15.83494, 
    15.97997, 16.12502, 16.27008, 16.41515, 16.56023, 16.70533, 16.85043, 
    16.99555, 17.14067, 17.28579, 17.43092, 17.57606, 17.7212, 17.86634, 
    18.01148, 18.15662, 18.30176, 18.4469, 18.59204, 18.73717, 18.88229, 
    19.02741, 19.17252, 19.31762, 19.46272, 19.6078, 19.75287, 19.89793, 
    20.04297, 20.188, 20.33302, 20.47801, 20.62299, 20.76795, 20.91289, 
    21.05781, 21.2027, 21.34757, 21.49242, 21.63725, 21.78204, 21.92681, 
    22.07155, 22.21626, 22.36094, 22.50559, 22.65021, 22.79479, 22.93934, 
    23.08385, 23.22833, 23.37277, 23.51717, 23.66153, 23.80585, 23.95012, 
    24.09436, 24.23855, 24.3827, 24.5268, 24.67085, 24.81485, 24.95881, 
    25.10272, 25.24657, 25.39038, 25.53413, 25.67783, 25.82147, 25.96506, 
    26.10859, 26.25206, 26.39548, 26.53883, 26.68213, 26.82536, 26.96853, 
    27.11164, 27.25468, 27.39766, 27.54057, 27.68341, 27.82619, 27.96889, 
    28.11153, 28.2541, 28.39659, 28.53901, 28.68136, 28.82364, 28.96583, 
    29.10795, 29.25, 29.39197, 29.53385, 29.67566, 29.81739, 29.95903, 
    30.10059, 30.24207, 30.38347, 30.52478, 30.666, 30.80714, 30.94818, 
    31.08915, 31.23002, 31.3708, 31.51149, 31.65209, 31.79259, 31.933, 
    32.07332, 32.21354, 32.35367, 32.4937, 32.63363, 32.77347, 32.9132, 
    33.05284, 33.19237, 33.33181, 33.47114, 33.61037, 33.74949, 33.88851, 
    34.02743, 34.16624, 34.30494, 34.44353, 34.58202, 34.7204, 34.85867, 
    34.99683, 35.13487, 35.27281, 35.41063, 35.54834, 35.68594, 35.82343, 
    35.96079, 36.09805, 36.23518, 36.3722, 36.5091, 36.64589, 36.78255, 
    36.91909, 37.05552, 37.19182, 37.328, 37.46406, 37.6, 37.73581, 37.8715, 
    38.00706, 38.14251, 38.27782, 38.41301, 38.54807, 38.68301, 38.81781, 
    38.95249, 39.08704, 39.22146, 39.35575, 39.48991, 39.62393, 39.75783, 
    39.89159, 40.02522, 40.15872, 40.29208, 40.42531, 40.55841, 40.69136, 
    40.82419, 40.95688, 41.08943, 41.22184, 41.35412, 41.48626, 41.61826, 
    41.75012, 41.88184, 42.01342,
  -17.6394, -17.52184, -17.40412, -17.28624, -17.1682, -17.05, -16.93164, 
    -16.81313, -16.69446, -16.57562, -16.45663, -16.33748, -16.21817, 
    -16.0987, -15.97907, -15.85928, -15.73934, -15.61923, -15.49897, 
    -15.37855, -15.25797, -15.13723, -15.01633, -14.89528, -14.77407, 
    -14.65269, -14.53117, -14.40948, -14.28763, -14.16563, -14.04347, 
    -13.92115, -13.79867, -13.67604, -13.55325, -13.4303, -13.3072, 
    -13.18394, -13.06052, -12.93695, -12.81322, -12.68933, -12.56529, 
    -12.44109, -12.31674, -12.19223, -12.06756, -11.94274, -11.81777, 
    -11.69264, -11.56736, -11.44192, -11.31632, -11.19058, -11.06468, 
    -10.93862, -10.81242, -10.68606, -10.55954, -10.43288, -10.30606, 
    -10.17909, -10.05197, -9.924694, -9.79727, -9.669694, -9.541967, 
    -9.41409, -9.286063, -9.157887, -9.02956, -8.901084, -8.77246, -8.643686, 
    -8.514765, -8.385695, -8.256477, -8.127112, -7.9976, -7.867941, 
    -7.738136, -7.608186, -7.478089, -7.347847, -7.21746, -7.086929, 
    -6.956254, -6.825435, -6.694472, -6.563366, -6.432118, -6.300728, 
    -6.169196, -6.037523, -5.905709, -5.773754, -5.641659, -5.509425, 
    -5.377051, -5.244539, -5.111888, -4.9791, -4.846174, -4.713112, 
    -4.579913, -4.446578, -4.313108, -4.179503, -4.045763, -3.91189, 
    -3.777883, -3.643743, -3.509471, -3.375067, -3.240531, -3.105865, 
    -2.971069, -2.836143, -2.701087, -2.565904, -2.430592, -2.295152, 
    -2.159586, -2.023894, -1.888076, -1.752132, -1.616065, -1.479873, 
    -1.343558, -1.20712, -1.07056, -0.933879, -0.7970768, -0.6601545, 
    -0.5231126, -0.3859518, -0.2486728, -0.1112761, 0.02623751, 0.1638674, 
    0.3016129, 0.4394734, 0.5774481, 0.7155363, 0.8537375, 0.9920508, 
    1.130476, 1.269011, 1.407657, 1.546412, 1.685275, 1.824247, 1.963325, 
    2.10251, 2.241801, 2.381196, 2.520696, 2.6603, 2.800005, 2.939813, 
    3.079722, 3.219731, 3.35984, 3.500047, 3.640353, 3.780755, 3.921254, 
    4.061849, 4.202538, 4.343321, 4.484198, 4.625166, 4.766226, 4.907377, 
    5.048617, 5.189947, 5.331364, 5.472869, 5.61446, 5.756137, 5.897898, 
    6.039743, 6.181671, 6.323681, 6.465773, 6.607944, 6.750195, 6.892524, 
    7.034931, 7.177415, 7.319974, 7.462609, 7.605317, 7.748098, 7.890952, 
    8.033876, 8.176871, 8.319935, 8.463068, 8.606268, 8.749534, 8.892866, 
    9.036263, 9.179723, 9.323246, 9.46683, 9.610476, 9.754182, 9.897945, 
    10.04177, 10.18565, 10.32958, 10.47357, 10.61761, 10.76171, 10.90586, 
    11.05006, 11.19431, 11.33861, 11.48295, 11.62735, 11.77179, 11.91627, 
    12.0608, 12.20537, 12.34998, 12.49464, 12.63933, 12.78406, 12.92883, 
    13.07364, 13.21848, 13.36336, 13.50827, 13.65321, 13.79819, 13.94319, 
    14.08823, 14.23329, 14.37839, 14.5235, 14.66865, 14.81381, 14.959, 
    15.10422, 15.24945, 15.3947, 15.53998, 15.68527, 15.83058, 15.9759, 
    16.12124, 16.26659, 16.41195, 16.55733, 16.70272, 16.84812, 16.99352, 
    17.13893, 17.28435, 17.42978, 17.5752, 17.72063, 17.86607, 18.0115, 
    18.15694, 18.30237, 18.4478, 18.59323, 18.73865, 18.88407, 19.02948, 
    19.17488, 19.32028, 19.46567, 19.61104, 19.7564, 19.90175, 20.04709, 
    20.19241, 20.33772, 20.483, 20.62827, 20.77353, 20.91875, 21.06396, 
    21.20915, 21.35431, 21.49945, 21.64457, 21.78966, 21.93471, 22.07974, 
    22.22475, 22.36972, 22.51466, 22.65956, 22.80443, 22.94927, 23.09407, 
    23.23884, 23.38356, 23.52825, 23.6729, 23.8175, 23.96207, 24.10659, 
    24.25107, 24.3955, 24.53988, 24.68422, 24.82851, 24.97276, 25.11695, 
    25.26109, 25.40517, 25.54921, 25.69319, 25.83712, 25.98099, 26.1248, 
    26.26855, 26.41225, 26.55589, 26.69946, 26.84297, 26.98643, 27.12981, 
    27.27313, 27.41639, 27.55958, 27.7027, 27.84575, 27.98874, 28.13165, 
    28.27449, 28.41726, 28.55996, 28.70258, 28.84513, 28.9876, 29.13, 
    29.27231, 29.41455, 29.55671, 29.69879, 29.84078, 29.9827, 30.12453, 
    30.26628, 30.40794, 30.54952, 30.69101, 30.83241, 30.97373, 31.11496, 
    31.25609, 31.39714, 31.53809, 31.67896, 31.81972, 31.9604, 32.10098, 
    32.24146, 32.38185, 32.52214, 32.66233, 32.80242, 32.94242, 33.08231, 
    33.2221, 33.36179, 33.50138, 33.64086, 33.78024, 33.91951, 34.05868, 
    34.19774, 34.3367, 34.47554, 34.61428, 34.75291, 34.89143, 35.02983, 
    35.16813, 35.30632, 35.44439, 35.58234, 35.72018, 35.85791, 35.99552, 
    36.13302, 36.2704, 36.40766, 36.5448, 36.68182, 36.81873, 36.95551, 
    37.09217, 37.22871, 37.36513, 37.50142, 37.6376, 37.77364, 37.90957, 
    38.04537, 38.18104, 38.31659, 38.452, 38.5873, 38.72246, 38.85749, 
    38.9924, 39.12717, 39.26182, 39.39634, 39.53072, 39.66497, 39.79909, 
    39.93307, 40.06693, 40.20065, 40.33423, 40.46768, 40.60099, 40.73417, 
    40.86721, 41.00011, 41.13288, 41.26551, 41.398, 41.53035, 41.66256, 
    41.79464, 41.92657, 42.05836,
  -17.70059, -17.58289, -17.46503, -17.34701, -17.22883, -17.11049, 
    -16.99199, -16.87333, -16.75451, -16.63554, -16.5164, -16.3971, 
    -16.27765, -16.15803, -16.03825, -15.91832, -15.79822, -15.67797, 
    -15.55755, -15.43698, -15.31625, -15.19536, -15.07431, -14.9531, 
    -14.83173, -14.7102, -14.58851, -14.46667, -14.34466, -14.2225, 
    -14.10018, -13.9777, -13.85506, -13.73227, -13.60932, -13.4862, 
    -13.36294, -13.23951, -13.11593, -12.99218, -12.86829, -12.74423, 
    -12.62002, -12.49565, -12.37113, -12.24645, -12.12161, -11.99661, 
    -11.87147, -11.74616, -11.6207, -11.49509, -11.36932, -11.24339, 
    -11.11731, -10.99108, -10.86469, -10.73815, -10.61145, -10.48461, 
    -10.3576, -10.23045, -10.10314, -9.975683, -9.848072, -9.720309, 
    -9.592394, -9.464328, -9.336111, -9.207744, -9.079225, -8.950557, 
    -8.821739, -8.692771, -8.563655, -8.434389, -8.304976, -8.175413, 
    -8.045703, -7.915846, -7.785841, -7.65569, -7.525393, -7.394948, 
    -7.264359, -7.133624, -7.002744, -6.87172, -6.740551, -6.60924, 
    -6.477784, -6.346185, -6.214444, -6.082561, -5.950536, -5.81837, 
    -5.686063, -5.553616, -5.421028, -5.288301, -5.155435, -5.022431, 
    -4.889288, -4.756008, -4.622591, -4.489037, -4.355346, -4.22152, 
    -4.087559, -3.953463, -3.819233, -3.68487, -3.550373, -3.415743, 
    -3.280982, -3.146089, -3.011065, -2.87591, -2.740626, -2.605212, 
    -2.469669, -2.333999, -2.1982, -2.062275, -1.926223, -1.790045, 
    -1.653742, -1.517315, -1.380763, -1.244088, -1.10729, -0.9703702, 
    -0.8333285, -0.696166, -0.5588832, -0.4214808, -0.2839594, -0.1463197, 
    -0.00856236, 0.129312, 0.2673026, 0.4054089, 0.5436301, 0.6819656, 
    0.8204146, 0.9589765, 1.097651, 1.236436, 1.375332, 1.514338, 1.653454, 
    1.792678, 1.93201, 2.071449, 2.210994, 2.350645, 2.4904, 2.63026, 
    2.770223, 2.910288, 3.050456, 3.190724, 3.331092, 3.47156, 3.612126, 
    3.75279, 3.893551, 4.034408, 4.175361, 4.316408, 4.457548, 4.598782, 
    4.740108, 4.881524, 5.023031, 5.164628, 5.306313, 5.448086, 5.589946, 
    5.731893, 5.873924, 6.016039, 6.158238, 6.30052, 6.442883, 6.585327, 
    6.727851, 6.870454, 7.013135, 7.155893, 7.298728, 7.441638, 7.584621, 
    7.727679, 7.87081, 8.014011, 8.157284, 8.300627, 8.444037, 8.587517, 
    8.731063, 8.874675, 9.018352, 9.162093, 9.305897, 9.449763, 9.593691, 
    9.737679, 9.881725, 10.02583, 10.16999, 10.31421, 10.45849, 10.60281, 
    10.7472, 10.89163, 11.03611, 11.18065, 11.32523, 11.46987, 11.61455, 
    11.75927, 11.90404, 12.04886, 12.19372, 12.33862, 12.48356, 12.62854, 
    12.77357, 12.91863, 13.06372, 13.20885, 13.35402, 13.49922, 13.64446, 
    13.78972, 13.93502, 14.08035, 14.2257, 14.37109, 14.51649, 14.66193, 
    14.80739, 14.95287, 15.09838, 15.2439, 15.38945, 15.53501, 15.6806, 
    15.8262, 15.97182, 16.11745, 16.26309, 16.40875, 16.55442, 16.7001, 
    16.84579, 16.99149, 17.1372, 17.28291, 17.42863, 17.57435, 17.72007, 
    17.8658, 18.01153, 18.15725, 18.30298, 18.44871, 18.59443, 18.74014, 
    18.88585, 19.03156, 19.17726, 19.32294, 19.46862, 19.61429, 19.75995, 
    19.90559, 20.05122, 20.19683, 20.34243, 20.48801, 20.63358, 20.77912, 
    20.92464, 21.07014, 21.21562, 21.36108, 21.50651, 21.65191, 21.79729, 
    21.94264, 22.08797, 22.23326, 22.37852, 22.52375, 22.66894, 22.8141, 
    22.95923, 23.10432, 23.24938, 23.39439, 23.53937, 23.6843, 23.8292, 
    23.97405, 24.11886, 24.26362, 24.40834, 24.55301, 24.69764, 24.84222, 
    24.98675, 25.13122, 25.27565, 25.42002, 25.56434, 25.7086, 25.85282, 
    25.99697, 26.14106, 26.2851, 26.42908, 26.573, 26.71685, 26.86065, 
    27.00438, 27.14805, 27.29165, 27.43518, 27.57865, 27.72205, 27.86539, 
    28.00865, 28.15184, 28.29495, 28.438, 28.58097, 28.72387, 28.86669, 
    29.00944, 29.15211, 29.2947, 29.43721, 29.57964, 29.72199, 29.86426, 
    30.00645, 30.14855, 30.29057, 30.4325, 30.57435, 30.7161, 30.85778, 
    30.99936, 31.14085, 31.28226, 31.42356, 31.56479, 31.70591, 31.84694, 
    31.98788, 32.12872, 32.26947, 32.41011, 32.55067, 32.69112, 32.83147, 
    32.97172, 33.11187, 33.25192, 33.39187, 33.53172, 33.67145, 33.81109, 
    33.95061, 34.09004, 34.22935, 34.36856, 34.50766, 34.64664, 34.78553, 
    34.92429, 35.06295, 35.20149, 35.33992, 35.47824, 35.61644, 35.75453, 
    35.89251, 36.03036, 36.1681, 36.30572, 36.44322, 36.58061, 36.71787, 
    36.85501, 36.99204, 37.12894, 37.26572, 37.40237, 37.5389, 37.67531, 
    37.8116, 37.94775, 38.08379, 38.21969, 38.35547, 38.49112, 38.62664, 
    38.76204, 38.8973, 39.03243, 39.16743, 39.30231, 39.43705, 39.57166, 
    39.70613, 39.84048, 39.97469, 40.10876, 40.2427, 40.3765, 40.51017, 
    40.6437, 40.7771, 40.91036, 41.04348, 41.17646, 41.30931, 41.44201, 
    41.57458, 41.707, 41.83929, 41.97143, 42.10343,
  -17.76192, -17.64408, -17.52608, -17.40792, -17.2896, -17.17112, -17.05248, 
    -16.93368, -16.81472, -16.6956, -16.57631, -16.45687, -16.33727, 
    -16.2175, -16.09758, -15.9775, -15.85725, -15.73685, -15.61628, 
    -15.49556, -15.37467, -15.25363, -15.13242, -15.01106, -14.88953, 
    -14.76785, -14.64601, -14.524, -14.40184, -14.27952, -14.15704, -14.0344, 
    -13.9116, -13.78864, -13.66552, -13.54225, -13.41881, -13.29522, 
    -13.17147, -13.04756, -12.9235, -12.79927, -12.67489, -12.55035, 
    -12.42566, -12.30081, -12.1758, -12.05063, -11.92531, -11.79983, 
    -11.67419, -11.5484, -11.42245, -11.29635, -11.17009, -11.04368, 
    -10.91711, -10.79039, -10.66351, -10.53648, -10.40929, -10.28195, 
    -10.15446, -10.02681, -9.899015, -9.771064, -9.642961, -9.514705, 
    -9.386297, -9.257739, -9.129028, -9.000168, -8.871157, -8.741995, 
    -8.612683, -8.483222, -8.353611, -8.223851, -8.093944, -7.963887, 
    -7.833682, -7.70333, -7.572831, -7.442185, -7.311392, -7.180454, 
    -7.049369, -6.918139, -6.786765, -6.655245, -6.523582, -6.391775, 
    -6.259824, -6.12773, -5.995494, -5.863117, -5.730597, -5.597936, 
    -5.465135, -5.332193, -5.199111, -5.06589, -4.93253, -4.799032, 
    -4.665395, -4.531621, -4.397711, -4.263664, -4.12948, -3.995162, 
    -3.860708, -3.72612, -3.591398, -3.456543, -3.321555, -3.186434, 
    -3.051182, -2.915798, -2.780284, -2.64464, -2.508866, -2.372964, 
    -2.236933, -2.100774, -1.964488, -1.828075, -1.691537, -1.554873, 
    -1.418084, -1.281171, -1.144134, -1.006975, -0.8696932, -0.7322899, 
    -0.5947656, -0.457121, -0.3193567, -0.1814733, -0.04347157, 0.09464783, 
    0.2328842, 0.371237, 0.5097054, 0.6482887, 0.7869862, 0.9257973, 
    1.064721, 1.203757, 1.342905, 1.482163, 1.621531, 1.761008, 1.900594, 
    2.040288, 2.180088, 2.319995, 2.460007, 2.600124, 2.740345, 2.880668, 
    3.021095, 3.161623, 3.302251, 3.44298, 3.583807, 3.724734, 3.865757, 
    4.006878, 4.148094, 4.289406, 4.430812, 4.572311, 4.713903, 4.855587, 
    4.997361, 5.139226, 5.28118, 5.423222, 5.565351, 5.707568, 5.84987, 
    5.992257, 6.134727, 6.277282, 6.419918, 6.562635, 6.705433, 6.84831, 
    6.991266, 7.1343, 7.27741, 7.420596, 7.563857, 7.707192, 7.8506, 
    7.994081, 8.137631, 8.281253, 8.424944, 8.568703, 8.712529, 8.856422, 
    9.000381, 9.144403, 9.288489, 9.432638, 9.576849, 9.72112, 9.865451, 
    10.00984, 10.15429, 10.29879, 10.44335, 10.58796, 10.73263, 10.87735, 
    11.02212, 11.16694, 11.31182, 11.45674, 11.6017, 11.74672, 11.89178, 
    12.03688, 12.18203, 12.32722, 12.47245, 12.61772, 12.76304, 12.90839, 
    13.05377, 13.1992, 13.34465, 13.49015, 13.63567, 13.78123, 13.92682, 
    14.07244, 14.21808, 14.36376, 14.50946, 14.65519, 14.80094, 14.94672, 
    15.09251, 15.23833, 15.38417, 15.53003, 15.67591, 15.82181, 15.96772, 
    16.11364, 16.25958, 16.40553, 16.5515, 16.69747, 16.84346, 16.98945, 
    17.13545, 17.28146, 17.42747, 17.57349, 17.71951, 17.86553, 18.01155, 
    18.15757, 18.30359, 18.44961, 18.59563, 18.74164, 18.88765, 19.03364, 
    19.17964, 19.32562, 19.47159, 19.61756, 19.76351, 19.90944, 20.05537, 
    20.20127, 20.34717, 20.49304, 20.6389, 20.78473, 20.93055, 21.07634, 
    21.22212, 21.36786, 21.51359, 21.65929, 21.80496, 21.9506, 22.09621, 
    22.2418, 22.38735, 22.53287, 22.67836, 22.82381, 22.96923, 23.11461, 
    23.25995, 23.40526, 23.55052, 23.69575, 23.84093, 23.98607, 24.13117, 
    24.27622, 24.42123, 24.56619, 24.71111, 24.85597, 25.00078, 25.14555, 
    25.29026, 25.43492, 25.57952, 25.72407, 25.86857, 26.013, 26.15738, 
    26.30171, 26.44597, 26.59017, 26.73431, 26.87838, 27.0224, 27.16634, 
    27.31023, 27.45404, 27.59779, 27.74147, 27.88508, 28.02862, 28.17209, 
    28.31549, 28.45881, 28.60206, 28.74523, 28.88833, 29.03135, 29.1743, 
    29.31716, 29.45995, 29.60265, 29.74527, 29.88781, 30.03027, 30.17265, 
    30.31493, 30.45714, 30.59925, 30.74128, 30.88322, 31.02507, 31.16683, 
    31.3085, 31.45008, 31.59156, 31.73295, 31.87425, 32.01545, 32.15656, 
    32.29757, 32.43848, 32.57929, 32.72, 32.86061, 33.00113, 33.14154, 
    33.28184, 33.42205, 33.56215, 33.70214, 33.84203, 33.98182, 34.12149, 
    34.26106, 34.40052, 34.53987, 34.67912, 34.81824, 34.95726, 35.09617, 
    35.23496, 35.37364, 35.51221, 35.65066, 35.78899, 35.92721, 36.06531, 
    36.20329, 36.34116, 36.4789, 36.61653, 36.75403, 36.89142, 37.02868, 
    37.16582, 37.30284, 37.43973, 37.5765, 37.71314, 37.84966, 37.98605, 
    38.12232, 38.25846, 38.39447, 38.53035, 38.66611, 38.80173, 38.93722, 
    39.07259, 39.20782, 39.34291, 39.47788, 39.61272, 39.74742, 39.88198, 
    40.01642, 40.15071, 40.28488, 40.4189, 40.55279, 40.68654, 40.82016, 
    40.95364, 41.08697, 41.22017, 41.35323, 41.48615, 41.61893, 41.75157, 
    41.88407, 42.01642, 42.14864,
  -17.8234, -17.70542, -17.58728, -17.46898, -17.35052, -17.2319, -17.11312, 
    -16.99418, -16.87507, -16.75581, -16.63638, -16.51679, -16.39704, 
    -16.27713, -16.15705, -16.03682, -15.91643, -15.79587, -15.67516, 
    -15.55428, -15.43324, -15.31204, -15.19069, -15.06917, -14.94749, 
    -14.82565, -14.70364, -14.58148, -14.45916, -14.33668, -14.21404, 
    -14.09124, -13.96828, -13.84516, -13.72188, -13.59844, -13.47484, 
    -13.35108, -13.22717, -13.10309, -12.97886, -12.85446, -12.72991, 
    -12.6052, -12.48034, -12.35531, -12.23013, -12.10479, -11.97929, 
    -11.85363, -11.72782, -11.60185, -11.47573, -11.34945, -11.22301, 
    -11.09642, -10.96967, -10.84276, -10.7157, -10.58849, -10.46112, 
    -10.3336, -10.20592, -10.07808, -9.950099, -9.821959, -9.693667, 
    -9.565222, -9.436625, -9.307874, -9.178972, -9.049918, -8.920713, 
    -8.791357, -8.66185, -8.532192, -8.402385, -8.272428, -8.142321, 
    -8.012065, -7.88166, -7.751107, -7.620406, -7.489557, -7.358561, 
    -7.227418, -7.096129, -6.964693, -6.833112, -6.701385, -6.569513, 
    -6.437497, -6.305336, -6.173033, -6.040585, -5.907995, -5.775262, 
    -5.642388, -5.509371, -5.376214, -5.242917, -5.109478, -4.975901, 
    -4.842184, -4.708328, -4.574334, -4.440202, -4.305933, -4.171528, 
    -4.036986, -3.902308, -3.767495, -3.632548, -3.497466, -3.362251, 
    -3.226902, -3.091422, -2.955809, -2.820064, -2.684189, -2.548184, 
    -2.412049, -2.275784, -2.139391, -2.002871, -1.866223, -1.729448, 
    -1.592547, -1.45552, -1.318369, -1.181093, -1.043694, -0.9061716, 
    -0.7685269, -0.6307605, -0.492873, -0.3548652, -0.2167376, -0.07849086, 
    0.05987422, 0.198357, 0.3369569, 0.475673, 0.6145048, 0.7534516, 
    0.8925126, 1.031687, 1.170974, 1.310374, 1.449885, 1.589506, 1.729237, 
    1.869078, 2.009026, 2.149083, 2.289246, 2.429515, 2.56989, 2.710369, 
    2.850952, 2.991638, 3.132427, 3.273316, 3.414307, 3.555397, 3.696586, 
    3.837873, 3.979258, 4.120739, 4.262316, 4.403988, 4.545753, 4.687613, 
    4.829564, 4.971607, 5.11374, 5.255963, 5.398275, 5.540676, 5.683163, 
    5.825737, 5.968396, 6.111139, 6.253966, 6.396876, 6.539868, 6.68294, 
    6.826093, 6.969325, 7.112634, 7.256021, 7.399485, 7.543023, 7.686636, 
    7.830323, 7.974082, 8.117913, 8.261815, 8.405786, 8.549826, 8.693933, 
    8.838108, 8.982348, 9.126655, 9.271024, 9.415456, 9.55995, 9.704505, 
    9.84912, 9.993794, 10.13853, 10.28332, 10.42816, 10.57306, 10.71801, 
    10.86302, 11.00808, 11.15319, 11.29835, 11.44356, 11.58882, 11.73412, 
    11.87947, 12.02486, 12.1703, 12.31578, 12.4613, 12.60687, 12.75247, 
    12.89811, 13.04379, 13.1895, 13.33525, 13.48104, 13.62686, 13.77271, 
    13.91859, 14.0645, 14.21044, 14.35641, 14.5024, 14.64843, 14.79447, 
    14.94054, 15.08663, 15.23275, 15.37888, 15.52504, 15.67121, 15.8174, 
    15.9636, 16.10982, 16.25606, 16.40231, 16.54856, 16.69484, 16.84112, 
    16.9874, 17.1337, 17.28, 17.42631, 17.57262, 17.71894, 17.86525, 
    18.01157, 18.15789, 18.30421, 18.45052, 18.59683, 18.74314, 18.88944, 
    19.03574, 19.18202, 19.3283, 19.47457, 19.62083, 19.76707, 19.91331, 
    20.05953, 20.20573, 20.35192, 20.49809, 20.64424, 20.79037, 20.93648, 
    21.08257, 21.22863, 21.37467, 21.52069, 21.66668, 21.81265, 21.95858, 
    22.10449, 22.25037, 22.39621, 22.54202, 22.6878, 22.83355, 22.97926, 
    23.12493, 23.27057, 23.41616, 23.56172, 23.70723, 23.85271, 23.99814, 
    24.14353, 24.28887, 24.43416, 24.57941, 24.72462, 24.86977, 25.01487, 
    25.15992, 25.30492, 25.44986, 25.59476, 25.73959, 25.88437, 26.02909, 
    26.17376, 26.31837, 26.46291, 26.6074, 26.75182, 26.89618, 27.04047, 
    27.1847, 27.32887, 27.47296, 27.61699, 27.76095, 27.90484, 28.04866, 
    28.19241, 28.33609, 28.47969, 28.62321, 28.76667, 28.91004, 29.05334, 
    29.19656, 29.3397, 29.48276, 29.62574, 29.76863, 29.91145, 30.05418, 
    30.19682, 30.33938, 30.48186, 30.62424, 30.76654, 30.90875, 31.05087, 
    31.1929, 31.33483, 31.47668, 31.61843, 31.76009, 31.90165, 32.04311, 
    32.18448, 32.32576, 32.46693, 32.608, 32.74898, 32.88985, 33.03062, 
    33.17129, 33.31186, 33.45232, 33.59268, 33.73293, 33.87308, 34.01312, 
    34.15305, 34.29287, 34.43259, 34.57219, 34.71169, 34.85107, 34.99034, 
    35.12949, 35.26854, 35.40746, 35.54628, 35.68497, 35.82355, 35.96202, 
    36.10037, 36.23859, 36.37671, 36.51469, 36.65256, 36.79031, 36.92793, 
    37.06544, 37.20282, 37.34007, 37.4772, 37.61421, 37.75109, 37.88785, 
    38.02448, 38.16098, 38.29735, 38.43359, 38.56971, 38.70569, 38.84155, 
    38.97727, 39.11286, 39.24832, 39.38365, 39.51884, 39.6539, 39.78883, 
    39.92362, 40.05828, 40.1928, 40.32718, 40.46143, 40.59554, 40.72951, 
    40.86335, 40.99704, 41.1306, 41.26401, 41.39729, 41.53042, 41.66341, 
    41.79627, 41.92898, 42.06155, 42.19397,
  -17.88503, -17.76691, -17.64863, -17.53019, -17.41159, -17.29283, 
    -17.17391, -17.05482, -16.93557, -16.81616, -16.69659, -16.57685, 
    -16.45696, -16.3369, -16.21668, -16.0963, -15.97575, -15.85505, 
    -15.73418, -15.61315, -15.49196, -15.37061, -15.2491, -15.12742, 
    -15.00559, -14.88359, -14.76143, -14.63911, -14.51663, -14.39399, 
    -14.27119, -14.14823, -14.0251, -13.90182, -13.77838, -13.65477, 
    -13.53101, -13.40709, -13.283, -13.15876, -13.03436, -12.9098, -12.78508, 
    -12.6602, -12.53516, -12.40996, -12.28461, -12.15909, -12.03342, 
    -11.90759, -11.7816, -11.65545, -11.52915, -11.40269, -11.27607, 
    -11.1493, -11.02237, -10.89528, -10.76804, -10.64064, -10.51309, 
    -10.38538, -10.25752, -10.1295, -10.00132, -9.872997, -9.744515, 
    -9.615881, -9.487092, -9.35815, -9.229055, -9.099809, -8.970409, 
    -8.840858, -8.711156, -8.581302, -8.451297, -8.321142, -8.190836, 
    -8.060381, -7.929775, -7.799021, -7.668118, -7.537066, -7.405867, 
    -7.274519, -7.143024, -7.011383, -6.879594, -6.74766, -6.615579, 
    -6.483354, -6.350983, -6.218468, -6.085809, -5.953006, -5.82006, 
    -5.686971, -5.55374, -5.420367, -5.286852, -5.153197, -5.019401, 
    -4.885465, -4.75139, -4.617175, -4.482822, -4.348331, -4.213702, 
    -4.078937, -3.944035, -3.808996, -3.673823, -3.538514, -3.403071, 
    -3.267494, -3.131784, -2.995942, -2.859967, -2.72386, -2.587622, 
    -2.451254, -2.314756, -2.178129, -2.041373, -1.904489, -1.767477, 
    -1.630338, -1.493074, -1.355683, -1.218168, -1.080528, -0.9427645, 
    -0.8048778, -0.6668687, -0.5287378, -0.3904858, -0.2521133, -0.113621, 
    0.02499039, 0.1637202, 0.3025678, 0.4415324, 0.5806133, 0.7198099, 
    0.8591214, 0.9985471, 1.138086, 1.277738, 1.417502, 1.557378, 1.697364, 
    1.837459, 1.977664, 2.117977, 2.258398, 2.398925, 2.539558, 2.680297, 
    2.82114, 2.962086, 3.103136, 3.244287, 3.38554, 3.526893, 3.668346, 
    3.809897, 3.951547, 4.093294, 4.235137, 4.377075, 4.519108, 4.661235, 
    4.803455, 4.945767, 5.08817, 5.230663, 5.373246, 5.515918, 5.658677, 
    5.801523, 5.944455, 6.087472, 6.230573, 6.373757, 6.517024, 6.660372, 
    6.803801, 6.947309, 7.090896, 7.23456, 7.378302, 7.522119, 7.666011, 
    7.809978, 7.954017, 8.098128, 8.242311, 8.386563, 8.530885, 8.675275, 
    8.819733, 8.964256, 9.108845, 9.253498, 9.398214, 9.542994, 9.687834, 
    9.832735, 9.977695, 10.12271, 10.26779, 10.41292, 10.55811, 10.70335, 
    10.84865, 10.99399, 11.13939, 11.28484, 11.43034, 11.57588, 11.72148, 
    11.86712, 12.0128, 12.15853, 12.3043, 12.45012, 12.59597, 12.74187, 
    12.8878, 13.03377, 13.17978, 13.32582, 13.4719, 13.61801, 13.76415, 
    13.91033, 14.05654, 14.20277, 14.34903, 14.49532, 14.64164, 14.78798, 
    14.93435, 15.08073, 15.22714, 15.37357, 15.52002, 15.66649, 15.81297, 
    15.95948, 16.10599, 16.25252, 16.39907, 16.54562, 16.69219, 16.83877, 
    16.98535, 17.13194, 17.27854, 17.42515, 17.57175, 17.71837, 17.86498, 
    18.0116, 18.15821, 18.30482, 18.45144, 18.59804, 18.74465, 18.89125, 
    19.03784, 19.18442, 19.331, 19.47756, 19.62411, 19.77066, 19.91718, 
    20.0637, 20.2102, 20.35668, 20.50315, 20.64959, 20.79602, 20.94242, 
    21.08881, 21.23517, 21.38151, 21.52782, 21.6741, 21.82036, 21.96659, 
    22.11279, 22.25896, 22.4051, 22.55121, 22.69728, 22.84332, 22.98932, 
    23.13529, 23.28121, 23.4271, 23.57295, 23.71876, 23.86452, 24.01024, 
    24.15592, 24.30156, 24.44714, 24.59268, 24.73817, 24.88361, 25.029, 
    25.17434, 25.31963, 25.46486, 25.61004, 25.75516, 25.90023, 26.04524, 
    26.19019, 26.33508, 26.47991, 26.62468, 26.76939, 26.91403, 27.05861, 
    27.20312, 27.34757, 27.49195, 27.63626, 27.7805, 27.92467, 28.06877, 
    28.2128, 28.35675, 28.50064, 28.64444, 28.78817, 28.93182, 29.0754, 
    29.21889, 29.36231, 29.50564, 29.6489, 29.79207, 29.93516, 30.07816, 
    30.22108, 30.36391, 30.50666, 30.64931, 30.79188, 30.93436, 31.07675, 
    31.21905, 31.36125, 31.50336, 31.64538, 31.78731, 31.92913, 32.07087, 
    32.2125, 32.35403, 32.49547, 32.63681, 32.77805, 32.91918, 33.06021, 
    33.20115, 33.34197, 33.4827, 33.62331, 33.76382, 33.90422, 34.04452, 
    34.18471, 34.32479, 34.46476, 34.60461, 34.74436, 34.884, 35.02351, 
    35.16292, 35.30222, 35.44139, 35.58046, 35.7194, 35.85823, 35.99694, 
    36.13554, 36.27401, 36.41236, 36.55059, 36.68871, 36.8267, 36.96457, 
    37.10231, 37.23993, 37.37743, 37.51479, 37.65204, 37.78916, 37.92615, 
    38.06301, 38.19975, 38.33636, 38.47284, 38.60918, 38.7454, 38.88148, 
    39.01744, 39.15326, 39.28895, 39.4245, 39.55993, 39.69521, 39.83037, 
    39.96538, 40.10027, 40.23501, 40.36961, 40.50409, 40.63842, 40.77261, 
    40.90666, 41.04057, 41.17435, 41.30798, 41.44147, 41.57483, 41.70803, 
    41.8411, 41.97402, 42.1068, 42.23944,
  -17.9468, -17.82854, -17.71013, -17.59155, -17.47281, -17.3539, -17.23484, 
    -17.11561, -16.99622, -16.87666, -16.75694, -16.63706, -16.51702, 
    -16.39682, -16.27645, -16.15592, -16.03522, -15.91437, -15.79335, 
    -15.67217, -15.55083, -15.42932, -15.30765, -15.18582, -15.06383, 
    -14.94168, -14.81936, -14.69689, -14.57425, -14.45145, -14.32849, 
    -14.20536, -14.08208, -13.95863, -13.83503, -13.71126, -13.58733, 
    -13.46324, -13.33899, -13.21458, -13.09001, -12.96528, -12.84039, 
    -12.71534, -12.59013, -12.46476, -12.33923, -12.21354, -12.08769, 
    -11.96169, -11.83552, -11.7092, -11.58272, -11.45608, -11.32928, 
    -11.20233, -11.07522, -10.94795, -10.82052, -10.69294, -10.5652, 
    -10.43731, -10.30926, -10.18105, -10.05269, -9.924177, -9.795506, 
    -9.666681, -9.537702, -9.408568, -9.279281, -9.14984, -9.020247, 
    -8.890501, -8.760602, -8.630552, -8.500349, -8.369996, -8.239491, 
    -8.108835, -7.978029, -7.847074, -7.715968, -7.584713, -7.453309, 
    -7.321757, -7.190056, -7.058208, -6.926212, -6.79407, -6.66178, 
    -6.529345, -6.396764, -6.264038, -6.131166, -5.99815, -5.86499, 
    -5.731687, -5.59824, -5.464651, -5.33092, -5.197046, -5.063032, 
    -4.928876, -4.794581, -4.660145, -4.52557, -4.390857, -4.256005, 
    -4.121015, -3.985888, -3.850624, -3.715224, -3.579688, -3.444017, 
    -3.308211, -3.172271, -3.036198, -2.899992, -2.763653, -2.627183, 
    -2.490581, -2.353849, -2.216986, -2.079994, -1.942874, -1.805625, 
    -1.668248, -1.530745, -1.393115, -1.255359, -1.117478, -0.9794725, 
    -0.8413433, -0.7030909, -0.564716, -0.4262192, -0.2876012, -0.1488627, 
    -0.01000442, 0.128973, 0.268069, 0.4072827, 0.5466134, 0.6860604, 
    0.8256232, 0.9653008, 1.105093, 1.244998, 1.385016, 1.525146, 1.665387, 
    1.805739, 1.9462, 2.086771, 2.227449, 2.368235, 2.509128, 2.650126, 
    2.79123, 2.932438, 3.073749, 3.215163, 3.356679, 3.498296, 3.640013, 
    3.78183, 3.923745, 4.065758, 4.207868, 4.350074, 4.492375, 4.63477, 
    4.77726, 4.919841, 5.062515, 5.205279, 5.348134, 5.491077, 5.634109, 
    5.777228, 5.920434, 6.063725, 6.207101, 6.350561, 6.494104, 6.637728, 
    6.781434, 6.92522, 7.069085, 7.213027, 7.357048, 7.501145, 7.645317, 
    7.789564, 7.933884, 8.078277, 8.22274, 8.367275, 8.51188, 8.656553, 
    8.801294, 8.946101, 9.090975, 9.235913, 9.380915, 9.525979, 9.671105, 
    9.816293, 9.96154, 10.10685, 10.25221, 10.39763, 10.54311, 10.68864, 
    10.83422, 10.97986, 11.12554, 11.27128, 11.41707, 11.56291, 11.70879, 
    11.85472, 12.0007, 12.14672, 12.29279, 12.43889, 12.58504, 12.73123, 
    12.87745, 13.02372, 13.17002, 13.31636, 13.46273, 13.60913, 13.75557, 
    13.90204, 14.04854, 14.19507, 14.34163, 14.48822, 14.63483, 14.78147, 
    14.92813, 15.07481, 15.22152, 15.36824, 15.51499, 15.66175, 15.80854, 
    15.95533, 16.10215, 16.24898, 16.39582, 16.54267, 16.68953, 16.83641, 
    16.98329, 17.13018, 17.27708, 17.42398, 17.57088, 17.71779, 17.86471, 
    18.01162, 18.15853, 18.30544, 18.45235, 18.59926, 18.74616, 18.89305, 
    19.03995, 19.18683, 19.3337, 19.48056, 19.62741, 19.77425, 19.92108, 
    20.06789, 20.21468, 20.36146, 20.50823, 20.65497, 20.80169, 20.94839, 
    21.09507, 21.24173, 21.38836, 21.53497, 21.68155, 21.82811, 21.97463, 
    22.12113, 22.26759, 22.41403, 22.56043, 22.70679, 22.85313, 22.99942, 
    23.14568, 23.2919, 23.43808, 23.58422, 23.73032, 23.87638, 24.02239, 
    24.16836, 24.31429, 24.46016, 24.60599, 24.75177, 24.8975, 25.04318, 
    25.18881, 25.33439, 25.47991, 25.62538, 25.77079, 25.91614, 26.06144, 
    26.20668, 26.35185, 26.49697, 26.64203, 26.78702, 26.93195, 27.07681, 
    27.22161, 27.36634, 27.511, 27.65559, 27.80012, 27.94457, 28.08895, 
    28.23326, 28.37749, 28.52165, 28.66574, 28.80975, 28.95368, 29.09753, 
    29.2413, 29.385, 29.52861, 29.67214, 29.81558, 29.95895, 30.10222, 
    30.24542, 30.38852, 30.53154, 30.67447, 30.81731, 30.96006, 31.10272, 
    31.24529, 31.38776, 31.53014, 31.67243, 31.81462, 31.95671, 32.09871, 
    32.24061, 32.38241, 32.52411, 32.66571, 32.80721, 32.94861, 33.0899, 
    33.2311, 33.37218, 33.51316, 33.65404, 33.79481, 33.93547, 34.07603, 
    34.21647, 34.3568, 34.49703, 34.63714, 34.77714, 34.91703, 35.0568, 
    35.19646, 35.33601, 35.47543, 35.61475, 35.75394, 35.89302, 36.03198, 
    36.17082, 36.30954, 36.44814, 36.58661, 36.72497, 36.8632, 37.00131, 
    37.1393, 37.27716, 37.41489, 37.55251, 37.68999, 37.82734, 37.96457, 
    38.10167, 38.23864, 38.37548, 38.5122, 38.64878, 38.78523, 38.92155, 
    39.05773, 39.19378, 39.3297, 39.46549, 39.60114, 39.73665, 39.87203, 
    40.00727, 40.14238, 40.27734, 40.41217, 40.54687, 40.68142, 40.81583, 
    40.95011, 41.08424, 41.21823, 41.35209, 41.48579, 41.61936, 41.75278, 
    41.88606, 42.0192, 42.15219, 42.28504,
  -18.00872, -17.89033, -17.77177, -17.65306, -17.53417, -17.41513, 
    -17.29592, -17.17655, -17.05701, -16.93731, -16.81745, -16.69742, 
    -16.57724, -16.45688, -16.33637, -16.21569, -16.09484, -15.97384, 
    -15.85267, -15.73134, -15.60984, -15.48818, -15.36636, -15.24438, 
    -15.12223, -14.99992, -14.87745, -14.75481, -14.63201, -14.50905, 
    -14.38593, -14.26265, -14.1392, -14.01559, -13.89182, -13.76789, 
    -13.6438, -13.51954, -13.39512, -13.27055, -13.14581, -13.02091, 
    -12.89585, -12.77062, -12.64524, -12.5197, -12.394, -12.26814, -12.14211, 
    -12.01593, -11.88959, -11.76309, -11.63643, -11.50961, -11.38264, 
    -11.2555, -11.12821, -11.00076, -10.87315, -10.74539, -10.61746, 
    -10.48938, -10.36115, -10.23275, -10.10421, -9.975501, -9.846641, 
    -9.717625, -9.588454, -9.459128, -9.329649, -9.200014, -9.070227, 
    -8.940285, -8.81019, -8.679943, -8.549542, -8.41899, -8.288286, -8.15743, 
    -8.026423, -7.895265, -7.763957, -7.632498, -7.50089, -7.369133, 
    -7.237226, -7.105171, -6.972968, -6.840616, -6.708118, -6.575472, 
    -6.44268, -6.309742, -6.176658, -6.043429, -5.910055, -5.776536, 
    -5.642874, -5.509068, -5.375119, -5.241027, -5.106794, -4.972419, 
    -4.837903, -4.703246, -4.568449, -4.433512, -4.298436, -4.163221, 
    -4.027869, -3.892379, -3.756752, -3.620988, -3.485088, -3.349053, 
    -3.212883, -3.076579, -2.940141, -2.80357, -2.666866, -2.53003, 
    -2.393063, -2.255965, -2.118737, -1.981379, -1.843892, -1.706277, 
    -1.568534, -1.430664, -1.292667, -1.154544, -1.016297, -0.8779243, 
    -0.739428, -0.6008084, -0.4620663, -0.3232022, -0.1842169, -0.04511097, 
    0.09411478, 0.2334597, 0.3729231, 0.5125043, 0.6522025, 0.792017, 
    0.9319472, 1.071992, 1.212152, 1.352424, 1.492809, 1.633307, 1.773915, 
    1.914634, 2.055462, 2.1964, 2.337445, 2.478598, 2.619857, 2.761222, 
    2.902692, 3.044266, 3.185943, 3.327723, 3.469604, 3.611587, 3.75367, 
    3.895851, 4.038131, 4.180509, 4.322983, 4.465553, 4.608218, 4.750977, 
    4.893829, 5.036774, 5.179811, 5.322937, 5.466154, 5.609459, 5.752852, 
    5.896333, 6.039899, 6.183551, 6.327287, 6.471107, 6.615008, 6.758992, 
    6.903056, 7.047199, 7.191422, 7.335722, 7.480099, 7.624552, 7.76908, 
    7.913682, 8.058357, 8.203104, 8.347921, 8.49281, 8.637767, 8.782793, 
    8.927885, 9.073044, 9.218267, 9.363556, 9.508907, 9.654321, 9.799795, 
    9.94533, 10.09092, 10.23658, 10.38228, 10.52805, 10.67387, 10.81974, 
    10.96567, 11.11165, 11.25768, 11.40376, 11.54989, 11.69607, 11.84229, 
    11.98856, 12.13487, 12.28123, 12.42763, 12.57407, 12.72055, 12.86707, 
    13.01363, 13.16023, 13.30686, 13.45353, 13.60023, 13.74696, 13.89373, 
    14.04052, 14.18735, 14.3342, 14.48109, 14.628, 14.77493, 14.92189, 
    15.06887, 15.21587, 15.3629, 15.50994, 15.657, 15.80408, 15.95118, 
    16.09829, 16.24542, 16.39256, 16.53971, 16.68687, 16.83404, 16.98122, 
    17.12841, 17.27561, 17.42281, 17.57001, 17.71722, 17.86443, 18.01164, 
    18.15886, 18.30606, 18.45327, 18.60048, 18.74768, 18.89487, 19.04206, 
    19.18924, 19.33641, 19.48357, 19.63072, 19.77786, 19.92498, 20.07209, 
    20.21918, 20.36626, 20.51332, 20.66036, 20.80738, 20.95438, 21.10136, 
    21.24832, 21.39524, 21.54215, 21.68903, 21.83588, 21.9827, 22.12949, 
    22.27625, 22.42298, 22.56968, 22.71634, 22.86296, 23.00956, 23.15611, 
    23.30262, 23.4491, 23.59553, 23.74193, 23.88828, 24.03458, 24.18085, 
    24.32706, 24.47323, 24.61935, 24.76542, 24.91145, 25.05742, 25.20333, 
    25.3492, 25.49501, 25.64077, 25.78647, 25.93211, 26.0777, 26.22322, 
    26.36869, 26.51409, 26.65943, 26.80471, 26.94992, 27.09507, 27.24015, 
    27.38517, 27.53011, 27.67499, 27.8198, 27.96453, 28.1092, 28.25379, 
    28.3983, 28.54274, 28.68711, 28.8314, 28.97561, 29.11974, 29.26379, 
    29.40776, 29.55165, 29.69546, 29.83918, 29.98282, 30.12637, 30.26984, 
    30.41322, 30.55651, 30.69971, 30.84282, 30.98584, 31.12877, 31.27161, 
    31.41436, 31.557, 31.69956, 31.84202, 31.98438, 32.12665, 32.26881, 
    32.41088, 32.55285, 32.69471, 32.83648, 32.97813, 33.11969, 33.26115, 
    33.4025, 33.54374, 33.68487, 33.8259, 33.96682, 34.10763, 34.24833, 
    34.38892, 34.5294, 34.66977, 34.81003, 34.95017, 35.09019, 35.23011, 
    35.3699, 35.50958, 35.64915, 35.78859, 35.92792, 36.06712, 36.20621, 
    36.34518, 36.48402, 36.62275, 36.76134, 36.89982, 37.03817, 37.1764, 
    37.3145, 37.45248, 37.59033, 37.72805, 37.86565, 38.00312, 38.14045, 
    38.27766, 38.41474, 38.55169, 38.6885, 38.82518, 38.96173, 39.09815, 
    39.23443, 39.37058, 39.5066, 39.64247, 39.77821, 39.91382, 40.04929, 
    40.18462, 40.31981, 40.45486, 40.58978, 40.72456, 40.85919, 40.99368, 
    41.12804, 41.26225, 41.39632, 41.53024, 41.66403, 41.79766, 41.93116, 
    42.06451, 42.19772, 42.33078,
  -18.07079, -17.95226, -17.83357, -17.71471, -17.59569, -17.4765, -17.35715, 
    -17.23764, -17.11796, -16.99811, -16.87811, -16.75793, -16.6376, 
    -16.5171, -16.39643, -16.27561, -16.15462, -16.03346, -15.91214, 
    -15.79065, -15.66901, -15.54719, -15.42522, -15.30308, -15.18078, 
    -15.05831, -14.93568, -14.81289, -14.68993, -14.56681, -14.44353, 
    -14.32008, -14.19647, -14.0727, -13.94877, -13.82467, -13.70041, 
    -13.57599, -13.45141, -13.32666, -13.20175, -13.07668, -12.95145, 
    -12.82606, -12.70051, -12.57479, -12.44892, -12.32288, -12.19668, 
    -12.07033, -11.94381, -11.81713, -11.69029, -11.5633, -11.43614, 
    -11.30882, -11.18135, -11.05372, -10.92593, -10.79798, -10.66987, 
    -10.5416, -10.41318, -10.2846, -10.15586, -10.02697, -9.897919, 
    -9.768712, -9.63935, -9.509832, -9.380159, -9.250331, -9.120348, 
    -8.990211, -8.859921, -8.729475, -8.598877, -8.468125, -8.337222, 
    -8.206165, -8.074957, -7.943597, -7.812085, -7.680423, -7.54861, 
    -7.416647, -7.284534, -7.152272, -7.01986, -6.8873, -6.754592, -6.621736, 
    -6.488733, -6.355582, -6.222286, -6.088842, -5.955254, -5.82152, 
    -5.687642, -5.553618, -5.419452, -5.285141, -5.150689, -5.016093, 
    -4.881356, -4.746477, -4.611457, -4.476297, -4.340997, -4.205557, 
    -4.069978, -3.934262, -3.798407, -3.662415, -3.526286, -3.390021, 
    -3.253621, -3.117085, -2.980415, -2.843611, -2.706673, -2.569602, 
    -2.4324, -2.295066, -2.157601, -2.020005, -1.88228, -1.744425, -1.606442, 
    -1.468331, -1.330093, -1.191728, -1.053238, -0.9146215, -0.7758807, 
    -0.6370159, -0.4980277, -0.3589169, -0.2196841, -0.08033003, 0.05914465, 
    0.1987392, 0.338453, 0.4782853, 0.6182353, 0.7583024, 0.8984858, 
    1.038785, 1.179199, 1.319727, 1.460368, 1.601122, 1.741988, 1.882965, 
    2.024052, 2.165249, 2.306554, 2.447968, 2.589488, 2.731115, 2.872848, 
    3.014685, 3.156627, 3.298671, 3.440818, 3.583066, 3.725416, 3.867864, 
    4.010412, 4.153059, 4.295802, 4.438642, 4.581577, 4.724607, 4.867731, 
    5.010947, 5.154256, 5.297656, 5.441146, 5.584726, 5.728395, 5.87215, 
    6.015993, 6.159921, 6.303934, 6.448031, 6.592211, 6.736474, 6.880816, 
    7.02524, 7.169743, 7.314324, 7.458982, 7.603717, 7.748527, 7.893411, 
    8.038369, 8.1834, 8.328502, 8.473675, 8.618917, 8.764228, 8.909606, 
    9.055052, 9.200562, 9.346137, 9.491776, 9.637477, 9.78324, 9.929064, 
    10.07495, 10.22089, 10.36689, 10.51294, 10.65905, 10.80522, 10.95144, 
    11.09771, 11.24403, 11.3904, 11.53682, 11.68329, 11.82981, 11.97637, 
    12.12298, 12.26963, 12.41632, 12.56306, 12.70984, 12.85665, 13.00351, 
    13.1504, 13.29733, 13.44429, 13.59129, 13.73832, 13.88538, 14.03248, 
    14.1796, 14.32675, 14.47393, 14.62114, 14.76837, 14.91563, 15.06291, 
    15.21021, 15.35753, 15.50487, 15.65223, 15.79961, 15.94701, 16.09442, 
    16.24184, 16.38928, 16.53673, 16.68419, 16.83167, 16.97915, 17.12664, 
    17.27413, 17.42163, 17.56914, 17.71665, 17.86415, 18.01167, 18.15918, 
    18.30669, 18.4542, 18.6017, 18.7492, 18.89669, 19.04418, 19.19166, 
    19.33913, 19.48659, 19.63404, 19.78148, 19.9289, 20.07631, 20.2237, 
    20.37108, 20.51844, 20.66578, 20.8131, 20.96039, 21.10767, 21.25492, 
    21.40215, 21.54935, 21.69653, 21.84368, 21.99079, 22.13788, 22.28494, 
    22.43197, 22.57896, 22.72592, 22.87284, 23.01973, 23.16657, 23.31338, 
    23.46015, 23.60688, 23.75357, 23.90022, 24.04682, 24.19337, 24.33988, 
    24.48634, 24.63276, 24.77912, 24.92543, 25.0717, 25.21791, 25.36406, 
    25.51016, 25.65621, 25.8022, 25.94813, 26.09401, 26.23982, 26.38557, 
    26.53127, 26.6769, 26.82246, 26.96796, 27.11339, 27.25876, 27.40406, 
    27.54929, 27.69446, 27.83955, 27.98457, 28.12951, 28.27439, 28.41918, 
    28.56391, 28.70855, 28.85312, 28.99761, 29.14202, 29.28635, 29.4306, 
    29.57477, 29.71885, 29.86285, 30.00677, 30.15059, 30.29434, 30.43799, 
    30.58156, 30.72503, 30.86842, 31.01171, 31.15491, 31.29803, 31.44104, 
    31.58396, 31.72678, 31.86951, 32.01214, 32.15467, 32.29711, 32.43944, 
    32.58167, 32.7238, 32.86583, 33.00776, 33.14958, 33.29129, 33.43291, 
    33.57441, 33.71581, 33.85709, 33.99827, 34.13934, 34.2803, 34.42115, 
    34.56189, 34.70251, 34.84302, 34.98342, 35.1237, 35.26386, 35.40391, 
    35.54384, 35.68365, 35.82335, 35.96292, 36.10238, 36.24172, 36.38093, 
    36.52002, 36.65899, 36.79784, 36.93656, 37.07515, 37.21362, 37.35197, 
    37.49019, 37.62828, 37.76624, 37.90408, 38.04178, 38.17936, 38.3168, 
    38.45411, 38.59129, 38.72834, 38.86526, 39.00204, 39.13869, 39.27521, 
    39.41159, 39.54783, 39.68394, 39.8199, 39.95574, 40.09143, 40.22699, 
    40.36241, 40.49768, 40.63282, 40.76782, 40.90268, 41.03739, 41.17197, 
    41.3064, 41.44069, 41.57483, 41.70883, 41.84269, 41.97639, 42.10996, 
    42.24338, 42.37666,
  -18.13301, -18.01435, -17.89551, -17.77652, -17.65735, -17.53803, 
    -17.41853, -17.29888, -17.17905, -17.05907, -16.93891, -16.8186, 
    -16.69811, -16.57747, -16.45666, -16.33568, -16.21454, -16.09323, 
    -15.97176, -15.85012, -15.72832, -15.60636, -15.48423, -15.36193, 
    -15.23947, -15.11685, -14.99406, -14.87111, -14.748, -14.62472, 
    -14.50127, -14.37767, -14.25389, -14.12996, -14.00586, -13.8816, 
    -13.75718, -13.63259, -13.50784, -13.38292, -13.25785, -13.13261, 
    -13.00721, -12.88164, -12.75592, -12.63003, -12.50398, -12.37777, 
    -12.2514, -12.12487, -11.99817, -11.87132, -11.7443, -11.61713, 
    -11.48979, -11.36229, -11.23464, -11.10682, -10.97885, -10.85071, 
    -10.72242, -10.59397, -10.46536, -10.33659, -10.20767, -10.07858, 
    -9.949342, -9.819945, -9.690391, -9.56068, -9.430814, -9.300792, 
    -9.170614, -9.040281, -8.909793, -8.779151, -8.648354, -8.517404, 
    -8.386299, -8.255042, -8.123632, -7.992069, -7.860354, -7.728488, 
    -7.59647, -7.464301, -7.331981, -7.199512, -7.066892, -6.934123, 
    -6.801204, -6.668138, -6.534923, -6.40156, -6.268049, -6.134392, 
    -6.000588, -5.866639, -5.732544, -5.598303, -5.463918, -5.329389, 
    -5.194716, -5.0599, -4.924941, -4.78984, -4.654597, -4.519213, -4.383687, 
    -4.248023, -4.112217, -3.976274, -3.840191, -3.70397, -3.567612, 
    -3.431116, -3.294485, -3.157717, -3.020814, -2.883776, -2.746604, 
    -2.609299, -2.47186, -2.33429, -2.196587, -2.058753, -1.920789, 
    -1.782694, -1.644471, -1.506119, -1.367638, -1.229031, -1.090296, 
    -0.9514357, -0.8124498, -0.6733391, -0.5341043, -0.3947462, -0.2552653, 
    -0.1156624, 0.02406188, 0.1639068, 0.3038716, 0.4439556, 0.5841581, 
    0.7244784, 0.8649157, 1.005469, 1.146138, 1.286922, 1.427821, 1.568832, 
    1.709956, 1.851192, 1.992538, 2.133995, 2.275561, 2.417237, 2.559019, 
    2.700909, 2.842905, 2.985007, 3.127213, 3.269523, 3.411936, 3.554451, 
    3.697068, 3.839785, 3.982601, 4.125516, 4.268529, 4.41164, 4.554846, 
    4.698148, 4.841544, 4.985034, 5.128616, 5.27229, 5.416055, 5.55991, 
    5.703854, 5.847886, 5.992005, 6.136211, 6.280502, 6.424878, 6.569337, 
    6.713879, 6.858502, 7.003206, 7.14799, 7.292852, 7.437793, 7.58281, 
    7.727903, 7.873072, 8.018313, 8.163629, 8.309016, 8.454474, 8.600002, 
    8.7456, 8.891265, 9.036997, 9.182796, 9.328658, 9.474586, 9.620576, 
    9.766628, 9.912742, 10.05891, 10.20515, 10.35144, 10.49778, 10.64419, 
    10.79064, 10.93715, 11.08372, 11.23033, 11.377, 11.52371, 11.67048, 
    11.81729, 11.96414, 12.11105, 12.25799, 12.40498, 12.55201, 12.69909, 
    12.8462, 12.99335, 13.14054, 13.28776, 13.43502, 13.58232, 13.72965, 
    13.87701, 14.0244, 14.17182, 14.31927, 14.46675, 14.61426, 14.76179, 
    14.90934, 15.05692, 15.20452, 15.35214, 15.49979, 15.64745, 15.79513, 
    15.94282, 16.09053, 16.23826, 16.386, 16.53375, 16.68151, 16.82928, 
    16.97707, 17.12486, 17.27265, 17.42045, 17.56826, 17.71607, 17.86388, 
    18.01169, 18.1595, 18.30731, 18.45512, 18.60293, 18.75073, 18.89852, 
    19.04631, 19.19409, 19.34186, 19.48962, 19.63737, 19.78511, 19.93283, 
    20.08054, 20.22824, 20.37591, 20.52357, 20.67121, 20.81883, 20.96642, 
    21.114, 21.26155, 21.40908, 21.55658, 21.70405, 21.8515, 21.99892, 
    22.14631, 22.29366, 22.44098, 22.58827, 22.73553, 22.88275, 23.02993, 
    23.17707, 23.32418, 23.47125, 23.61827, 23.76525, 23.9122, 24.05909, 
    24.20594, 24.35274, 24.4995, 24.64621, 24.79286, 24.93947, 25.08603, 
    25.23253, 25.37898, 25.52537, 25.67171, 25.81799, 25.96421, 26.11038, 
    26.25648, 26.40252, 26.5485, 26.69442, 26.84027, 26.98606, 27.13178, 
    27.27744, 27.42302, 27.56854, 27.71399, 27.85936, 28.00467, 28.1499, 
    28.29505, 28.44013, 28.58514, 28.73007, 28.87492, 29.01969, 29.16438, 
    29.30899, 29.45352, 29.59797, 29.74233, 29.88661, 30.0308, 30.1749, 
    30.31892, 30.46285, 30.60669, 30.75044, 30.8941, 31.03767, 31.18114, 
    31.32453, 31.46781, 31.611, 31.7541, 31.8971, 32.04, 32.1828, 32.3255, 
    32.4681, 32.6106, 32.75299, 32.89529, 33.03748, 33.17956, 33.32154, 
    33.46342, 33.60518, 33.74684, 33.88839, 34.02983, 34.17116, 34.31237, 
    34.45348, 34.59447, 34.73536, 34.87612, 35.01677, 35.15731, 35.29773, 
    35.43803, 35.57821, 35.71828, 35.85822, 35.99805, 36.13775, 36.27734, 
    36.4168, 36.55614, 36.69535, 36.83444, 36.97341, 37.11225, 37.25097, 
    37.38955, 37.52801, 37.66634, 37.80455, 37.94262, 38.08057, 38.21838, 
    38.35606, 38.49361, 38.63103, 38.76831, 38.90546, 39.04248, 39.17936, 
    39.3161, 39.45272, 39.58919, 39.72553, 39.86172, 39.99779, 40.13371, 
    40.26949, 40.40514, 40.54064, 40.676, 40.81122, 40.9463, 41.08123, 
    41.21603, 41.35068, 41.48518, 41.61955, 41.75377, 41.88784, 42.02176, 
    42.15554, 42.28918, 42.42266,
  -18.19539, -18.07658, -17.95761, -17.83847, -17.71917, -17.5997, -17.48007, 
    -17.36027, -17.2403, -17.12017, -16.99987, -16.87941, -16.75878, 
    -16.63799, -16.51702, -16.3959, -16.27461, -16.15315, -16.03153, 
    -15.90974, -15.78779, -15.66567, -15.54339, -15.42094, -15.29832, 
    -15.17554, -15.0526, -14.92949, -14.80621, -14.68277, -14.55917, 
    -14.4354, -14.31147, -14.18737, -14.06311, -13.93868, -13.81409, 
    -13.68934, -13.56442, -13.43934, -13.31409, -13.18869, -13.06311, 
    -12.93738, -12.81148, -12.68542, -12.5592, -12.43281, -12.30627, 
    -12.17956, -12.05269, -11.92565, -11.79846, -11.6711, -11.54359, 
    -11.41591, -11.28807, -11.16007, -11.03191, -10.9036, -10.77512, 
    -10.64648, -10.51768, -10.38873, -10.25961, -10.13034, -10.00091, 
    -9.871324, -9.741577, -9.611674, -9.481614, -9.351398, -9.221025, 
    -9.090495, -8.95981, -8.82897, -8.697974, -8.566824, -8.43552, -8.304062, 
    -8.172449, -8.040684, -7.908765, -7.776694, -7.644471, -7.512096, 
    -7.379569, -7.246891, -7.114063, -6.981084, -6.847956, -6.714677, 
    -6.58125, -6.447675, -6.313951, -6.180079, -6.04606, -5.911894, 
    -5.777582, -5.643124, -5.50852, -5.373771, -5.238878, -5.10384, 
    -4.968659, -4.833335, -4.697869, -4.56226, -4.42651, -4.290619, 
    -4.154587, -4.018415, -3.882104, -3.745654, -3.609066, -3.472339, 
    -3.335476, -3.198476, -3.06134, -2.924068, -2.786661, -2.64912, 
    -2.511445, -2.373637, -2.235696, -2.097624, -1.959419, -1.821085, 
    -1.68262, -1.544026, -1.405303, -1.266452, -1.127473, -0.9883678, 
    -0.8491361, -0.709779, -0.5702969, -0.4306908, -0.2909612, -0.1511088, 
    -0.01113432, 0.1289615, 0.269178, 0.4095144, 0.5499701, 0.6905442, 
    0.8312361, 0.9720451, 1.11297, 1.254011, 1.395166, 1.536436, 1.677819, 
    1.819314, 1.960921, 2.102639, 2.244467, 2.386404, 2.52845, 2.670603, 
    2.812864, 2.95523, 3.097702, 3.240278, 3.382958, 3.525741, 3.668625, 
    3.811611, 3.954697, 4.097882, 4.241166, 4.384548, 4.528026, 4.6716, 
    4.815269, 4.959033, 5.102889, 5.246838, 5.390879, 5.53501, 5.67923, 
    5.82354, 5.967937, 6.112421, 6.25699, 6.401646, 6.546384, 6.691206, 
    6.836111, 6.981096, 7.126163, 7.271307, 7.416531, 7.561832, 7.707209, 
    7.852662, 7.998189, 8.143789, 8.289462, 8.435207, 8.581022, 8.726907, 
    8.87286, 9.01888, 9.164967, 9.311119, 9.457336, 9.603616, 9.749959, 
    9.896362, 10.04283, 10.18935, 10.33593, 10.48257, 10.62927, 10.77602, 
    10.92282, 11.06968, 11.21659, 11.36355, 11.51056, 11.65761, 11.80472, 
    11.95187, 12.09907, 12.24631, 12.3936, 12.54093, 12.6883, 12.83571, 
    12.98316, 13.13064, 13.27816, 13.42572, 13.57332, 13.72094, 13.8686, 
    14.0163, 14.16402, 14.31177, 14.45955, 14.60735, 14.75518, 14.90304, 
    15.05092, 15.19882, 15.34674, 15.49468, 15.64264, 15.79062, 15.93862, 
    16.08663, 16.23466, 16.3827, 16.53076, 16.67882, 16.82689, 16.97498, 
    17.12307, 17.27117, 17.41927, 17.56738, 17.71549, 17.8636, 18.01171, 
    18.15983, 18.30794, 18.45605, 18.60416, 18.75226, 18.90036, 19.04845, 
    19.19653, 19.3446, 19.49266, 19.64072, 19.78876, 19.93678, 20.08479, 
    20.23278, 20.38076, 20.52872, 20.67666, 20.82458, 20.97248, 21.12035, 
    21.26821, 21.41603, 21.56383, 21.71161, 21.85935, 22.00707, 22.15475, 
    22.30241, 22.45003, 22.59762, 22.74517, 22.89269, 23.04017, 23.18761, 
    23.33502, 23.48238, 23.6297, 23.77698, 23.92422, 24.07141, 24.21855, 
    24.36565, 24.5127, 24.6597, 24.80666, 24.95356, 25.10041, 25.2472, 
    25.39394, 25.54063, 25.68726, 25.83383, 25.98034, 26.1268, 26.2732, 
    26.41953, 26.5658, 26.712, 26.85815, 27.00422, 27.15023, 27.29618, 
    27.44205, 27.58785, 27.73359, 27.87925, 28.02484, 28.17035, 28.31579, 
    28.46116, 28.60645, 28.75166, 28.89679, 29.04184, 29.18682, 29.33171, 
    29.47652, 29.62124, 29.76588, 29.91044, 30.05491, 30.19929, 30.34359, 
    30.48779, 30.63191, 30.77594, 30.91987, 31.06371, 31.20746, 31.35112, 
    31.49468, 31.63814, 31.78151, 31.92477, 32.06794, 32.21101, 32.35398, 
    32.49685, 32.63962, 32.78228, 32.92484, 33.0673, 33.20965, 33.35189, 
    33.49403, 33.63605, 33.77798, 33.91978, 34.06149, 34.20308, 34.34455, 
    34.48592, 34.62717, 34.76831, 34.90933, 35.05024, 35.19103, 35.3317, 
    35.47226, 35.61269, 35.75301, 35.89321, 36.03328, 36.17324, 36.31307, 
    36.45278, 36.59237, 36.73183, 36.87117, 37.01038, 37.14947, 37.28843, 
    37.42725, 37.56596, 37.70453, 37.84298, 37.98129, 38.11947, 38.25753, 
    38.39544, 38.53323, 38.67089, 38.80841, 38.94579, 39.08304, 39.22016, 
    39.35714, 39.49398, 39.63068, 39.76725, 39.90368, 40.03997, 40.17611, 
    40.31212, 40.44799, 40.58372, 40.71931, 40.85475, 40.99005, 41.12521, 
    41.26023, 41.3951, 41.52982, 41.6644, 41.79884, 41.93313, 42.06727, 
    42.20126, 42.33511, 42.46881,
  -18.25791, -18.13897, -18.01986, -17.90058, -17.78114, -17.66153, 
    -17.54175, -17.42181, -17.3017, -17.18143, -17.06098, -16.94037, 
    -16.8196, -16.69866, -16.57755, -16.45628, -16.33484, -16.21323, 
    -16.09145, -15.96951, -15.84741, -15.72513, -15.6027, -15.48009, 
    -15.35732, -15.23439, -15.11128, -14.98802, -14.86458, -14.74098, 
    -14.61722, -14.49329, -14.36919, -14.24493, -14.12051, -13.99592, 
    -13.87116, -13.74624, -13.62115, -13.4959, -13.37049, -13.24491, 
    -13.11917, -12.99327, -12.8672, -12.74096, -12.61457, -12.48801, 
    -12.36128, -12.2344, -12.10735, -11.98014, -11.85277, -11.72523, 
    -11.59753, -11.46968, -11.34165, -11.21347, -11.08513, -10.95663, 
    -10.82796, -10.69914, -10.57016, -10.44101, -10.31171, -10.18225, 
    -10.05263, -9.922848, -9.79291, -9.662814, -9.532559, -9.402148, 
    -9.27158, -9.140854, -9.009972, -8.878934, -8.747739, -8.616389, 
    -8.484884, -8.353225, -8.22141, -8.089441, -7.957319, -7.825043, 
    -7.692614, -7.560032, -7.427298, -7.294412, -7.161374, -7.028186, 
    -6.894846, -6.761357, -6.627717, -6.493928, -6.35999, -6.225904, 
    -6.091669, -5.957286, -5.822756, -5.68808, -5.553257, -5.418288, 
    -5.283175, -5.147915, -5.012512, -4.876965, -4.741274, -4.605441, 
    -4.469465, -4.333347, -4.197088, -4.060688, -3.924148, -3.787468, 
    -3.650649, -3.513691, -3.376596, -3.239362, -3.101992, -2.964486, 
    -2.826844, -2.689066, -2.551154, -2.413109, -2.274929, -2.136617, 
    -1.998173, -1.859598, -1.720891, -1.582054, -1.443088, -1.303993, 
    -1.16477, -1.025419, -0.8859405, -0.7463362, -0.6066063, -0.4667515, 
    -0.3267726, -0.1866701, -0.04644471, 0.09390273, 0.2343716, 0.3749611, 
    0.5156705, 0.6564992, 0.7974464, 0.9385113, 1.079693, 1.220991, 1.362405, 
    1.503933, 1.645576, 1.787331, 1.929199, 2.071178, 2.213269, 2.355469, 
    2.497778, 2.640196, 2.782722, 2.925354, 3.068092, 3.210935, 3.353883, 
    3.496934, 3.640087, 3.783343, 3.926699, 4.070155, 4.21371, 4.357364, 
    4.501115, 4.644962, 4.788906, 4.932944, 5.077075, 5.2213, 5.365617, 
    5.510025, 5.654523, 5.79911, 5.943786, 6.088549, 6.233398, 6.378334, 
    6.523354, 6.668457, 6.813643, 6.958911, 7.10426, 7.249689, 7.395196, 
    7.540781, 7.686443, 7.832181, 7.977994, 8.123881, 8.269841, 8.415874, 
    8.561976, 8.708149, 8.854391, 9.0007, 9.147077, 9.293519, 9.440026, 
    9.586597, 9.733231, 9.879927, 10.02668, 10.1735, 10.32037, 10.46731, 
    10.61429, 10.76134, 10.90844, 11.05559, 11.20279, 11.35005, 11.49735, 
    11.64471, 11.79211, 11.93956, 12.08705, 12.23459, 12.38218, 12.5298, 
    12.67747, 12.82518, 12.97293, 13.12071, 13.26853, 13.41639, 13.56428, 
    13.71221, 13.86017, 14.00816, 14.15618, 14.30423, 14.45231, 14.60042, 
    14.74855, 14.89671, 15.04489, 15.19309, 15.34132, 15.48956, 15.63783, 
    15.78611, 15.93441, 16.08272, 16.23105, 16.37939, 16.52775, 16.67612, 
    16.82449, 16.97288, 17.12127, 17.26967, 17.41808, 17.56649, 17.7149, 
    17.86332, 18.01174, 18.16016, 18.30857, 18.45699, 18.60539, 18.7538, 
    18.9022, 19.05059, 19.19898, 19.34735, 19.49572, 19.64407, 19.79241, 
    19.94074, 20.08905, 20.23735, 20.38563, 20.53389, 20.68213, 20.83035, 
    20.97855, 21.12673, 21.27488, 21.42301, 21.57111, 21.71919, 21.86723, 
    22.01525, 22.16324, 22.31119, 22.45911, 22.607, 22.75485, 22.90267, 
    23.05045, 23.19819, 23.34589, 23.49355, 23.64117, 23.78875, 23.93628, 
    24.08377, 24.23121, 24.3786, 24.52595, 24.67325, 24.8205, 24.96769, 
    25.11484, 25.26193, 25.40896, 25.55594, 25.70286, 25.84973, 25.99654, 
    26.14328, 26.28997, 26.43659, 26.58315, 26.72965, 26.87608, 27.02245, 
    27.16875, 27.31498, 27.46114, 27.60723, 27.75325, 27.8992, 28.04508, 
    28.19088, 28.3366, 28.48225, 28.62783, 28.77332, 28.91874, 29.06407, 
    29.20933, 29.3545, 29.49959, 29.6446, 29.78952, 29.93436, 30.07911, 
    30.22377, 30.36834, 30.51283, 30.65722, 30.80152, 30.94573, 31.08985, 
    31.23387, 31.3778, 31.52163, 31.66537, 31.809, 31.95254, 32.09599, 
    32.23933, 32.38256, 32.5257, 32.66874, 32.81167, 32.95449, 33.09721, 
    33.23983, 33.38234, 33.52474, 33.66703, 33.80922, 33.95129, 34.09325, 
    34.2351, 34.37684, 34.51846, 34.65997, 34.80137, 34.94265, 35.08381, 
    35.22486, 35.36578, 35.5066, 35.64729, 35.78786, 35.92831, 36.06863, 
    36.20884, 36.34892, 36.48888, 36.62872, 36.76843, 36.90801, 37.04747, 
    37.1868, 37.326, 37.46508, 37.60402, 37.74284, 37.88153, 38.02008, 
    38.1585, 38.29679, 38.43496, 38.57298, 38.71087, 38.84863, 38.98625, 
    39.12373, 39.26108, 39.39829, 39.53537, 39.6723, 39.8091, 39.94576, 
    40.08228, 40.21865, 40.35489, 40.49098, 40.62694, 40.76275, 40.89841, 
    41.03394, 41.16932, 41.30456, 41.43965, 41.57459, 41.70939, 41.84405, 
    41.97855, 42.11291, 42.24712, 42.38119, 42.5151,
  -18.32059, -18.20151, -18.08226, -17.96284, -17.84326, -17.72351, 
    -17.60359, -17.48351, -17.36325, -17.24283, -17.12225, -17.00149, 
    -16.88057, -16.75948, -16.63823, -16.5168, -16.39521, -16.27345, 
    -16.15153, -16.02944, -15.90718, -15.78475, -15.66216, -15.5394, 
    -15.41648, -15.29338, -15.17012, -15.0467, -14.9231, -14.79935, 
    -14.67542, -14.55133, -14.42707, -14.30265, -14.17806, -14.0533, 
    -13.92838, -13.80329, -13.67804, -13.55262, -13.42704, -13.30129, 
    -13.17538, -13.0493, -12.92306, -12.79666, -12.67008, -12.54335, 
    -12.41645, -12.28939, -12.16216, -12.03478, -11.90722, -11.77951, 
    -11.65163, -11.52359, -11.39539, -11.26702, -11.1385, -11.00981, 
    -10.88096, -10.75195, -10.62278, -10.49345, -10.36396, -10.2343, 
    -10.10449, -9.974521, -9.84439, -9.714101, -9.583652, -9.453046, 
    -9.322281, -9.19136, -9.06028, -8.929043, -8.797649, -8.6661, -8.534393, 
    -8.402532, -8.270514, -8.138342, -8.006015, -7.873534, -7.740899, 
    -7.60811, -7.475169, -7.342074, -7.208827, -7.075428, -6.941878, 
    -6.808176, -6.674324, -6.540321, -6.406168, -6.271867, -6.137415, 
    -6.002816, -5.868069, -5.733173, -5.598131, -5.462942, -5.327607, 
    -5.192126, -5.056499, -4.920729, -4.784813, -4.648755, -4.512553, 
    -4.376208, -4.239721, -4.103092, -3.966323, -3.829412, -3.692362, 
    -3.555173, -3.417844, -3.280378, -3.142773, -3.005032, -2.867153, 
    -2.729139, -2.59099, -2.452706, -2.314287, -2.175735, -2.03705, 
    -1.898233, -1.759284, -1.620205, -1.480995, -1.341655, -1.202186, 
    -1.062589, -0.9228637, -0.7830117, -0.6430333, -0.5029293, -0.3627003, 
    -0.222347, -0.08187011, 0.0587296, 0.1994514, 0.3402947, 0.4812587, 
    0.6223426, 0.7635457, 0.9048673, 1.046307, 1.187863, 1.329535, 1.471323, 
    1.613226, 1.755242, 1.897372, 2.039613, 2.181967, 2.324431, 2.467005, 
    2.609688, 2.752479, 2.895378, 3.038383, 3.181494, 3.32471, 3.46803, 
    3.611453, 3.754979, 3.898606, 4.042334, 4.186162, 4.330088, 4.474113, 
    4.618235, 4.762453, 4.906766, 5.051174, 5.195675, 5.340269, 5.484954, 
    5.629731, 5.774597, 5.919552, 6.064596, 6.209726, 6.354942, 6.500244, 
    6.645629, 6.791098, 6.936649, 7.082282, 7.227995, 7.373787, 7.519658, 
    7.665606, 7.811631, 7.95773, 8.103905, 8.250153, 8.396473, 8.542864, 
    8.689326, 8.835857, 8.982457, 9.129125, 9.275858, 9.422656, 9.569519, 
    9.716445, 9.863433, 10.01048, 10.15759, 10.30476, 10.45199, 10.59927, 
    10.74661, 10.894, 11.04145, 11.18895, 11.3365, 11.4841, 11.63175, 
    11.77945, 11.9272, 12.07499, 12.22283, 12.37071, 12.51864, 12.66661, 
    12.81461, 12.96266, 13.11074, 13.25887, 13.40703, 13.55522, 13.70345, 
    13.85171, 14, 14.14832, 14.29668, 14.44506, 14.59346, 14.7419, 14.89036, 
    15.03884, 15.18735, 15.33587, 15.48442, 15.63299, 15.78157, 15.93018, 
    16.0788, 16.22743, 16.37608, 16.52473, 16.6734, 16.82209, 16.97078, 
    17.11947, 17.26818, 17.41689, 17.5656, 17.71432, 17.86304, 18.01176, 
    18.16048, 18.3092, 18.45792, 18.60664, 18.75534, 18.90405, 19.05275, 
    19.20143, 19.35011, 19.49878, 19.64744, 19.79608, 19.94472, 20.09333, 
    20.24193, 20.39051, 20.53908, 20.68762, 20.83615, 20.98465, 21.13313, 
    21.28158, 21.43001, 21.57842, 21.72679, 21.87514, 22.02346, 22.17175, 
    22.32, 22.46822, 22.61641, 22.76457, 22.91268, 23.06076, 23.2088, 
    23.3568, 23.50476, 23.65268, 23.80056, 23.94839, 24.09617, 24.24391, 
    24.39161, 24.53925, 24.68684, 24.83439, 24.98188, 25.12932, 25.2767, 
    25.42403, 25.57131, 25.71852, 25.86568, 26.01278, 26.15982, 26.3068, 
    26.45372, 26.60057, 26.74736, 26.89408, 27.04074, 27.18733, 27.33385, 
    27.4803, 27.62668, 27.77299, 27.91922, 28.06539, 28.21147, 28.35748, 
    28.50342, 28.64928, 28.79506, 28.94076, 29.08638, 29.23192, 29.37737, 
    29.52275, 29.66804, 29.81324, 29.95835, 30.10338, 30.24833, 30.39318, 
    30.53794, 30.68261, 30.82719, 30.97168, 31.11607, 31.26037, 31.40457, 
    31.54868, 31.69268, 31.8366, 31.98041, 32.12412, 32.26773, 32.41124, 
    32.55465, 32.69795, 32.84115, 32.98425, 33.12724, 33.27011, 33.41289, 
    33.55556, 33.69811, 33.84056, 33.98289, 34.12512, 34.26723, 34.40923, 
    34.55111, 34.69288, 34.83454, 34.97607, 35.1175, 35.2588, 35.39998, 
    35.54105, 35.68199, 35.82281, 35.96352, 36.1041, 36.24456, 36.38489, 
    36.5251, 36.66518, 36.80514, 36.94497, 37.08468, 37.22425, 37.3637, 
    37.50303, 37.64221, 37.78127, 37.9202, 38.059, 38.19766, 38.33619, 
    38.47459, 38.61285, 38.75098, 38.88897, 39.02683, 39.16455, 39.30213, 
    39.43958, 39.57689, 39.71405, 39.85108, 39.98797, 40.12471, 40.26132, 
    40.39779, 40.53411, 40.67029, 40.80632, 40.94221, 41.07796, 41.21357, 
    41.34903, 41.48434, 41.6195, 41.75452, 41.88939, 42.02412, 42.1587, 
    42.29312, 42.4274, 42.56153,
  -18.38342, -18.2642, -18.14481, -18.02526, -17.90553, -17.78564, -17.66558, 
    -17.54536, -17.42496, -17.3044, -17.18367, -17.06277, -16.9417, 
    -16.82046, -16.69906, -16.57749, -16.45575, -16.33384, -16.21176, 
    -16.08952, -15.96711, -15.84453, -15.72178, -15.59887, -15.47578, 
    -15.35253, -15.22912, -15.10553, -14.98178, -14.85786, -14.73378, 
    -14.60952, -14.4851, -14.36051, -14.23576, -14.11084, -13.98575, 
    -13.8605, -13.73508, -13.6095, -13.48374, -13.35783, -13.23174, 
    -13.10549, -12.97908, -12.8525, -12.72576, -12.59885, -12.47177, 
    -12.34453, -12.21713, -12.08956, -11.96183, -11.83394, -11.70588, 
    -11.57766, -11.44927, -11.32073, -11.19201, -11.06314, -10.93411, 
    -10.80491, -10.67555, -10.54603, -10.41635, -10.28651, -10.1565, 
    -10.02634, -9.896018, -9.765535, -9.634892, -9.504091, -9.373131, 
    -9.242011, -9.110734, -8.979299, -8.847705, -8.715955, -8.584047, 
    -8.451983, -8.319764, -8.187387, -8.054856, -7.92217, -7.789328, 
    -7.656332, -7.523182, -7.389879, -7.256422, -7.122813, -6.989051, 
    -6.855137, -6.721071, -6.586854, -6.452487, -6.317969, -6.183302, 
    -6.048485, -5.913519, -5.778405, -5.643143, -5.507733, -5.372176, 
    -5.236472, -5.100623, -4.964628, -4.828487, -4.692203, -4.555774, 
    -4.419202, -4.282487, -4.145629, -4.008629, -3.871489, -3.734207, 
    -3.596785, -3.459223, -3.321522, -3.183683, -3.045706, -2.907591, 
    -2.76934, -2.630952, -2.492429, -2.353771, -2.214978, -2.076052, 
    -1.936993, -1.797801, -1.658478, -1.519023, -1.379438, -1.239723, 
    -1.099879, -0.9599065, -0.8198062, -0.6795787, -0.5392247, -0.398745, 
    -0.2581403, -0.1174113, 0.02344135, 0.1644169, 0.3055146, 0.4467337, 
    0.5880736, 0.7295333, 0.8711123, 1.01281, 1.154625, 1.296557, 1.438605, 
    1.580769, 1.723047, 1.865439, 2.007944, 2.150561, 2.293289, 2.436128, 
    2.579077, 2.722135, 2.865301, 3.008574, 3.151954, 3.295439, 3.439029, 
    3.582723, 3.72652, 3.870419, 4.014419, 4.15852, 4.30272, 4.447019, 
    4.591416, 4.735909, 4.880499, 5.025184, 5.169962, 5.314834, 5.459798, 
    5.604854, 5.75, 5.895236, 6.04056, 6.185971, 6.33147, 6.477054, 6.622723, 
    6.768476, 6.914311, 7.060228, 7.206226, 7.352304, 7.498461, 7.644696, 
    7.791008, 7.937396, 8.083858, 8.230395, 8.377005, 8.523685, 8.670438, 
    8.81726, 8.96415, 9.111109, 9.258134, 9.405225, 9.552381, 9.6996, 
    9.846882, 9.994226, 10.14163, 10.28909, 10.43661, 10.58419, 10.73183, 
    10.87952, 11.02726, 11.17506, 11.32291, 11.47081, 11.61876, 11.76675, 
    11.9148, 12.06289, 12.21103, 12.35921, 12.50744, 12.6557, 12.80401, 
    12.95236, 13.10074, 13.24917, 13.39763, 13.54612, 13.69465, 13.84321, 
    13.99181, 14.14044, 14.28909, 14.43777, 14.58648, 14.73522, 14.88399, 
    15.03277, 15.18158, 15.33041, 15.47926, 15.62814, 15.77703, 15.92593, 
    16.07486, 16.22379, 16.37274, 16.52171, 16.67068, 16.81967, 16.96866, 
    17.11767, 17.26668, 17.41569, 17.56471, 17.71374, 17.86276, 18.01179, 
    18.16081, 18.30984, 18.45886, 18.60788, 18.7569, 18.9059, 19.0549, 
    19.2039, 19.35288, 19.50186, 19.65082, 19.79977, 19.9487, 20.09762, 
    20.24653, 20.39541, 20.54428, 20.69313, 20.84196, 20.99076, 21.13955, 
    21.28831, 21.43704, 21.58575, 21.73443, 21.88308, 22.0317, 22.18029, 
    22.32885, 22.47737, 22.62586, 22.77431, 22.92273, 23.07111, 23.21945, 
    23.36775, 23.51601, 23.66423, 23.81241, 23.96054, 24.10862, 24.25666, 
    24.40465, 24.55259, 24.70048, 24.84832, 24.99611, 25.14385, 25.29153, 
    25.43916, 25.58673, 25.73424, 25.88169, 26.02909, 26.17642, 26.32369, 
    26.4709, 26.61805, 26.76513, 26.91214, 27.05909, 27.20597, 27.35278, 
    27.49952, 27.64619, 27.79279, 27.93931, 28.08577, 28.23214, 28.37844, 
    28.52466, 28.67081, 28.81687, 28.96286, 29.10876, 29.25459, 29.40033, 
    29.54598, 29.69155, 29.83704, 29.98243, 30.12774, 30.27297, 30.4181, 
    30.56314, 30.70809, 30.85295, 30.99771, 31.14238, 31.28695, 31.43143, 
    31.57581, 31.7201, 31.86428, 32.00837, 32.15235, 32.29623, 32.44001, 
    32.58369, 32.72726, 32.87074, 33.0141, 33.15735, 33.3005, 33.44354, 
    33.58648, 33.72929, 33.87201, 34.01461, 34.15709, 34.29947, 34.44173, 
    34.58387, 34.7259, 34.86782, 35.00961, 35.15129, 35.29285, 35.43429, 
    35.57561, 35.71681, 35.85789, 35.99885, 36.13968, 36.28039, 36.42097, 
    36.56144, 36.70177, 36.84198, 36.98206, 37.12201, 37.26183, 37.40153, 
    37.54109, 37.68053, 37.81983, 37.959, 38.09804, 38.23694, 38.37571, 
    38.51435, 38.65285, 38.79122, 38.92945, 39.06754, 39.2055, 39.34332, 
    39.48099, 39.61853, 39.75593, 39.89319, 40.03031, 40.16729, 40.30412, 
    40.44081, 40.57737, 40.71377, 40.85003, 40.98615, 41.12212, 41.25795, 
    41.39363, 41.52916, 41.66455, 41.79979, 41.93488, 42.06982, 42.20461, 
    42.33926, 42.47375, 42.6081,
  -18.44641, -18.32705, -18.20752, -18.08783, -17.96797, -17.84793, 
    -17.72773, -17.60736, -17.48682, -17.36612, -17.24524, -17.12419, 
    -17.00298, -16.8816, -16.76004, -16.63832, -16.51643, -16.39438, 
    -16.27215, -16.14975, -16.02719, -15.90446, -15.78156, -15.65849, 
    -15.53525, -15.41184, -15.28827, -15.16452, -15.04061, -14.91653, 
    -14.79229, -14.66787, -14.54329, -14.41854, -14.29362, -14.16853, 
    -14.04328, -13.91786, -13.79228, -13.66652, -13.5406, -13.41451, 
    -13.28826, -13.16184, -13.03525, -12.9085, -12.78158, -12.6545, 
    -12.52725, -12.39983, -12.27225, -12.1445, -12.01659, -11.88852, 
    -11.76028, -11.63188, -11.50331, -11.37458, -11.24568, -11.11662, 
    -10.9874, -10.85802, -10.72847, -10.59876, -10.46889, -10.33886, 
    -10.20867, -10.07831, -9.947796, -9.81712, -9.686282, -9.555285, 
    -9.424128, -9.292811, -9.161336, -9.029701, -8.897908, -8.765958, 
    -8.633848, -8.501582, -8.369159, -8.236579, -8.103843, -7.97095, 
    -7.837902, -7.704699, -7.57134, -7.437827, -7.304161, -7.17034, 
    -7.036366, -6.902239, -6.767961, -6.633529, -6.498947, -6.364213, 
    -6.229328, -6.094294, -5.959109, -5.823775, -5.688293, -5.552661, 
    -5.416883, -5.280956, -5.144883, -5.008663, -4.872298, -4.735786, 
    -4.599131, -4.46233, -4.325387, -4.188299, -4.051069, -3.913697, 
    -3.776183, -3.638528, -3.500733, -3.362797, -3.224723, -3.086509, 
    -2.948157, -2.809668, -2.671042, -2.532279, -2.393381, -2.254347, 
    -2.115179, -1.975877, -1.836442, -1.696874, -1.557175, -1.417344, 
    -1.277382, -1.137291, -0.9970698, -0.8567205, -0.7162432, -0.5756387, 
    -0.4349077, -0.294051, -0.1530691, -0.01196284, 0.1292671, 0.2706199, 
    0.4120948, 0.5536913, 0.6954084, 0.8372455, 0.9792017, 1.121276, 
    1.263469, 1.405778, 1.548203, 1.690744, 1.833399, 1.976168, 2.119049, 
    2.262043, 2.405148, 2.548363, 2.691689, 2.835123, 2.978664, 3.122313, 
    3.266069, 3.40993, 3.553895, 3.697963, 3.842135, 3.986409, 4.130784, 
    4.275259, 4.419833, 4.564505, 4.709275, 4.854142, 4.999104, 5.144161, 
    5.289312, 5.434556, 5.579891, 5.725318, 5.870835, 6.016441, 6.162135, 
    6.307916, 6.453784, 6.599737, 6.745774, 6.891895, 7.038098, 7.184382, 
    7.330747, 7.477191, 7.623713, 7.770314, 7.91699, 8.063742, 8.210568, 
    8.357468, 8.504439, 8.651483, 8.798596, 8.94578, 9.09303, 9.240349, 
    9.387733, 9.535182, 9.682695, 9.830273, 9.977911, 10.12561, 10.27337, 
    10.42119, 10.56906, 10.71699, 10.86498, 11.01302, 11.16112, 11.30927, 
    11.45746, 11.60571, 11.75401, 11.90236, 12.05075, 12.19918, 12.34767, 
    12.49619, 12.64476, 12.79337, 12.94202, 13.09071, 13.23943, 13.3882, 
    13.53699, 13.68583, 13.83469, 13.98359, 14.13252, 14.28148, 14.43046, 
    14.57948, 14.72852, 14.87759, 15.02668, 15.17579, 15.32493, 15.47409, 
    15.62326, 15.77246, 15.92167, 16.0709, 16.22014, 16.3694, 16.51867, 
    16.66795, 16.81724, 16.96655, 17.11585, 17.26517, 17.41449, 17.56382, 
    17.71315, 17.86248, 18.01181, 18.16114, 18.31047, 18.4598, 18.60913, 
    18.75845, 18.90776, 19.05707, 19.20637, 19.35566, 19.50494, 19.65421, 
    19.80346, 19.95271, 20.10193, 20.25114, 20.40033, 20.54951, 20.69866, 
    20.84779, 20.9969, 21.14599, 21.29506, 21.44409, 21.59311, 21.74209, 
    21.89104, 22.03997, 22.18886, 22.33772, 22.48655, 22.63534, 22.7841, 
    22.93282, 23.0815, 23.23014, 23.37874, 23.52731, 23.67582, 23.8243, 
    23.97273, 24.12111, 24.26945, 24.41774, 24.56598, 24.71417, 24.86231, 
    25.0104, 25.15843, 25.30641, 25.45433, 25.6022, 25.75001, 25.89776, 
    26.04545, 26.19308, 26.34064, 26.48815, 26.63559, 26.78296, 26.93027, 
    27.07751, 27.22468, 27.37178, 27.51881, 27.66577, 27.81266, 27.95948, 
    28.10622, 28.25288, 28.39947, 28.54598, 28.69241, 28.83876, 28.98503, 
    29.13123, 29.27733, 29.42336, 29.5693, 29.71515, 29.86092, 30.0066, 
    30.15219, 30.29769, 30.4431, 30.58843, 30.73365, 30.87879, 31.02383, 
    31.16878, 31.31363, 31.45839, 31.60304, 31.7476, 31.89206, 32.03642, 
    32.18068, 32.32483, 32.46888, 32.61283, 32.75668, 32.90042, 33.04405, 
    33.18757, 33.33099, 33.4743, 33.6175, 33.76058, 33.90356, 34.04642, 
    34.18917, 34.33181, 34.47433, 34.61674, 34.75903, 34.90121, 35.04326, 
    35.1852, 35.32702, 35.46872, 35.61029, 35.75175, 35.89308, 36.03429, 
    36.17538, 36.31634, 36.45718, 36.59789, 36.73847, 36.87893, 37.01926, 
    37.15946, 37.29953, 37.43947, 37.57928, 37.71896, 37.85851, 37.99792, 
    38.1372, 38.27635, 38.41536, 38.55424, 38.69298, 38.83158, 38.97005, 
    39.10838, 39.24657, 39.38462, 39.52254, 39.66031, 39.79795, 39.93544, 
    40.07279, 40.21, 40.34706, 40.48398, 40.62076, 40.75739, 40.89388, 
    41.03022, 41.16642, 41.30247, 41.43837, 41.57413, 41.70973, 41.84519, 
    41.9805, 42.11567, 42.25068, 42.38554, 42.52024, 42.6548,
  -18.50955, -18.39005, -18.27039, -18.15055, -18.03055, -17.91038, 
    -17.79004, -17.66952, -17.54884, -17.42799, -17.30697, -17.18578, 
    -17.06442, -16.94289, -16.82119, -16.69932, -16.57728, -16.45507, 
    -16.33269, -16.21014, -16.08743, -15.96454, -15.84149, -15.71826, 
    -15.59487, -15.4713, -15.34757, -15.22367, -15.0996, -14.97536, 
    -14.85095, -14.72638, -14.60163, -14.47672, -14.35163, -14.22638, 
    -14.10097, -13.97538, -13.84962, -13.7237, -13.59761, -13.47135, 
    -13.34493, -13.21834, -13.09158, -12.96465, -12.83756, -12.7103, 
    -12.58287, -12.45528, -12.32752, -12.1996, -12.07151, -11.94325, 
    -11.81483, -11.68625, -11.5575, -11.42858, -11.2995, -11.17026, 
    -11.04085, -10.91128, -10.78155, -10.65165, -10.52159, -10.39137, 
    -10.26098, -10.13043, -9.999723, -9.868853, -9.737821, -9.606627, 
    -9.475274, -9.34376, -9.212087, -9.080253, -8.948259, -8.816108, 
    -8.683797, -8.551328, -8.418701, -8.285916, -8.152975, -8.019876, 
    -7.886621, -7.75321, -7.619643, -7.48592, -7.352043, -7.218011, 
    -7.083825, -6.949485, -6.814992, -6.680346, -6.545548, -6.410598, 
    -6.275496, -6.140243, -6.004839, -5.869285, -5.733582, -5.597729, 
    -5.461728, -5.325578, -5.189281, -5.052835, -4.916244, -4.779507, 
    -4.642623, -4.505594, -4.368421, -4.231104, -4.093643, -3.956039, 
    -3.818292, -3.680404, -3.542374, -3.404204, -3.265893, -3.127443, 
    -2.988853, -2.850126, -2.71126, -2.572258, -2.433118, -2.293843, 
    -2.154433, -2.014887, -1.875208, -1.735395, -1.59545, -1.455373, 
    -1.315164, -1.174824, -1.034354, -0.8937555, -0.7530278, -0.6121721, 
    -0.4711892, -0.3300797, -0.1888443, -0.04748377, 0.09400116, 0.2356098, 
    0.3773413, 0.519195, 0.6611702, 0.803266, 0.9454818, 1.087817, 1.23027, 
    1.372841, 1.515529, 1.658332, 1.801251, 1.944285, 2.087432, 2.230692, 
    2.374063, 2.517546, 2.661139, 2.804842, 2.948654, 3.092573, 3.236599, 
    3.380731, 3.524968, 3.66931, 3.813756, 3.958303, 4.102952, 4.247703, 
    4.392553, 4.537502, 4.68255, 4.827694, 4.972935, 5.118271, 5.263702, 
    5.409226, 5.554843, 5.700551, 5.84635, 5.992239, 6.138216, 6.284281, 
    6.430433, 6.576671, 6.722994, 6.869401, 7.01589, 7.162462, 7.309114, 
    7.455846, 7.602658, 7.749547, 7.896513, 8.043555, 8.190672, 8.337863, 
    8.485126, 8.632462, 8.779868, 8.927343, 9.074888, 9.2225, 9.370179, 
    9.517923, 9.665731, 9.813604, 9.961538, 10.10953, 10.25759, 10.4057, 
    10.55388, 10.70211, 10.85039, 10.99873, 11.14713, 11.29558, 11.44407, 
    11.59262, 11.74122, 11.88986, 12.03856, 12.1873, 12.33608, 12.48491, 
    12.63378, 12.78269, 12.93164, 13.08063, 13.22966, 13.37873, 13.52783, 
    13.67697, 13.82614, 13.97534, 14.12457, 14.27384, 14.42313, 14.57245, 
    14.7218, 14.87117, 15.02057, 15.16999, 15.31943, 15.46889, 15.61838, 
    15.76788, 15.9174, 16.06693, 16.21648, 16.36604, 16.51562, 16.66521, 
    16.81481, 16.96442, 17.11403, 17.26366, 17.41329, 17.56292, 17.71256, 
    17.8622, 18.01184, 18.16148, 18.31111, 18.46075, 18.61038, 18.76001, 
    18.90963, 19.05925, 19.20885, 19.35845, 19.50804, 19.65761, 19.80718, 
    19.95672, 20.10626, 20.25577, 20.40527, 20.55475, 20.70421, 20.85365, 
    21.00307, 21.15246, 21.30183, 21.45117, 21.60049, 21.74978, 21.89903, 
    22.04826, 22.19746, 22.34663, 22.49576, 22.64485, 22.79391, 22.94294, 
    23.09192, 23.24087, 23.38977, 23.53864, 23.68746, 23.83623, 23.98497, 
    24.13365, 24.28229, 24.43088, 24.57942, 24.72791, 24.87635, 25.02473, 
    25.17307, 25.32134, 25.46956, 25.61773, 25.76583, 25.91388, 26.06187, 
    26.20979, 26.35765, 26.50545, 26.65318, 26.80085, 26.94846, 27.09599, 
    27.24345, 27.39085, 27.53817, 27.68542, 27.83261, 27.97971, 28.12674, 
    28.27369, 28.42057, 28.56737, 28.71409, 28.86073, 29.00729, 29.15376, 
    29.30016, 29.44647, 29.59269, 29.73883, 29.88488, 30.03084, 30.17672, 
    30.3225, 30.4682, 30.6138, 30.75931, 30.90472, 31.05005, 31.19527, 
    31.3404, 31.48543, 31.63037, 31.7752, 31.91994, 32.06457, 32.2091, 
    32.35353, 32.49786, 32.64207, 32.78619, 32.9302, 33.0741, 33.2179, 
    33.36158, 33.50516, 33.64862, 33.79198, 33.93522, 34.07835, 34.22136, 
    34.36427, 34.50705, 34.64972, 34.79227, 34.93471, 35.07702, 35.21922, 
    35.3613, 35.50325, 35.64509, 35.7868, 35.92839, 36.06985, 36.21119, 
    36.35241, 36.4935, 36.63446, 36.7753, 36.916, 37.05658, 37.19703, 
    37.33735, 37.47754, 37.6176, 37.75752, 37.89731, 38.03697, 38.17649, 
    38.31588, 38.45514, 38.59425, 38.73323, 38.87208, 39.01078, 39.14935, 
    39.28778, 39.42607, 39.56422, 39.70222, 39.84009, 39.97781, 40.11539, 
    40.25283, 40.39013, 40.52728, 40.66428, 40.80115, 40.93786, 41.07443, 
    41.21085, 41.34713, 41.48325, 41.61923, 41.75506, 41.89074, 42.02627, 
    42.16165, 42.29688, 42.43195, 42.56688, 42.70166,
  -18.57285, -18.45321, -18.33341, -18.21344, -18.09329, -17.97298, -17.8525, 
    -17.73184, -17.61102, -17.49002, -17.36885, -17.24752, -17.12601, 
    -17.00433, -16.88249, -16.76047, -16.63828, -16.51592, -16.39339, 
    -16.27069, -16.14782, -16.02478, -15.90157, -15.77819, -15.65464, 
    -15.53092, -15.40703, -15.28297, -15.15874, -15.03434, -14.90978, 
    -14.78504, -14.66013, -14.53505, -14.40981, -14.28439, -14.15881, 
    -14.03305, -13.90713, -13.78104, -13.65478, -13.52835, -13.40176, 
    -13.27499, -13.14806, -13.02096, -12.89369, -12.76626, -12.63866, 
    -12.51089, -12.38295, -12.25485, -12.12658, -11.99814, -11.86954, 
    -11.74077, -11.61184, -11.48274, -11.35348, -11.22405, -11.09445, 
    -10.9647, -10.83477, -10.70469, -10.57444, -10.44402, -10.31345, 
    -10.18271, -10.0518, -9.920737, -9.789511, -9.658121, -9.52657, 
    -9.394859, -9.262986, -9.130953, -8.99876, -8.866406, -8.733894, 
    -8.601222, -8.468391, -8.335402, -8.202254, -8.06895, -7.935487, 
    -7.801867, -7.668091, -7.534159, -7.40007, -7.265827, -7.131428, 
    -6.996875, -6.862168, -6.727306, -6.592292, -6.457125, -6.321805, 
    -6.186334, -6.05071, -5.914936, -5.779012, -5.642937, -5.506712, 
    -5.370339, -5.233817, -5.097147, -4.960329, -4.823364, -4.686252, 
    -4.548995, -4.411592, -4.274044, -4.136351, -3.998515, -3.860535, 
    -3.722413, -3.584148, -3.445742, -3.307195, -3.168507, -3.02968, 
    -2.890713, -2.751608, -2.612365, -2.472984, -2.333466, -2.193813, 
    -2.054024, -1.9141, -1.774042, -1.63385, -1.493525, -1.353069, -1.21248, 
    -1.071761, -0.930912, -0.7899333, -0.6488258, -0.5075902, -0.3662273, 
    -0.2247377, -0.08312225, 0.05861839, 0.2004835, 0.3424723, 0.484584, 
    0.6268179, 0.7691733, 0.9116493, 1.054245, 1.19696, 1.339794, 1.482744, 
    1.625812, 1.768996, 1.912295, 2.055708, 2.199234, 2.342873, 2.486624, 
    2.630487, 2.774459, 2.918541, 3.062731, 3.207029, 3.351433, 3.495944, 
    3.640559, 3.785278, 3.930101, 4.075026, 4.220053, 4.36518, 4.510407, 
    4.655732, 4.801156, 4.946676, 5.092292, 5.238003, 5.383809, 5.529707, 
    5.675698, 5.82178, 5.967952, 6.114213, 6.260564, 6.407001, 6.553525, 
    6.700134, 6.846828, 6.993605, 7.140464, 7.287405, 7.434427, 7.581528, 
    7.728707, 7.875964, 8.023297, 8.170706, 8.318189, 8.465745, 8.613373, 
    8.761073, 8.908843, 9.056682, 9.204589, 9.352563, 9.500603, 9.648707, 
    9.796876, 9.945107, 10.0934, 10.24175, 10.39017, 10.53864, 10.68717, 
    10.83575, 10.98439, 11.13309, 11.28184, 11.43063, 11.57948, 11.72838, 
    11.87733, 12.02633, 12.17537, 12.32445, 12.47359, 12.62276, 12.77197, 
    12.92123, 13.07052, 13.21986, 13.36923, 13.51864, 13.66808, 13.81755, 
    13.96706, 14.1166, 14.26617, 14.41577, 14.5654, 14.71505, 14.86473, 
    15.01443, 15.16416, 15.31391, 15.46368, 15.61347, 15.76328, 15.91311, 
    16.06295, 16.21281, 16.36268, 16.51256, 16.66246, 16.81237, 16.96228, 
    17.11221, 17.26214, 17.41208, 17.56202, 17.71196, 17.86191, 18.01186, 
    18.16181, 18.31176, 18.4617, 18.61164, 18.76158, 18.91151, 19.06143, 
    19.21135, 19.36125, 19.51115, 19.66103, 19.8109, 19.96076, 20.1106, 
    20.26042, 20.41023, 20.56001, 20.70978, 20.85953, 21.00925, 21.15895, 
    21.30863, 21.45827, 21.6079, 21.75749, 21.90706, 22.05659, 22.20609, 
    22.35556, 22.505, 22.6544, 22.80377, 22.95309, 23.10238, 23.25163, 
    23.40084, 23.55001, 23.69913, 23.84821, 23.99725, 24.14623, 24.29517, 
    24.44407, 24.59291, 24.7417, 24.89044, 25.03912, 25.18775, 25.33633, 
    25.48485, 25.63331, 25.78172, 25.93006, 26.07834, 26.22657, 26.37473, 
    26.52282, 26.67085, 26.81881, 26.96671, 27.11454, 27.26229, 27.40998, 
    27.5576, 27.70514, 27.85262, 28.00001, 28.14734, 28.29458, 28.44175, 
    28.58883, 28.73584, 28.88277, 29.02962, 29.17638, 29.32306, 29.46966, 
    29.61617, 29.76259, 29.90893, 30.05518, 30.20133, 30.3474, 30.49338, 
    30.63926, 30.78505, 30.93075, 31.07635, 31.22186, 31.36726, 31.51257, 
    31.65778, 31.80289, 31.9479, 32.09282, 32.23762, 32.38232, 32.52692, 
    32.67142, 32.8158, 32.96009, 33.10426, 33.24832, 33.39228, 33.53612, 
    33.67986, 33.82348, 33.96698, 34.11038, 34.25366, 34.39683, 34.53988, 
    34.68281, 34.82562, 34.96832, 35.1109, 35.25335, 35.39569, 35.5379, 
    35.68, 35.82196, 35.96381, 36.10553, 36.24713, 36.3886, 36.52994, 
    36.67115, 36.81224, 36.9532, 37.09403, 37.23473, 37.37529, 37.51573, 
    37.65604, 37.79621, 37.93624, 38.07615, 38.21591, 38.35555, 38.49504, 
    38.6344, 38.77362, 38.9127, 39.05165, 39.19046, 39.32912, 39.46764, 
    39.60603, 39.74427, 39.88237, 40.02033, 40.15814, 40.29581, 40.43333, 
    40.57072, 40.70795, 40.84504, 40.98198, 41.11877, 41.25542, 41.39192, 
    41.52827, 41.66447, 41.80052, 41.93642, 42.07217, 42.20777, 42.34322, 
    42.47852, 42.61366, 42.74865,
  -18.6363, -18.51653, -18.39659, -18.27648, -18.15619, -18.03574, -17.91512, 
    -17.79432, -17.67335, -17.55221, -17.4309, -17.30942, -17.18776, 
    -17.06594, -16.94394, -16.82178, -16.69944, -16.57693, -16.45425, 
    -16.3314, -16.20838, -16.08518, -15.96182, -15.83828, -15.71458, 
    -15.5907, -15.46665, -15.34243, -15.21805, -15.09349, -14.96876, 
    -14.84386, -14.71879, -14.59354, -14.46813, -14.34255, -14.2168, 
    -14.09088, -13.96479, -13.83853, -13.7121, -13.58551, -13.45874, 
    -13.3318, -13.2047, -13.07743, -12.94998, -12.82237, -12.69459, 
    -12.56665, -12.43853, -12.31025, -12.1818, -12.05319, -11.9244, 
    -11.79545, -11.66634, -11.53706, -11.40761, -11.27799, -11.14821, 
    -11.01826, -10.88815, -10.75788, -10.62744, -10.49683, -10.36606, 
    -10.23513, -10.10403, -9.972775, -9.841352, -9.709766, -9.578018, 
    -9.446109, -9.314037, -9.181804, -9.04941, -8.916855, -8.78414, 
    -8.651265, -8.518229, -8.385036, -8.251682, -8.11817, -7.9845, -7.850672, 
    -7.716686, -7.582543, -7.448244, -7.313788, -7.179177, -7.04441, 
    -6.909488, -6.774411, -6.63918, -6.503796, -6.368258, -6.232567, 
    -6.096724, -5.960729, -5.824583, -5.688285, -5.551837, -5.415239, 
    -5.278492, -5.141596, -5.004551, -4.867359, -4.730019, -4.592532, 
    -4.454898, -4.317119, -4.179195, -4.041126, -3.902912, -3.764555, 
    -3.626056, -3.487413, -3.348629, -3.209704, -3.070637, -2.931431, 
    -2.792086, -2.652601, -2.512979, -2.373218, -2.233321, -2.093287, 
    -1.953118, -1.812814, -1.672375, -1.531803, -1.391098, -1.25026, 
    -1.109291, -0.9681909, -0.8269604, -0.6856005, -0.5441116, -0.4024946, 
    -0.2607502, -0.1188791, 0.02311794, 0.1652402, 0.3074869, 0.4498573, 
    0.5923507, 0.7349663, 0.8777032, 1.020561, 1.163538, 1.306635, 1.44985, 
    1.593182, 1.736631, 1.880196, 2.023876, 2.16767, 2.311578, 2.455598, 
    2.59973, 2.743972, 2.888325, 3.032787, 3.177357, 3.322035, 3.466819, 
    3.611709, 3.756703, 3.901802, 4.047004, 4.192307, 4.337712, 4.483217, 
    4.628822, 4.774525, 4.920325, 5.066223, 5.212215, 5.358303, 5.504484, 
    5.650758, 5.797124, 5.943581, 6.090127, 6.236763, 6.383487, 6.530297, 
    6.677194, 6.824175, 6.971241, 7.11839, 7.26562, 7.412932, 7.560323, 
    7.707794, 7.855342, 8.002968, 8.150669, 8.298445, 8.446295, 8.594217, 
    8.742211, 8.890276, 9.03841, 9.186614, 9.334884, 9.483221, 9.631623, 
    9.780089, 9.928618, 10.07721, 10.22586, 10.37458, 10.52335, 10.67218, 
    10.82106, 10.97, 11.119, 11.26805, 11.41715, 11.5663, 11.7155, 11.86475, 
    12.01405, 12.16339, 12.31279, 12.46222, 12.6117, 12.76122, 12.91078, 
    13.06038, 13.21002, 13.35969, 13.50941, 13.65915, 13.80894, 13.95875, 
    14.1086, 14.25847, 14.40838, 14.55831, 14.70828, 14.85826, 15.00828, 
    15.15831, 15.30837, 15.45845, 15.60855, 15.75866, 15.9088, 16.05895, 
    16.20912, 16.3593, 16.50949, 16.6597, 16.80992, 16.96014, 17.11037, 
    17.26062, 17.41086, 17.56111, 17.71137, 17.86163, 18.01188, 18.16214, 
    18.3124, 18.46265, 18.6129, 18.76315, 18.91339, 19.06362, 19.21385, 
    19.36406, 19.51427, 19.66446, 19.81464, 19.9648, 20.11495, 20.26508, 
    20.4152, 20.56529, 20.71537, 20.86543, 21.01546, 21.16546, 21.31545, 
    21.4654, 21.61533, 21.76524, 21.91511, 22.06495, 22.21476, 22.36454, 
    22.51428, 22.66398, 22.81366, 22.96329, 23.11288, 23.26244, 23.41195, 
    23.56142, 23.71085, 23.86023, 24.00957, 24.15886, 24.3081, 24.4573, 
    24.60644, 24.75554, 24.90458, 25.05356, 25.20249, 25.35137, 25.50019, 
    25.64895, 25.79766, 25.9463, 26.09488, 26.2434, 26.39186, 26.54025, 
    26.68857, 26.83683, 26.98503, 27.13315, 27.2812, 27.42919, 27.5771, 
    27.72494, 27.8727, 28.02039, 28.168, 28.31554, 28.463, 28.61038, 
    28.75768, 28.90489, 29.05203, 29.19908, 29.34605, 29.49293, 29.63973, 
    29.78644, 29.93306, 30.07959, 30.22603, 30.37239, 30.51865, 30.66481, 
    30.81088, 30.95686, 31.10275, 31.24853, 31.39422, 31.53981, 31.6853, 
    31.83068, 31.97597, 32.12116, 32.26624, 32.41122, 32.55609, 32.70086, 
    32.84552, 32.99007, 33.13452, 33.27885, 33.42308, 33.56719, 33.71119, 
    33.85508, 33.99886, 34.14252, 34.28607, 34.4295, 34.57281, 34.71601, 
    34.85909, 35.00204, 35.14488, 35.2876, 35.4302, 35.57267, 35.71502, 
    35.85725, 35.99935, 36.14133, 36.28318, 36.4249, 36.5665, 36.70797, 
    36.84931, 36.99052, 37.1316, 37.27255, 37.41336, 37.55405, 37.6946, 
    37.83502, 37.9753, 38.11545, 38.25546, 38.39534, 38.53507, 38.67467, 
    38.81414, 38.95346, 39.09264, 39.23169, 39.37059, 39.50935, 39.64797, 
    39.78645, 39.92479, 40.06298, 40.20102, 40.33892, 40.47668, 40.61429, 
    40.75175, 40.88907, 41.02624, 41.16326, 41.30013, 41.43686, 41.57343, 
    41.70985, 41.84613, 41.98225, 42.11822, 42.25404, 42.38971, 42.52522, 
    42.66058, 42.79579,
  -18.69992, -18.58001, -18.45993, -18.33968, -18.21925, -18.09866, 
    -17.97789, -17.85695, -17.73584, -17.61456, -17.4931, -17.37148, 
    -17.24968, -17.1277, -17.00556, -16.88325, -16.76076, -16.6381, 
    -16.51527, -16.39226, -16.26909, -16.14574, -16.02222, -15.89853, 
    -15.77467, -15.65064, -15.52643, -15.40205, -15.27751, -15.15279, 
    -15.0279, -14.90283, -14.7776, -14.6522, -14.52662, -14.40088, -14.27496, 
    -14.14887, -14.02261, -13.89618, -13.76959, -13.64282, -13.51588, 
    -13.38877, -13.26149, -13.13405, -13.00643, -12.87864, -12.75069, 
    -12.62257, -12.49427, -12.36581, -12.23718, -12.10839, -11.97942, 
    -11.85029, -11.72099, -11.59152, -11.46189, -11.33209, -11.20212, 
    -11.07199, -10.94169, -10.81122, -10.68059, -10.5498, -10.41883, 
    -10.28771, -10.15642, -10.02496, -9.893345, -9.761563, -9.629618, 
    -9.49751, -9.365239, -9.232806, -9.100211, -8.967455, -8.834537, 
    -8.701458, -8.568218, -8.434818, -8.301259, -8.16754, -8.033661, 
    -7.899624, -7.765429, -7.631075, -7.496564, -7.361897, -7.227071, 
    -7.09209, -6.956953, -6.821661, -6.686213, -6.55061, -6.414854, 
    -6.278944, -6.14288, -6.006664, -5.870296, -5.733775, -5.597104, 
    -5.460281, -5.323308, -5.186186, -5.048913, -4.911493, -4.773924, 
    -4.636207, -4.498343, -4.360332, -4.222175, -4.083873, -3.945425, 
    -3.806833, -3.668097, -3.529218, -3.390197, -3.251033, -3.111727, 
    -2.972281, -2.832695, -2.692968, -2.553103, -2.4131, -2.272958, 
    -2.132679, -1.992264, -1.851713, -1.711027, -1.570207, -1.429252, 
    -1.288165, -1.146945, -1.005593, -0.8641102, -0.722497, -0.5807542, 
    -0.4388825, -0.2968825, -0.1547551, -0.01250102, 0.1298791, 0.2723844, 
    0.4150143, 0.5577678, 0.7006443, 0.843643, 0.9867631, 1.130004, 1.273364, 
    1.416844, 1.560442, 1.704157, 1.847988, 1.991936, 2.135998, 2.280175, 
    2.424465, 2.568867, 2.713381, 2.858006, 3.00274, 3.147584, 3.292535, 
    3.437594, 3.582759, 3.72803, 3.873405, 4.018884, 4.164466, 4.310149, 
    4.455934, 4.601818, 4.747802, 4.893883, 5.040062, 5.186337, 5.332708, 
    5.479173, 5.625731, 5.772382, 5.919124, 6.065957, 6.212879, 6.35989, 
    6.506989, 6.654173, 6.801444, 6.948799, 7.096237, 7.243758, 7.391361, 
    7.539044, 7.686807, 7.834648, 7.982566, 8.130561, 8.278631, 8.426775, 
    8.574993, 8.723283, 8.871643, 9.020074, 9.168574, 9.317142, 9.465776, 
    9.614477, 9.763242, 9.91207, 10.06096, 10.20991, 10.35893, 10.508, 
    10.65713, 10.80632, 10.95556, 11.10486, 11.25421, 11.40361, 11.55307, 
    11.70257, 11.85213, 12.00173, 12.15138, 12.30107, 12.45081, 12.6006, 
    12.75042, 12.90029, 13.0502, 13.20014, 13.35013, 13.50014, 13.6502, 
    13.80029, 13.95041, 14.10057, 14.25075, 14.40097, 14.55121, 14.70148, 
    14.85177, 15.0021, 15.15244, 15.30281, 15.4532, 15.6036, 15.75403, 
    15.90448, 16.05494, 16.20542, 16.35591, 16.50641, 16.65693, 16.80746, 
    16.95799, 17.10854, 17.25909, 17.40965, 17.56021, 17.71077, 17.86134, 
    18.01191, 18.16248, 18.31305, 18.46361, 18.61417, 18.76473, 18.91528, 
    19.06582, 19.21636, 19.36688, 19.5174, 19.6679, 19.81839, 19.96886, 
    20.11932, 20.26977, 20.42019, 20.57059, 20.72098, 20.87134, 21.02168, 
    21.172, 21.32229, 21.47256, 21.6228, 21.77301, 21.92319, 22.07334, 
    22.22346, 22.37354, 22.52359, 22.6736, 22.82358, 22.97352, 23.12342, 
    23.27328, 23.4231, 23.57288, 23.72261, 23.8723, 24.02194, 24.17153, 
    24.32108, 24.47058, 24.62003, 24.76942, 24.91876, 25.06805, 25.21729, 
    25.36646, 25.51558, 25.66465, 25.81365, 25.96259, 26.11147, 26.26029, 
    26.40905, 26.55774, 26.70636, 26.85492, 27.00341, 27.15183, 27.30018, 
    27.44846, 27.59666, 27.7448, 27.89285, 28.04084, 28.18874, 28.33657, 
    28.48432, 28.63199, 28.77958, 28.92709, 29.07452, 29.22186, 29.36912, 
    29.51629, 29.66337, 29.81037, 29.95728, 30.10409, 30.25082, 30.39746, 
    30.544, 30.69045, 30.83681, 30.98307, 31.12923, 31.2753, 31.42126, 
    31.56713, 31.7129, 31.85857, 32.00414, 32.1496, 32.29496, 32.44021, 
    32.58536, 32.7304, 32.87534, 33.02016, 33.16488, 33.30949, 33.45398, 
    33.59837, 33.74264, 33.8868, 34.03084, 34.17477, 34.31858, 34.46228, 
    34.60586, 34.74932, 34.89266, 35.03588, 35.17899, 35.32196, 35.46482, 
    35.60756, 35.75017, 35.89265, 36.03501, 36.17725, 36.31936, 36.46133, 
    36.60318, 36.74491, 36.8865, 37.02796, 37.16929, 37.31049, 37.45156, 
    37.59249, 37.73329, 37.87395, 38.01448, 38.15488, 38.29514, 38.43526, 
    38.57524, 38.71508, 38.85479, 38.99435, 39.13377, 39.27306, 39.4122, 
    39.5512, 39.69005, 39.82877, 39.96733, 40.10576, 40.24404, 40.38217, 
    40.52016, 40.658, 40.7957, 40.93324, 41.07064, 41.20789, 41.34499, 
    41.48193, 41.61873, 41.75538, 41.89188, 42.02822, 42.16441, 42.30045, 
    42.43634, 42.57207, 42.70765, 42.84307,
  -18.76369, -18.64364, -18.52343, -18.40303, -18.28247, -18.16174, 
    -18.04083, -17.91975, -17.79849, -17.67706, -17.55546, -17.43369, 
    -17.31175, -17.18963, -17.06734, -16.94487, -16.82224, -16.69943, 
    -16.57644, -16.45329, -16.32996, -16.20646, -16.08279, -15.95894, 
    -15.83492, -15.71073, -15.58637, -15.46183, -15.33713, -15.21225, 
    -15.08719, -14.96197, -14.83657, -14.71101, -14.58527, -14.45936, 
    -14.33327, -14.20702, -14.08059, -13.954, -13.82723, -13.70029, 
    -13.57318, -13.4459, -13.31845, -13.19083, -13.06304, -12.93507, 
    -12.80694, -12.67864, -12.55017, -12.42153, -12.29272, -12.16374, 
    -12.0346, -11.90528, -11.7758, -11.64615, -11.51633, -11.38634, 
    -11.25619, -11.12587, -10.99538, -10.86472, -10.7339, -10.60291, 
    -10.47176, -10.34044, -10.20896, -10.07731, -9.945492, -9.813514, 
    -9.681371, -9.549064, -9.416594, -9.28396, -9.151164, -9.018206, 
    -8.885084, -8.751801, -8.618357, -8.484752, -8.350986, -8.217059, 
    -8.082973, -7.948726, -7.81432, -7.679756, -7.545033, -7.410152, 
    -7.275113, -7.139917, -7.004565, -6.869056, -6.733391, -6.59757, 
    -6.461595, -6.325465, -6.189181, -6.052743, -5.916152, -5.779408, 
    -5.642512, -5.505465, -5.368266, -5.230916, -5.093416, -4.955767, 
    -4.817968, -4.680021, -4.541926, -4.403683, -4.265293, -4.126757, 
    -3.988075, -3.849247, -3.710275, -3.571159, -3.431899, -3.292496, 
    -3.152951, -3.013264, -2.873436, -2.733467, -2.593359, -2.453111, 
    -2.312725, -2.1722, -2.031539, -1.890741, -1.749806, -1.608737, 
    -1.467533, -1.326195, -1.184723, -1.043119, -0.9013833, -0.7595164, 
    -0.6175189, -0.4753918, -0.3331356, -0.1907512, -0.04823933, 0.09439934, 
    0.237164, 0.380054, 0.5230684, 0.6662065, 0.8094677, 0.9528509, 1.096356, 
    1.239981, 1.383726, 1.52759, 1.671572, 1.815671, 1.959887, 2.104219, 
    2.248665, 2.393226, 2.537899, 2.682685, 2.827582, 2.97259, 3.117708, 
    3.262934, 3.408268, 3.55371, 3.699257, 3.84491, 3.990667, 4.136528, 
    4.28249, 4.428555, 4.57472, 4.720985, 4.867349, 5.013811, 5.160369, 
    5.307024, 5.453773, 5.600616, 5.747553, 5.894582, 6.041701, 6.188911, 
    6.33621, 6.483597, 6.631071, 6.778631, 6.926277, 7.074006, 7.221819, 
    7.369713, 7.517689, 7.665745, 7.813879, 7.962091, 8.110381, 8.258746, 
    8.407187, 8.5557, 8.704287, 8.852944, 9.001673, 9.150471, 9.299336, 
    9.44827, 9.59727, 9.746334, 9.895463, 10.04465, 10.19391, 10.34322, 
    10.4926, 10.64203, 10.79152, 10.94106, 11.09066, 11.24032, 11.39003, 
    11.53979, 11.6896, 11.83946, 11.98936, 12.13932, 12.28932, 12.43937, 
    12.58946, 12.73959, 12.88976, 13.03998, 13.19023, 13.34052, 13.49085, 
    13.64121, 13.79161, 13.94204, 14.09251, 14.243, 14.39352, 14.54408, 
    14.69466, 14.84526, 14.99589, 15.14655, 15.29723, 15.44792, 15.59864, 
    15.74938, 15.90014, 16.05091, 16.2017, 16.3525, 16.50332, 16.65415, 
    16.80499, 16.95583, 17.10669, 17.25755, 17.40842, 17.5593, 17.71017, 
    17.86105, 18.01193, 18.16282, 18.31369, 18.46457, 18.61544, 18.76631, 
    18.91718, 19.06803, 19.21888, 19.36971, 19.52054, 19.67135, 19.82215, 
    19.97294, 20.12371, 20.27446, 20.4252, 20.57591, 20.72661, 20.87729, 
    21.02794, 21.17856, 21.32916, 21.47974, 21.63029, 21.78081, 21.9313, 
    22.08176, 22.23218, 22.38257, 22.53293, 22.68325, 22.83354, 22.98379, 
    23.134, 23.28416, 23.43429, 23.58437, 23.73441, 23.8844, 24.03435, 
    24.18425, 24.3341, 24.48391, 24.63366, 24.78336, 24.933, 25.0826, 
    25.23213, 25.38161, 25.53104, 25.6804, 25.82971, 25.97895, 26.12813, 
    26.27725, 26.4263, 26.57529, 26.72422, 26.87307, 27.02186, 27.17058, 
    27.31922, 27.4678, 27.6163, 27.76473, 27.91308, 28.06136, 28.20956, 
    28.35768, 28.50572, 28.65369, 28.80157, 28.94937, 29.09708, 29.24472, 
    29.39226, 29.53972, 29.6871, 29.83438, 29.98158, 30.12868, 30.2757, 
    30.42262, 30.56945, 30.71618, 30.86282, 31.00936, 31.15581, 31.30216, 
    31.44841, 31.59456, 31.74061, 31.88655, 32.0324, 32.17814, 32.32377, 
    32.4693, 32.61473, 32.76004, 32.90525, 33.05035, 33.19535, 33.34023, 
    33.48499, 33.62965, 33.77419, 33.91862, 34.06293, 34.20713, 34.35121, 
    34.49517, 34.63902, 34.78275, 34.92635, 35.06984, 35.2132, 35.35645, 
    35.49956, 35.64256, 35.78543, 35.92817, 36.07079, 36.21328, 36.35565, 
    36.49788, 36.63999, 36.78197, 36.92381, 37.06553, 37.20711, 37.34856, 
    37.48988, 37.63106, 37.77211, 37.91302, 38.0538, 38.19444, 38.33494, 
    38.4753, 38.61553, 38.75562, 38.89557, 39.03537, 39.17503, 39.31456, 
    39.45394, 39.59317, 39.73227, 39.87122, 40.01002, 40.14868, 40.28719, 
    40.42556, 40.56378, 40.70185, 40.83978, 40.97755, 41.11518, 41.25265, 
    41.38998, 41.52715, 41.66418, 41.80105, 41.93777, 42.07434, 42.21075, 
    42.34701, 42.48312, 42.61906, 42.75486, 42.8905,
  -18.82762, -18.70744, -18.58708, -18.46655, -18.34585, -18.22497, 
    -18.10392, -17.9827, -17.8613, -17.73973, -17.61799, -17.49607, 
    -17.37398, -17.25171, -17.12927, -17.00666, -16.88387, -16.76092, 
    -16.63778, -16.51447, -16.39099, -16.26734, -16.14351, -16.01951, 
    -15.89534, -15.77099, -15.64647, -15.52178, -15.39691, -15.27187, 
    -15.14665, -15.02127, -14.89571, -14.76998, -14.64407, -14.518, 
    -14.39175, -14.26533, -14.13873, -14.01197, -13.88503, -13.75792, 
    -13.63064, -13.50319, -13.37556, -13.24777, -13.1198, -12.99166, 
    -12.86336, -12.73488, -12.60623, -12.47741, -12.34842, -12.21926, 
    -12.08993, -11.96043, -11.83077, -11.70093, -11.57093, -11.44075, 
    -11.31041, -11.1799, -11.04922, -10.91838, -10.78737, -10.65619, 
    -10.52484, -10.39333, -10.26165, -10.1298, -9.997794, -9.865618, 
    -9.733277, -9.600772, -9.468102, -9.335268, -9.20227, -9.069109, 
    -8.935784, -8.802298, -8.668648, -8.534837, -8.400863, -8.266728, 
    -8.132433, -7.997977, -7.863361, -7.728585, -7.59365, -7.458556, 
    -7.323303, -7.187892, -7.052324, -6.916598, -6.780716, -6.644677, 
    -6.508482, -6.372131, -6.235626, -6.098966, -5.962152, -5.825185, 
    -5.688064, -5.550791, -5.413365, -5.275788, -5.138061, -5.000182, 
    -4.862153, -4.723975, -4.585648, -4.447173, -4.308549, -4.169778, 
    -4.030861, -3.891798, -3.752589, -3.613235, -3.473736, -3.334094, 
    -3.194308, -3.05438, -2.91431, -2.774098, -2.633746, -2.493254, 
    -2.352622, -2.211852, -2.070943, -1.929897, -1.788714, -1.647395, 
    -1.50594, -1.364351, -1.222627, -1.08077, -0.9387807, -0.7966593, 
    -0.6544065, -0.5120233, -0.3695103, -0.2268682, -0.08409782, 0.05880012, 
    0.2018249, 0.3449756, 0.4882517, 0.6316522, 0.7751765, 0.9188237, 
    1.062593, 1.206484, 1.350495, 1.494626, 1.638875, 1.783243, 1.927728, 
    2.07233, 2.217047, 2.361879, 2.506824, 2.651883, 2.797054, 2.942336, 
    3.087729, 3.23323, 3.378841, 3.524559, 3.670384, 3.816315, 3.962352, 
    4.108492, 4.254735, 4.401081, 4.547528, 4.694075, 4.840722, 4.987467, 
    5.13431, 5.281249, 5.428284, 5.575413, 5.722637, 5.869952, 6.01736, 
    6.164858, 6.312446, 6.460123, 6.607887, 6.755738, 6.903675, 7.051696, 
    7.199801, 7.347989, 7.496258, 7.644608, 7.793036, 7.941544, 8.090129, 
    8.238791, 8.387527, 8.536338, 8.685222, 8.834178, 8.983205, 9.132301, 
    9.281466, 9.4307, 9.58, 9.729365, 9.878796, 10.02829, 10.17784, 10.32746, 
    10.47714, 10.62687, 10.77667, 10.92652, 11.07642, 11.22638, 11.37639, 
    11.52646, 11.67657, 11.82674, 11.97695, 12.12722, 12.27752, 12.42788, 
    12.57828, 12.72872, 12.8792, 13.02972, 13.18028, 13.33088, 13.48152, 
    13.63219, 13.7829, 13.93364, 14.08442, 14.23522, 14.38605, 14.53692, 
    14.68781, 14.83873, 14.98967, 15.14063, 15.29162, 15.44263, 15.59367, 
    15.74472, 15.89578, 16.04687, 16.19797, 16.34909, 16.50021, 16.65136, 
    16.80251, 16.95367, 17.10484, 17.25601, 17.40719, 17.55838, 17.70957, 
    17.86076, 18.01196, 18.16315, 18.31434, 18.46553, 18.61672, 18.7679, 
    18.91908, 19.07025, 19.22141, 19.37255, 19.52369, 19.67482, 19.82593, 
    19.97703, 20.12811, 20.27918, 20.43023, 20.58125, 20.73226, 20.88325, 
    21.03421, 21.18515, 21.33606, 21.48695, 21.63781, 21.78864, 21.93944, 
    22.09021, 22.24094, 22.39164, 22.54231, 22.69294, 22.84354, 22.99409, 
    23.14461, 23.29508, 23.44552, 23.59591, 23.74625, 23.89655, 24.04681, 
    24.19702, 24.34717, 24.49728, 24.64734, 24.79734, 24.94729, 25.09719, 
    25.24703, 25.39682, 25.54654, 25.69621, 25.84582, 25.99536, 26.14485, 
    26.29427, 26.44362, 26.59291, 26.74213, 26.89129, 27.04037, 27.18939, 
    27.33834, 27.48721, 27.63601, 27.78473, 27.93338, 28.08195, 28.23045, 
    28.37886, 28.5272, 28.67546, 28.82363, 28.97172, 29.11973, 29.26765, 
    29.41549, 29.56324, 29.71091, 29.85848, 30.00596, 30.15336, 30.30066, 
    30.44787, 30.59498, 30.742, 30.88893, 31.03575, 31.18248, 31.32911, 
    31.47565, 31.62208, 31.76841, 31.91463, 32.06076, 32.20678, 32.35269, 
    32.4985, 32.6442, 32.78979, 32.93528, 33.08065, 33.22592, 33.37107, 
    33.51611, 33.66104, 33.80585, 33.95055, 34.09513, 34.2396, 34.38395, 
    34.52818, 34.67229, 34.81628, 34.96016, 35.10391, 35.24754, 35.39104, 
    35.53442, 35.67768, 35.82081, 35.96381, 36.10669, 36.24944, 36.39206, 
    36.53455, 36.67692, 36.81915, 36.96125, 37.10322, 37.24506, 37.38676, 
    37.52832, 37.66976, 37.81105, 37.95222, 38.09324, 38.23413, 38.37488, 
    38.51549, 38.65596, 38.79629, 38.93648, 39.07652, 39.21643, 39.35619, 
    39.49581, 39.63529, 39.77462, 39.91381, 40.05285, 40.19174, 40.33049, 
    40.46909, 40.60754, 40.74584, 40.884, 41.022, 41.15986, 41.29756, 
    41.43512, 41.57251, 41.70977, 41.84686, 41.9838, 42.12059, 42.25723, 
    42.39371, 42.53004, 42.66621, 42.80222, 42.93808,
  -18.89171, -18.77139, -18.6509, -18.53023, -18.40939, -18.28837, -18.16718, 
    -18.04582, -17.92428, -17.80256, -17.68067, -17.55861, -17.43637, 
    -17.31396, -17.19137, -17.06861, -16.94567, -16.82257, -16.69928, 
    -16.57582, -16.45219, -16.32838, -16.2044, -16.08024, -15.95591, 
    -15.83141, -15.70673, -15.58188, -15.45685, -15.33165, -15.20627, 
    -15.08073, -14.95501, -14.82911, -14.70304, -14.5768, -14.45038, 
    -14.3238, -14.19703, -14.0701, -13.94299, -13.81571, -13.68826, 
    -13.56063, -13.43284, -13.30487, -13.17673, -13.04841, -12.91993, 
    -12.79127, -12.66244, -12.53345, -12.40428, -12.27494, -12.14542, 
    -12.01574, -11.88589, -11.75587, -11.62568, -11.49532, -11.36479, 
    -11.23409, -11.10323, -10.97219, -10.84099, -10.70962, -10.57808, 
    -10.44637, -10.3145, -10.18246, -10.05025, -9.917878, -9.785339, 
    -9.652635, -9.519764, -9.386729, -9.25353, -9.120166, -8.986638, 
    -8.852946, -8.719091, -8.585073, -8.450892, -8.31655, -8.182046, 
    -8.047379, -7.912553, -7.777565, -7.642417, -7.50711, -7.371643, 
    -7.236016, -7.100232, -6.964289, -6.828188, -6.69193, -6.555515, 
    -6.418944, -6.282218, -6.145335, -6.008297, -5.871106, -5.73376, 
    -5.596261, -5.458608, -5.320804, -5.182847, -5.044738, -4.906479, 
    -4.76807, -4.62951, -4.490802, -4.351945, -4.212939, -4.073786, 
    -3.934486, -3.795039, -3.655447, -3.515709, -3.375827, -3.2358, -3.09563, 
    -2.955318, -2.814863, -2.674266, -2.533529, -2.392651, -2.251633, 
    -2.110477, -1.969182, -1.82775, -1.686181, -1.544475, -1.402634, 
    -1.260658, -1.118547, -0.9763033, -0.8339267, -0.691418, -0.5487779, 
    -0.4060073, -0.2631069, -0.1200773, 0.02308058, 0.1663661, 0.3097784, 
    0.4533168, 0.5969805, 0.7407686, 0.8846804, 1.028715, 1.172872, 1.31715, 
    1.461549, 1.606067, 1.750704, 1.895459, 2.040331, 2.18532, 2.330424, 
    2.475642, 2.620975, 2.76642, 2.911977, 3.057645, 3.203424, 3.349311, 
    3.495307, 3.641411, 3.787621, 3.933937, 4.080358, 4.226882, 4.37351, 
    4.520239, 4.66707, 4.814001, 4.96103, 5.108158, 5.255383, 5.402704, 
    5.550121, 5.697632, 5.845236, 5.992932, 6.14072, 6.288598, 6.436565, 
    6.58462, 6.732763, 6.880992, 7.029306, 7.177705, 7.326186, 7.47475, 
    7.623395, 7.77212, 7.920923, 8.069804, 8.218763, 8.367797, 8.516906, 
    8.666088, 8.815344, 8.96467, 9.114067, 9.263533, 9.413067, 9.562669, 
    9.712336, 9.862068, 10.01186, 10.16172, 10.31164, 10.46162, 10.61166, 
    10.76176, 10.91192, 11.06213, 11.21239, 11.36271, 11.51308, 11.6635, 
    11.81398, 11.9645, 12.11507, 12.26569, 12.41635, 12.56705, 12.7178, 
    12.86859, 13.01943, 13.1703, 13.32121, 13.47216, 13.62314, 13.77416, 
    13.92521, 14.0763, 14.22741, 14.37856, 14.52973, 14.68094, 14.83217, 
    14.98342, 15.1347, 15.286, 15.43733, 15.58867, 15.74003, 15.89141, 
    16.04281, 16.19423, 16.34566, 16.4971, 16.64855, 16.80002, 16.95149, 
    17.10298, 17.25447, 17.40596, 17.55746, 17.70897, 17.86048, 18.01198, 
    18.16349, 18.315, 18.4665, 18.618, 18.7695, 18.92099, 19.07247, 19.22394, 
    19.37541, 19.52686, 19.6783, 19.82973, 19.98114, 20.13253, 20.28391, 
    20.43527, 20.58661, 20.73793, 20.88923, 21.04051, 21.19176, 21.34298, 
    21.49418, 21.64535, 21.7965, 21.94761, 22.09869, 22.24973, 22.40075, 
    22.55172, 22.70267, 22.85357, 23.00443, 23.15526, 23.30605, 23.45679, 
    23.60749, 23.75814, 23.90875, 24.05931, 24.20983, 24.36029, 24.51071, 
    24.66107, 24.81138, 24.96164, 25.11184, 25.26199, 25.41208, 25.56211, 
    25.71208, 25.86199, 26.01184, 26.16162, 26.31134, 26.461, 26.61059, 
    26.76011, 26.90957, 27.05896, 27.20827, 27.35752, 27.50669, 27.65578, 
    27.80481, 27.95375, 28.10262, 28.25141, 28.40012, 28.54876, 28.69731, 
    28.84578, 28.99416, 29.14246, 29.29068, 29.4388, 29.58685, 29.7348, 
    29.88266, 30.03044, 30.17812, 30.32571, 30.4732, 30.62061, 30.76791, 
    30.91512, 31.06223, 31.20925, 31.35616, 31.50298, 31.64969, 31.7963, 
    31.94281, 32.08921, 32.23552, 32.38171, 32.52779, 32.67377, 32.81964, 
    32.9654, 33.11106, 33.2566, 33.40202, 33.54734, 33.69254, 33.83762, 
    33.98259, 34.12745, 34.27218, 34.4168, 34.5613, 34.70568, 34.84994, 
    34.99408, 35.13809, 35.28199, 35.42575, 35.5694, 35.71292, 35.85631, 
    35.99957, 36.14271, 36.28572, 36.4286, 36.57135, 36.71397, 36.85646, 
    36.99881, 37.14104, 37.28312, 37.42508, 37.5669, 37.70858, 37.85013, 
    37.99154, 38.13282, 38.27395, 38.41494, 38.5558, 38.69651, 38.83709, 
    38.97752, 39.11781, 39.25796, 39.39796, 39.53782, 39.67754, 39.81711, 
    39.95653, 40.09581, 40.23494, 40.37392, 40.51275, 40.65144, 40.78997, 
    40.92836, 41.0666, 41.20468, 41.34261, 41.48039, 41.61802, 41.7555, 
    41.89282, 42.02998, 42.167, 42.30386, 42.44056, 42.57711, 42.71349, 
    42.84973, 42.9858,
  -18.95597, -18.83551, -18.71488, -18.59407, -18.47309, -18.35193, -18.2306, 
    -18.10909, -17.98741, -17.86555, -17.74352, -17.62131, -17.49893, 
    -17.37637, -17.25363, -17.13072, -17.00764, -16.88438, -16.76094, 
    -16.63733, -16.51355, -16.38959, -16.26545, -16.14114, -16.01665, 
    -15.89199, -15.76715, -15.64214, -15.51696, -15.39159, -15.26606, 
    -15.14035, -15.01446, -14.8884, -14.76217, -14.63576, -14.50918, 
    -14.38243, -14.2555, -14.12839, -14.00111, -13.87366, -13.74604, 
    -13.61824, -13.49027, -13.36213, -13.23381, -13.10532, -12.97666, 
    -12.84783, -12.71882, -12.58964, -12.46029, -12.33077, -12.20108, 
    -12.07121, -11.94118, -11.81097, -11.6806, -11.55005, -11.41933, 
    -11.28845, -11.15739, -11.02616, -10.89477, -10.76321, -10.63147, 
    -10.49957, -10.36751, -10.23527, -10.10287, -9.970294, -9.837557, 
    -9.704653, -9.571582, -9.438346, -9.304944, -9.171377, -9.037645, 
    -8.903749, -8.769688, -8.635464, -8.501076, -8.366525, -8.231811, 
    -8.096934, -7.961896, -7.826696, -7.691336, -7.555814, -7.420132, 
    -7.28429, -7.148289, -7.012128, -6.875809, -6.739332, -6.602697, 
    -6.465905, -6.328956, -6.19185, -6.054589, -5.917172, -5.779601, 
    -5.641875, -5.503995, -5.365963, -5.227777, -5.089438, -4.950948, 
    -4.812306, -4.673514, -4.534572, -4.395481, -4.256239, -4.11685, 
    -3.977313, -3.837628, -3.697797, -3.55782, -3.417696, -3.277429, 
    -3.137016, -2.99646, -2.855761, -2.71492, -2.573936, -2.432812, 
    -2.291547, -2.150142, -2.008599, -1.866916, -1.725096, -1.583139, 
    -1.441045, -1.298815, -1.156451, -1.013952, -0.8713194, -0.7285541, 
    -0.5856566, -0.4426277, -0.2994682, -0.1561787, -0.01276013, 0.1307869, 
    0.2744614, 0.4182629, 0.5621904, 0.7062432, 0.8504204, 0.9947214, 
    1.139145, 1.283691, 1.428358, 1.573146, 1.718053, 1.863078, 2.008222, 
    2.153483, 2.29886, 2.444352, 2.589959, 2.735679, 2.881512, 3.027457, 
    3.173512, 3.319678, 3.465953, 3.612336, 3.758826, 3.905423, 4.052125, 
    4.198932, 4.345842, 4.492855, 4.63997, 4.787185, 4.9345, 5.081914, 
    5.229426, 5.377034, 5.524739, 5.672538, 5.820431, 5.968418, 6.116496, 
    6.264665, 6.412923, 6.561271, 6.709706, 6.858229, 7.006836, 7.155529, 
    7.304306, 7.453165, 7.602106, 7.751127, 7.900228, 8.049407, 8.198664, 
    8.347996, 8.497404, 8.646886, 8.796441, 8.946068, 9.095766, 9.245534, 
    9.39537, 9.545274, 9.695244, 9.84528, 9.995378, 10.14554, 10.29577, 
    10.44605, 10.5964, 10.7468, 10.89726, 11.04778, 11.19835, 11.34898, 
    11.49966, 11.65039, 11.80117, 11.952, 12.10288, 12.2538, 12.40477, 
    12.55579, 12.70685, 12.85795, 13.00909, 13.16028, 13.3115, 13.46276, 
    13.61405, 13.76538, 13.91675, 14.06815, 14.21957, 14.37103, 14.52252, 
    14.67404, 14.82558, 14.97715, 15.12874, 15.28036, 15.432, 15.58365, 
    15.73533, 15.88703, 16.03874, 16.19047, 16.34221, 16.49397, 16.64574, 
    16.79752, 16.94931, 17.10111, 17.25291, 17.40473, 17.55654, 17.70836, 
    17.86018, 18.01201, 18.16383, 18.31565, 18.46747, 18.61929, 18.7711, 
    18.9229, 19.0747, 19.22649, 19.37827, 19.53004, 19.68179, 19.83353, 
    19.98526, 20.13697, 20.28866, 20.44034, 20.59199, 20.74363, 20.89524, 
    21.04683, 21.19839, 21.34993, 21.50144, 21.65293, 21.80438, 21.9558, 
    22.1072, 22.25856, 22.40988, 22.56117, 22.71243, 22.86364, 23.01482, 
    23.16595, 23.31705, 23.4681, 23.61911, 23.77007, 23.92099, 24.07186, 
    24.22269, 24.37346, 24.52418, 24.67485, 24.82547, 24.97603, 25.12654, 
    25.27699, 25.42739, 25.57772, 25.728, 25.87822, 26.02837, 26.17846, 
    26.32848, 26.47844, 26.62834, 26.77816, 26.92792, 27.0776, 27.22722, 
    27.37676, 27.52624, 27.67563, 27.82495, 27.9742, 28.12336, 28.27245, 
    28.42146, 28.57039, 28.71923, 28.868, 29.01668, 29.16527, 29.31378, 
    29.4622, 29.61053, 29.75878, 29.90693, 30.055, 30.20297, 30.35085, 
    30.49863, 30.64632, 30.79391, 30.94141, 31.08881, 31.23611, 31.38331, 
    31.53041, 31.6774, 31.8243, 31.97109, 32.11777, 32.26435, 32.41083, 
    32.55719, 32.70345, 32.8496, 32.99564, 33.14156, 33.28738, 33.43308, 
    33.57867, 33.72414, 33.8695, 34.01474, 34.15987, 34.30488, 34.44976, 
    34.59454, 34.73918, 34.88371, 35.02811, 35.17239, 35.31655, 35.46059, 
    35.60449, 35.74828, 35.89193, 36.03545, 36.17885, 36.32212, 36.46526, 
    36.60827, 36.75114, 36.89389, 37.0365, 37.17898, 37.32132, 37.46353, 
    37.6056, 37.74754, 37.88934, 38.031, 38.17252, 38.3139, 38.45515, 
    38.59625, 38.73721, 38.87803, 39.0187, 39.15924, 39.29963, 39.43987, 
    39.57997, 39.71992, 39.85973, 39.9994, 40.13891, 40.27827, 40.41749, 
    40.55656, 40.69548, 40.83425, 40.97287, 41.11133, 41.24965, 41.38781, 
    41.52582, 41.66367, 41.80137, 41.93892, 42.07631, 42.21355, 42.35063, 
    42.48755, 42.62432, 42.76093, 42.89738, 43.03368,
  -19.02039, -18.89979, -18.77902, -18.65808, -18.53696, -18.41566, 
    -18.29419, -18.17253, -18.05071, -17.92871, -17.80653, -17.68418, 
    -17.56165, -17.43894, -17.31606, -17.193, -17.06977, -16.94636, 
    -16.82277, -16.69901, -16.57507, -16.45095, -16.32666, -16.20219, 
    -16.07755, -15.95273, -15.82774, -15.70257, -15.57722, -15.4517, 
    -15.32601, -15.20013, -15.07409, -14.94786, -14.82146, -14.69489, 
    -14.56814, -14.44122, -14.31412, -14.18685, -14.0594, -13.93178, 
    -13.80398, -13.67601, -13.54787, -13.41955, -13.29106, -13.16239, 
    -13.03356, -12.90454, -12.77536, -12.646, -12.51647, -12.38677, 
    -12.25689, -12.12684, -11.99662, -11.86623, -11.73567, -11.60494, 
    -11.47403, -11.34296, -11.21171, -11.08029, -10.94871, -10.81695, 
    -10.68503, -10.55293, -10.42067, -10.28824, -10.15564, -10.02287, 
    -9.889931, -9.756827, -9.623556, -9.490119, -9.356514, -9.222744, 
    -9.088808, -8.954706, -8.820439, -8.686007, -8.551412, -8.416652, 
    -8.281729, -8.146642, -8.011392, -7.87598, -7.740406, -7.60467, 
    -7.468772, -7.332715, -7.196496, -7.060118, -6.92358, -6.786883, 
    -6.650027, -6.513013, -6.375842, -6.238513, -6.101027, -5.963386, 
    -5.825588, -5.687635, -5.549528, -5.411266, -5.27285, -5.134281, 
    -4.99556, -4.856686, -4.717661, -4.578485, -4.439157, -4.299681, 
    -4.160055, -4.020279, -3.880356, -3.740286, -3.600068, -3.459704, 
    -3.319194, -3.178538, -3.037739, -2.896795, -2.755708, -2.614478, 
    -2.473107, -2.331594, -2.18994, -2.048146, -1.906213, -1.764141, 
    -1.621932, -1.479585, -1.337101, -1.194482, -1.051727, -0.9088383, 
    -0.7658157, -0.62266, -0.4793722, -0.3359529, -0.1924029, -0.04872286, 
    0.09508632, 0.2390239, 0.3830892, 0.5272812, 0.6715994, 0.8160428, 
    0.9606107, 1.105302, 1.250116, 1.395053, 1.54011, 1.685288, 1.830586, 
    1.976002, 2.121535, 2.267186, 2.412953, 2.558835, 2.704831, 2.850941, 
    2.997163, 3.143497, 3.289941, 3.436496, 3.583159, 3.72993, 3.876809, 
    4.023793, 4.170883, 4.318077, 4.465374, 4.612773, 4.760274, 4.907876, 
    5.055577, 5.203376, 5.351273, 5.499266, 5.647355, 5.795538, 5.943815, 
    6.092185, 6.240645, 6.389197, 6.537838, 6.686566, 6.835383, 6.984286, 
    7.133274, 7.282347, 7.431502, 7.58074, 7.730059, 7.879457, 8.028935, 
    8.178491, 8.328123, 8.477832, 8.627614, 8.777471, 8.927399, 9.077399, 
    9.227469, 9.377608, 9.527816, 9.678089, 9.828429, 9.978834, 10.1293, 
    10.27983, 10.43042, 10.58107, 10.73179, 10.88255, 11.03338, 11.18426, 
    11.33519, 11.48618, 11.63722, 11.78831, 11.93945, 12.09064, 12.24188, 
    12.39316, 12.54449, 12.69586, 12.84727, 12.99872, 13.15022, 13.30175, 
    13.45333, 13.60493, 13.75658, 13.90825, 14.05997, 14.21171, 14.36348, 
    14.51528, 14.66711, 14.81897, 14.97086, 15.12276, 15.27469, 15.42665, 
    15.57862, 15.73061, 15.88263, 16.03465, 16.1867, 16.33876, 16.49083, 
    16.64292, 16.79502, 16.94712, 17.09924, 17.25136, 17.40348, 17.55562, 
    17.70775, 17.85989, 18.01203, 18.16417, 18.31631, 18.46845, 18.62058, 
    18.77271, 18.92483, 19.07694, 19.22905, 19.38114, 19.53322, 19.6853, 
    19.83735, 19.98939, 20.14142, 20.29343, 20.44542, 20.59739, 20.74934, 
    20.90127, 21.05317, 21.20505, 21.3569, 21.50873, 21.66053, 21.8123, 
    21.96404, 22.11574, 22.26741, 22.41905, 22.57065, 22.72222, 22.87375, 
    23.02524, 23.17668, 23.32809, 23.47945, 23.63078, 23.78205, 23.93328, 
    24.08446, 24.23559, 24.38667, 24.53771, 24.68869, 24.83961, 24.99048, 
    25.1413, 25.29206, 25.44276, 25.5934, 25.74398, 25.8945, 26.04496, 
    26.19536, 26.34569, 26.49595, 26.64615, 26.79627, 26.94633, 27.09632, 
    27.24624, 27.39608, 27.54585, 27.69555, 27.84517, 27.99471, 28.14418, 
    28.29357, 28.44287, 28.5921, 28.74124, 28.8903, 29.03927, 29.18816, 
    29.33697, 29.48568, 29.63431, 29.78284, 29.93129, 30.07965, 30.22791, 
    30.37608, 30.52415, 30.67213, 30.82001, 30.96779, 31.11548, 31.26307, 
    31.41055, 31.55793, 31.70521, 31.85239, 31.99946, 32.14643, 32.29329, 
    32.44005, 32.58669, 32.73323, 32.87966, 33.02597, 33.17218, 33.31827, 
    33.46425, 33.61011, 33.75586, 33.90149, 34.04701, 34.19241, 34.33768, 
    34.48285, 34.62788, 34.7728, 34.91759, 35.06227, 35.20681, 35.35124, 
    35.49554, 35.63971, 35.78375, 35.92767, 36.07146, 36.21512, 36.35865, 
    36.50205, 36.64531, 36.78845, 36.93145, 37.07432, 37.21705, 37.35965, 
    37.50211, 37.64444, 37.78662, 37.92867, 38.07058, 38.21236, 38.35399, 
    38.49548, 38.63683, 38.77803, 38.9191, 39.06002, 39.2008, 39.34143, 
    39.48192, 39.62226, 39.76245, 39.9025, 40.0424, 40.18215, 40.32175, 
    40.46121, 40.60051, 40.73966, 40.87866, 41.01751, 41.15621, 41.29475, 
    41.43315, 41.57138, 41.70947, 41.8474, 41.98517, 42.12279, 42.26025, 
    42.39755, 42.5347, 42.67168, 42.80852, 42.94519, 43.0817,
  -19.08497, -18.96424, -18.84333, -18.72225, -18.60098, -18.47955, 
    -18.35793, -18.23614, -18.11417, -17.99203, -17.86971, -17.74721, 
    -17.62453, -17.50168, -17.37865, -17.25544, -17.13206, -17.0085, 
    -16.88476, -16.76084, -16.63675, -16.51248, -16.38804, -16.26342, 
    -16.13862, -16.01364, -15.88849, -15.76316, -15.63766, -15.51198, 
    -15.38612, -15.26008, -15.13387, -15.00748, -14.88092, -14.75418, 
    -14.62727, -14.50018, -14.37291, -14.24547, -14.11785, -13.99006, 
    -13.86209, -13.73395, -13.60563, -13.47714, -13.34847, -13.21963, 
    -13.09061, -12.96142, -12.83206, -12.70252, -12.57281, -12.44292, 
    -12.31287, -12.18264, -12.05223, -11.92165, -11.79091, -11.65999, 
    -11.52889, -11.39763, -11.26619, -11.13459, -11.00281, -10.87086, 
    -10.73874, -10.60645, -10.47399, -10.34136, -10.20857, -10.0756, 
    -9.942464, -9.80916, -9.675688, -9.542048, -9.408241, -9.274267, 
    -9.140127, -9.005819, -8.871346, -8.736708, -8.601904, -8.466934, 
    -8.3318, -8.196503, -8.061042, -7.925416, -7.789629, -7.653678, 
    -7.517565, -7.38129, -7.244855, -7.108258, -6.971501, -6.834584, 
    -6.697507, -6.560271, -6.422877, -6.285324, -6.147614, -6.009747, 
    -5.871722, -5.733542, -5.595206, -5.456715, -5.318069, -5.179269, 
    -5.040316, -4.901209, -4.76195, -4.622539, -4.482977, -4.343264, -4.2034, 
    -4.063387, -3.923224, -3.782914, -3.642455, -3.501849, -3.361096, 
    -3.220198, -3.079154, -2.937965, -2.796632, -2.655155, -2.513535, 
    -2.371774, -2.22987, -2.087826, -1.945642, -1.803318, -1.660855, 
    -1.518255, -1.375516, -1.232641, -1.08963, -0.9464844, -0.8032037, 
    -0.6597892, -0.5162417, -0.3725619, -0.2287506, -0.08480848, 0.05926363, 
    0.203465, 0.3477947, 0.4922522, 0.6368364, 0.7815468, 0.9263824, 
    1.071342, 1.216426, 1.361632, 1.506961, 1.65241, 1.79798, 1.943669, 
    2.089476, 2.235402, 2.381444, 2.527602, 2.673875, 2.820262, 2.966763, 
    3.113375, 3.2601, 3.406934, 3.553879, 3.700932, 3.848093, 3.995361, 
    4.142735, 4.290213, 4.437795, 4.585481, 4.733268, 4.881157, 5.029146, 
    5.177234, 5.325419, 5.473702, 5.622082, 5.770556, 5.919125, 6.067786, 
    6.21654, 6.365385, 6.514319, 6.663343, 6.812455, 6.961654, 7.110939, 
    7.260308, 7.409761, 7.559297, 7.708914, 7.858612, 8.008389, 8.158245, 
    8.308178, 8.458187, 8.608272, 8.75843, 8.908662, 9.058965, 9.209338, 
    9.359782, 9.510294, 9.660872, 9.811518, 9.962228, 10.113, 10.26384, 
    10.41474, 10.5657, 10.71671, 10.86779, 11.01893, 11.17011, 11.32136, 
    11.47266, 11.62401, 11.77541, 11.92686, 12.07836, 12.22991, 12.3815, 
    12.53314, 12.68482, 12.83655, 12.98832, 13.14012, 13.29197, 13.44386, 
    13.59578, 13.74774, 13.89973, 14.05176, 14.20381, 14.3559, 14.50802, 
    14.66017, 14.81234, 14.96454, 15.11676, 15.26901, 15.42128, 15.57357, 
    15.72588, 15.87821, 16.03055, 16.18292, 16.33529, 16.48768, 16.64009, 
    16.7925, 16.94492, 17.09735, 17.24979, 17.40224, 17.55469, 17.70714, 
    17.8596, 18.01206, 18.16452, 18.31697, 18.46943, 18.62188, 18.77432, 
    18.92676, 19.07919, 19.23161, 19.38402, 19.53642, 19.68881, 19.84119, 
    19.99355, 20.14589, 20.29822, 20.45052, 20.60281, 20.75508, 20.90732, 
    21.05954, 21.21173, 21.3639, 21.51604, 21.66816, 21.82024, 21.97229, 
    22.12432, 22.2763, 22.42826, 22.58017, 22.73205, 22.88389, 23.03569, 
    23.18745, 23.33917, 23.49085, 23.64248, 23.79407, 23.94561, 24.0971, 
    24.24854, 24.39994, 24.55128, 24.70257, 24.85381, 25.00499, 25.15611, 
    25.30718, 25.45819, 25.60914, 25.76003, 25.91085, 26.06162, 26.21232, 
    26.36295, 26.51352, 26.66402, 26.81445, 26.96482, 27.11511, 27.26533, 
    27.41547, 27.56555, 27.71554, 27.86547, 28.01531, 28.16507, 28.31476, 
    28.46436, 28.61389, 28.76333, 28.91268, 29.06195, 29.21114, 29.36024, 
    29.50924, 29.65817, 29.807, 29.95574, 30.10438, 30.25294, 30.4014, 
    30.54976, 30.69803, 30.8462, 30.99427, 31.14224, 31.29012, 31.43789, 
    31.58556, 31.73312, 31.88058, 32.02794, 32.17519, 32.32234, 32.46937, 
    32.6163, 32.76312, 32.90982, 33.05642, 33.2029, 33.34927, 33.49553, 
    33.64167, 33.78769, 33.9336, 34.07938, 34.22506, 34.37061, 34.51604, 
    34.66135, 34.80653, 34.9516, 35.09654, 35.24135, 35.38604, 35.53061, 
    35.67505, 35.81936, 35.96354, 36.10759, 36.25151, 36.3953, 36.53896, 
    36.68248, 36.82588, 36.96914, 37.11226, 37.25525, 37.39811, 37.54082, 
    37.6834, 37.82584, 37.96814, 38.11031, 38.25233, 38.39421, 38.53595, 
    38.67754, 38.819, 38.96031, 39.10147, 39.2425, 39.38337, 39.5241, 
    39.66468, 39.80512, 39.9454, 40.08554, 40.22553, 40.36538, 40.50506, 
    40.6446, 40.78399, 40.92323, 41.06231, 41.20124, 41.34001, 41.47863, 
    41.6171, 41.75541, 41.89357, 42.03157, 42.16941, 42.30709, 42.44462, 
    42.58199, 42.7192, 42.85625, 42.99314, 43.12988,
  -19.14972, -19.02885, -18.9078, -18.78658, -18.66518, -18.5436, -18.42184, 
    -18.29991, -18.1778, -18.05551, -17.93305, -17.8104, -17.68758, 
    -17.56458, -17.4414, -17.31805, -17.19451, -17.0708, -16.94691, 
    -16.82285, -16.6986, -16.57418, -16.44958, -16.3248, -16.19985, 
    -16.07472, -15.94941, -15.82392, -15.69826, -15.57241, -15.44639, 
    -15.3202, -15.19382, -15.06727, -14.94054, -14.81364, -14.68656, 
    -14.5593, -14.43186, -14.30425, -14.17647, -14.0485, -13.92036, 
    -13.79205, -13.66356, -13.53489, -13.40604, -13.27703, -13.14783, 
    -13.01847, -12.88892, -12.7592, -12.62931, -12.49925, -12.369, -12.23859, 
    -12.108, -11.97724, -11.8463, -11.7152, -11.58391, -11.45246, -11.32084, 
    -11.18904, -11.05707, -10.92493, -10.79261, -10.66013, -10.52748, 
    -10.39465, -10.26165, -10.12849, -9.995155, -9.861651, -9.727978, 
    -9.594136, -9.460127, -9.325949, -9.191603, -9.05709, -8.92241, 
    -8.787564, -8.652551, -8.517372, -8.382029, -8.246519, -8.110846, 
    -7.975007, -7.839005, -7.702839, -7.566511, -7.430019, -7.293365, 
    -7.15655, -7.019573, -6.882436, -6.745138, -6.607679, -6.470061, 
    -6.332285, -6.194349, -6.056256, -5.918005, -5.779596, -5.641032, 
    -5.502311, -5.363434, -5.224403, -5.085217, -4.945877, -4.806384, 
    -4.666738, -4.526939, -4.386989, -4.246888, -4.106636, -3.966234, 
    -3.825682, -3.684982, -3.544134, -3.403138, -3.261995, -3.120706, 
    -2.979271, -2.837692, -2.695967, -2.554099, -2.412088, -2.269935, 
    -2.12764, -1.985203, -1.842627, -1.69991, -1.557055, -1.414061, -1.27093, 
    -1.127662, -0.9842584, -0.840719, -0.697045, -0.5532371, -0.4092962, 
    -0.2652228, -0.1210178, 0.02331792, 0.1677837, 0.3123788, 0.4571023, 
    0.6019534, 0.7469314, 0.8920355, 1.037265, 1.182618, 1.328096, 1.473696, 
    1.619417, 1.76526, 1.911223, 2.057305, 2.203506, 2.349824, 2.496259, 
    2.64281, 2.789476, 2.936255, 3.083148, 3.230153, 3.377269, 3.524495, 
    3.671831, 3.819276, 3.966827, 4.114486, 4.262249, 4.410118, 4.558091, 
    4.706166, 4.854342, 5.00262, 5.150997, 5.299473, 5.448047, 5.596718, 
    5.745484, 5.894345, 6.0433, 6.192348, 6.341487, 6.490717, 6.640036, 
    6.789444, 6.93894, 7.088521, 7.238189, 7.38794, 7.537776, 7.687693, 
    7.83769, 7.987769, 8.137925, 8.28816, 8.438472, 8.588859, 8.739321, 
    8.889855, 9.040462, 9.191141, 9.341889, 9.492707, 9.643592, 9.794544, 
    9.945561, 10.09664, 10.24779, 10.39899, 10.55026, 10.70159, 10.85298, 
    11.00442, 11.15592, 11.30747, 11.45908, 11.61074, 11.76246, 11.91422, 
    12.06603, 12.21789, 12.3698, 12.52175, 12.67375, 12.82579, 12.97787, 
    13.12999, 13.28215, 13.43435, 13.58659, 13.73886, 13.89117, 14.04351, 
    14.19589, 14.34829, 14.50073, 14.65319, 14.80568, 14.9582, 15.11074, 
    15.2633, 15.41589, 15.5685, 15.72113, 15.87377, 16.02644, 16.17912, 
    16.33181, 16.48452, 16.63724, 16.78997, 16.94272, 17.09547, 17.24822, 
    17.40099, 17.55376, 17.70653, 17.85931, 18.01208, 18.16486, 18.31763, 
    18.47041, 18.62318, 18.77594, 18.9287, 19.08145, 19.23419, 19.38692, 
    19.53964, 19.69234, 19.84504, 19.99771, 20.15038, 20.30302, 20.45564, 
    20.60825, 20.76083, 20.91339, 21.06593, 21.21844, 21.37093, 21.52339, 
    21.67582, 21.82822, 21.98059, 22.13292, 22.28522, 22.43749, 22.58972, 
    22.74192, 22.89407, 23.04619, 23.19827, 23.3503, 23.50229, 23.65423, 
    23.80613, 23.95799, 24.10979, 24.26155, 24.41325, 24.5649, 24.7165, 
    24.86805, 25.01954, 25.17097, 25.32235, 25.47367, 25.62493, 25.77612, 
    25.92726, 26.07833, 26.22934, 26.38028, 26.53115, 26.68196, 26.8327, 
    26.98337, 27.13396, 27.28448, 27.43493, 27.58531, 27.73561, 27.88583, 
    28.03598, 28.18604, 28.33603, 28.48593, 28.63575, 28.78549, 28.93515, 
    29.08471, 29.2342, 29.38359, 29.53289, 29.68211, 29.83124, 29.98027, 
    30.12921, 30.27806, 30.42681, 30.57546, 30.72402, 30.87248, 31.02084, 
    31.1691, 31.31726, 31.46532, 31.61328, 31.76113, 31.90888, 32.05652, 
    32.20406, 32.35148, 32.4988, 32.64601, 32.79311, 32.94009, 33.08697, 
    33.23373, 33.38038, 33.52691, 33.67333, 33.81963, 33.96581, 34.11187, 
    34.25782, 34.40364, 34.54934, 34.69492, 34.84038, 34.98572, 35.13092, 
    35.27601, 35.42097, 35.5658, 35.7105, 35.85508, 35.99952, 36.14384, 
    36.28802, 36.43208, 36.57599, 36.71978, 36.86343, 37.00695, 37.15033, 
    37.29358, 37.43669, 37.57966, 37.7225, 37.86519, 38.00774, 38.15016, 
    38.29243, 38.43456, 38.57655, 38.7184, 38.8601, 39.00166, 39.14307, 
    39.28433, 39.42545, 39.56643, 39.70725, 39.84793, 39.98845, 40.12883, 
    40.26906, 40.40914, 40.54906, 40.68884, 40.82846, 40.96793, 41.10724, 
    41.24641, 41.38541, 41.52427, 41.66296, 41.8015, 41.93988, 42.07811, 
    42.21618, 42.35409, 42.49184, 42.62943, 42.76686, 42.90414, 43.04125, 
    43.1782,
  -19.21463, -19.09362, -18.97244, -18.85108, -18.72954, -18.60782, 
    -18.48592, -18.36385, -18.24159, -18.11916, -17.99655, -17.87376, 
    -17.7508, -17.62765, -17.50432, -17.38082, -17.25714, -17.13328, 
    -17.00924, -16.88502, -16.76062, -16.63605, -16.51129, -16.38636, 
    -16.26125, -16.13596, -16.01049, -15.88484, -15.75902, -15.63302, 
    -15.50684, -15.38048, -15.25394, -15.12723, -15.00033, -14.87326, 
    -14.74601, -14.61859, -14.49098, -14.3632, -14.23525, -14.10711, 
    -13.9788, -13.85031, -13.72165, -13.5928, -13.46379, -13.33459, 
    -13.20522, -13.07567, -12.94595, -12.81605, -12.68598, -12.55573, 
    -12.42531, -12.29471, -12.16393, -12.03299, -11.90187, -11.77057, 
    -11.6391, -11.50746, -11.37564, -11.24365, -11.11149, -10.97916, 
    -10.84665, -10.71397, -10.58112, -10.4481, -10.31491, -10.18154, 
    -10.04801, -9.914302, -9.780428, -9.646384, -9.512171, -9.377789, 
    -9.243237, -9.108519, -8.973632, -8.838577, -8.703356, -8.567967, 
    -8.432412, -8.296692, -8.160805, -8.024754, -7.888537, -7.752156, 
    -7.615611, -7.478902, -7.34203, -7.204996, -7.067799, -6.93044, -6.79292, 
    -6.655239, -6.517397, -6.379395, -6.241235, -6.102915, -5.964436, 
    -5.825799, -5.687006, -5.548054, -5.408947, -5.269683, -5.130264, 
    -4.990691, -4.850963, -4.711081, -4.571045, -4.430858, -4.290518, 
    -4.150027, -4.009385, -3.868592, -3.72765, -3.586559, -3.445319, 
    -3.303932, -3.162397, -3.020716, -2.878889, -2.736916, -2.594799, 
    -2.452538, -2.310134, -2.167587, -2.024898, -1.882068, -1.739097, 
    -1.595987, -1.452737, -1.30935, -1.165824, -1.022161, -0.8783625, 
    -0.7344283, -0.5903593, -0.4461564, -0.3018204, -0.1573518, -0.01275169, 
    0.1319793, 0.2768404, 0.4218307, 0.5669495, 0.712196, 0.8575693, 
    1.003069, 1.148693, 1.294442, 1.440314, 1.586309, 1.732426, 1.878664, 
    2.025021, 2.171498, 2.318094, 2.464806, 2.611636, 2.75858, 2.90564, 
    3.052814, 3.2001, 3.347498, 3.495007, 3.642627, 3.790355, 3.938192, 
    4.086136, 4.234187, 4.382342, 4.530602, 4.678966, 4.827432, 4.975999, 
    5.124667, 5.273434, 5.422299, 5.571262, 5.720322, 5.869476, 6.018725, 
    6.168068, 6.317502, 6.467029, 6.616644, 6.76635, 6.916143, 7.066023, 
    7.21599, 7.366041, 7.516176, 7.666393, 7.816693, 7.967072, 8.117532, 
    8.268069, 8.418684, 8.569375, 8.72014, 8.87098, 9.021894, 9.172877, 
    9.323932, 9.475056, 9.626248, 9.777508, 9.928833, 10.08022, 10.23168, 
    10.38319, 10.53477, 10.68641, 10.8381, 10.98986, 11.14167, 11.29354, 
    11.44546, 11.59743, 11.74946, 11.90153, 12.05366, 12.20583, 12.35805, 
    12.51032, 12.66263, 12.81499, 12.96738, 13.11982, 13.2723, 13.42482, 
    13.57737, 13.72996, 13.88258, 14.03524, 14.18793, 14.34066, 14.49341, 
    14.64619, 14.799, 14.95183, 15.10469, 15.25758, 15.41048, 15.56341, 
    15.71636, 15.86932, 16.0223, 16.1753, 16.32832, 16.48135, 16.63439, 
    16.78744, 16.9405, 17.09357, 17.24665, 17.39973, 17.55282, 17.70592, 
    17.85901, 18.01211, 18.16521, 18.3183, 18.47139, 18.62448, 18.77757, 
    18.93064, 19.08371, 19.23677, 19.38982, 19.54286, 19.69589, 19.8489, 
    20.0019, 20.15488, 20.30784, 20.46078, 20.61371, 20.76661, 20.91949, 
    21.07235, 21.22518, 21.37798, 21.53076, 21.6835, 21.83622, 21.98891, 
    22.14156, 22.29418, 22.44676, 22.59931, 22.75182, 22.90429, 23.05673, 
    23.20912, 23.36147, 23.51377, 23.66603, 23.81824, 23.97041, 24.12253, 
    24.2746, 24.42661, 24.57858, 24.73049, 24.88235, 25.03415, 25.1859, 
    25.33758, 25.48921, 25.64078, 25.79229, 25.94373, 26.09511, 26.24642, 
    26.39767, 26.54885, 26.69997, 26.85101, 27.00198, 27.15289, 27.30371, 
    27.45447, 27.60515, 27.75575, 27.90627, 28.05672, 28.20709, 28.35737, 
    28.50758, 28.6577, 28.80774, 28.95769, 29.10756, 29.25734, 29.40703, 
    29.55663, 29.70614, 29.85556, 30.00489, 30.15412, 30.30326, 30.45231, 
    30.60126, 30.7501, 30.89886, 31.04751, 31.19606, 31.34451, 31.49286, 
    31.6411, 31.78924, 31.93727, 32.0852, 32.23302, 32.38073, 32.52834, 
    32.67583, 32.82321, 32.97047, 33.11763, 33.26467, 33.4116, 33.55841, 
    33.7051, 33.85168, 33.99814, 34.14448, 34.2907, 34.43679, 34.58277, 
    34.72862, 34.87435, 35.01995, 35.16544, 35.31079, 35.45601, 35.60111, 
    35.74608, 35.89092, 36.03563, 36.18021, 36.32466, 36.46898, 36.61316, 
    36.75721, 36.90112, 37.0449, 37.18854, 37.33204, 37.47541, 37.61863, 
    37.76172, 37.90467, 38.04748, 38.19014, 38.33267, 38.47505, 38.61729, 
    38.75938, 38.90133, 39.04314, 39.1848, 39.32631, 39.46767, 39.60889, 
    39.74995, 39.89087, 40.03164, 40.17226, 40.31273, 40.45304, 40.59321, 
    40.73322, 40.87308, 41.01278, 41.15233, 41.29172, 41.43096, 41.57005, 
    41.70897, 41.84774, 41.98635, 42.12481, 42.2631, 42.40124, 42.53921, 
    42.67703, 42.81469, 42.95218, 43.08951, 43.22668,
  -19.27971, -19.15857, -19.03724, -18.91574, -18.79407, -18.67221, 
    -18.55017, -18.42795, -18.30556, -18.18298, -18.06023, -17.93729, 
    -17.81418, -17.69089, -17.56741, -17.44376, -17.31993, -17.19592, 
    -17.07173, -16.94736, -16.82281, -16.69808, -16.57317, -16.44808, 
    -16.32281, -16.19737, -16.07174, -15.94594, -15.81995, -15.69379, 
    -15.56745, -15.44093, -15.31423, -15.18735, -15.06029, -14.93305, 
    -14.80564, -14.67804, -14.55027, -14.42232, -14.29419, -14.16589, 
    -14.0374, -13.90874, -13.7799, -13.65089, -13.52169, -13.39232, 
    -13.26277, -13.13305, -13.00315, -12.87307, -12.74281, -12.61238, 
    -12.48177, -12.35099, -12.22003, -12.0889, -11.95759, -11.82611, 
    -11.69445, -11.56262, -11.43061, -11.29843, -11.16607, -11.03355, 
    -10.90085, -10.76797, -10.63493, -10.50171, -10.36832, -10.23475, 
    -10.10102, -9.967114, -9.833038, -9.698792, -9.564374, -9.429788, 
    -9.295032, -9.160106, -9.025012, -8.889749, -8.754318, -8.61872, 
    -8.482954, -8.347021, -8.210921, -8.074656, -7.938224, -7.801627, 
    -7.664865, -7.527939, -7.390849, -7.253595, -7.116178, -6.978597, 
    -6.840855, -6.70295, -6.564885, -6.426658, -6.288271, -6.149724, 
    -6.011017, -5.872152, -5.733128, -5.593946, -5.454607, -5.315111, 
    -5.175459, -5.035651, -4.895688, -4.755569, -4.615297, -4.474872, 
    -4.334293, -4.193562, -4.052679, -3.911645, -3.77046, -3.629125, 
    -3.487641, -3.346009, -3.204228, -3.062299, -2.920224, -2.778003, 
    -2.635636, -2.493125, -2.350469, -2.20767, -2.064728, -1.921643, 
    -1.778418, -1.635052, -1.491545, -1.3479, -1.204116, -1.060194, 
    -0.9161352, -0.77194, -0.6276093, -0.4831437, -0.3385442, -0.1938114, 
    -0.04894607, 0.09605089, 0.2411787, 0.3864367, 0.5318239, 0.6773396, 
    0.8229828, 0.968753, 1.114649, 1.26067, 1.406816, 1.553085, 1.699476, 
    1.84599, 1.992624, 2.139378, 2.286251, 2.433242, 2.580351, 2.727576, 
    2.874916, 3.022371, 3.16994, 3.317621, 3.465414, 3.613318, 3.761332, 
    3.909454, 4.057685, 4.206023, 4.354466, 4.503015, 4.651668, 4.800424, 
    4.949282, 5.098241, 5.2473, 5.396458, 5.545715, 5.695068, 5.844517, 
    5.994061, 6.1437, 6.293431, 6.443254, 6.593168, 6.743171, 6.893263, 
    7.043443, 7.193709, 7.344061, 7.494497, 7.645016, 7.795618, 7.9463, 
    8.097063, 8.247904, 8.398823, 8.549819, 8.700891, 8.852036, 9.003255, 
    9.154546, 9.305908, 9.457339, 9.60884, 9.760408, 9.912043, 10.06374, 
    10.21551, 10.36733, 10.51922, 10.67117, 10.82318, 10.97524, 11.12737, 
    11.27955, 11.43178, 11.58407, 11.73641, 11.8888, 12.04124, 12.19373, 
    12.34626, 12.49885, 12.65147, 12.80414, 12.95686, 13.10961, 13.26241, 
    13.41524, 13.56811, 13.72102, 13.87396, 14.02694, 14.17995, 14.33299, 
    14.48606, 14.63916, 14.79229, 14.94544, 15.09862, 15.25183, 15.40505, 
    15.5583, 15.71157, 15.86485, 16.01816, 16.17148, 16.32481, 16.47816, 
    16.63152, 16.78489, 16.93828, 17.09167, 17.24507, 17.39848, 17.55189, 
    17.7053, 17.85872, 18.01213, 18.16555, 18.31897, 18.47238, 18.62579, 
    18.7792, 18.93259, 19.08599, 19.23937, 19.39274, 19.5461, 19.69944, 
    19.85278, 20.0061, 20.1594, 20.31268, 20.46594, 20.61919, 20.77241, 
    20.92561, 21.07878, 21.23194, 21.38506, 21.53815, 21.69122, 21.84426, 
    21.99726, 22.15023, 22.30317, 22.45607, 22.60894, 22.76176, 22.91455, 
    23.0673, 23.22001, 23.37267, 23.52529, 23.67787, 23.8304, 23.98288, 
    24.13531, 24.28769, 24.44003, 24.5923, 24.74453, 24.8967, 25.04881, 
    25.20087, 25.35287, 25.50481, 25.65669, 25.8085, 25.96026, 26.11195, 
    26.26357, 26.41513, 26.56662, 26.71804, 26.86939, 27.02067, 27.17188, 
    27.32301, 27.47407, 27.62506, 27.77596, 27.92679, 28.07754, 28.22821, 
    28.3788, 28.5293, 28.67973, 28.83007, 28.98032, 29.13049, 29.28056, 
    29.43055, 29.58045, 29.73026, 29.87998, 30.0296, 30.17913, 30.32856, 
    30.4779, 30.62714, 30.77629, 30.92533, 31.07427, 31.22311, 31.37185, 
    31.52049, 31.66902, 31.81745, 31.96577, 32.11398, 32.26209, 32.41008, 
    32.55797, 32.70575, 32.85341, 33.00096, 33.1484, 33.29572, 33.44293, 
    33.59002, 33.73699, 33.88385, 34.03058, 34.1772, 34.32369, 34.47006, 
    34.61631, 34.76244, 34.90844, 35.05431, 35.20007, 35.34569, 35.49118, 
    35.63655, 35.78179, 35.9269, 36.07187, 36.21671, 36.36143, 36.506, 
    36.65045, 36.79476, 36.93893, 37.08297, 37.22687, 37.37063, 37.51426, 
    37.65774, 37.80108, 37.94429, 38.08735, 38.23027, 38.37304, 38.51568, 
    38.65816, 38.80051, 38.94271, 39.08476, 39.22667, 39.36842, 39.51003, 
    39.65149, 39.7928, 39.93396, 40.07497, 40.21583, 40.35654, 40.49709, 
    40.6375, 40.77774, 40.91784, 41.05778, 41.19756, 41.33719, 41.47666, 
    41.61597, 41.75513, 41.89413, 42.03297, 42.17165, 42.31017, 42.44854, 
    42.58673, 42.72478, 42.86266, 43.00037, 43.13792, 43.27532,
  -19.34495, -19.22367, -19.10222, -18.98058, -18.85876, -18.73676, 
    -18.61458, -18.49222, -18.36969, -18.24697, -18.12407, -18.00099, 
    -17.87773, -17.75429, -17.63067, -17.50687, -17.38289, -17.25873, 
    -17.13438, -17.00986, -16.88516, -16.76028, -16.63522, -16.50997, 
    -16.38455, -16.25895, -16.13316, -16.0072, -15.88105, -15.75473, 
    -15.62823, -15.50154, -15.37468, -15.24764, -15.12041, -14.99301, 
    -14.86543, -14.73767, -14.60973, -14.48161, -14.35331, -14.22483, 
    -14.09618, -13.96734, -13.83833, -13.70914, -13.57977, -13.45022, 
    -13.32049, -13.19059, -13.06051, -12.93025, -12.79981, -12.6692, 
    -12.53841, -12.40744, -12.2763, -12.14498, -12.01348, -11.88181, 
    -11.74996, -11.61794, -11.48574, -11.35337, -11.22082, -11.0881, 
    -10.95521, -10.82214, -10.6889, -10.55548, -10.42189, -10.28813, 
    -10.15419, -10.02009, -9.88581, -9.75136, -9.616739, -9.481948, 
    -9.346986, -9.211853, -9.076551, -8.94108, -8.80544, -8.669631, 
    -8.533653, -8.397508, -8.261195, -8.124716, -7.988069, -7.851256, 
    -7.714277, -7.577132, -7.439823, -7.302349, -7.164711, -7.026909, 
    -6.888944, -6.750815, -6.612525, -6.474073, -6.335459, -6.196685, 
    -6.05775, -5.918655, -5.779401, -5.639988, -5.500417, -5.360688, 
    -5.220802, -5.080759, -4.940559, -4.800205, -4.659695, -4.519031, 
    -4.378212, -4.237241, -4.096117, -3.95484, -3.813413, -3.671834, 
    -3.530105, -3.388227, -3.246199, -3.104023, -2.961699, -2.819229, 
    -2.676611, -2.533849, -2.390941, -2.247889, -2.104692, -1.961354, 
    -1.817873, -1.67425, -1.530486, -1.386582, -1.242539, -1.098358, 
    -0.9540378, -0.809581, -0.6649877, -0.5202588, -0.3753951, -0.2303973, 
    -0.08526612, 0.05999754, 0.2053929, 0.3509192, 0.4965756, 0.6423612, 
    0.7882753, 0.9343171, 1.080486, 1.22678, 1.3732, 1.519743, 1.66641, 
    1.8132, 1.960111, 2.107143, 2.254295, 2.401566, 2.548954, 2.69646, 
    2.844083, 2.99182, 3.139672, 3.287637, 3.435715, 3.583904, 3.732204, 
    3.880614, 4.029132, 4.177758, 4.32649, 4.475328, 4.624272, 4.773319, 
    4.922468, 5.07172, 5.221072, 5.370523, 5.520074, 5.669723, 5.819467, 
    5.969308, 6.119243, 6.269271, 6.419392, 6.569605, 6.719907, 6.870299, 
    7.02078, 7.171347, 7.322, 7.472738, 7.62356, 7.774465, 7.925451, 
    8.076518, 8.227665, 8.378889, 8.53019, 8.681568, 8.833021, 8.984548, 
    9.136147, 9.287817, 9.439557, 9.591368, 9.743245, 9.89519, 10.0472, 
    10.19928, 10.35141, 10.50361, 10.65587, 10.8082, 10.96058, 11.11301, 
    11.26551, 11.41805, 11.57066, 11.72331, 11.87602, 12.02877, 12.18158, 
    12.33443, 12.48733, 12.64027, 12.79326, 12.94629, 13.09937, 13.25248, 
    13.40563, 13.55882, 13.71205, 13.86531, 14.01861, 14.17194, 14.3253, 
    14.47869, 14.63211, 14.78556, 14.93903, 15.09253, 15.24605, 15.3996, 
    15.55317, 15.70676, 15.86037, 16.01399, 16.16763, 16.32129, 16.47496, 
    16.62865, 16.78234, 16.93605, 17.08976, 17.24348, 17.39721, 17.55094, 
    17.70468, 17.85842, 18.01216, 18.1659, 18.31964, 18.47338, 18.62711, 
    18.78083, 18.93456, 19.08827, 19.24197, 19.39566, 19.54935, 19.70302, 
    19.85667, 20.01031, 20.16393, 20.31754, 20.47112, 20.62469, 20.77823, 
    20.93175, 21.08525, 21.23872, 21.39216, 21.54558, 21.69897, 21.85232, 
    22.00565, 22.15894, 22.31219, 22.46541, 22.6186, 22.77174, 22.92485, 
    23.07792, 23.23094, 23.38392, 23.53686, 23.68975, 23.8426, 23.9954, 
    24.14814, 24.30084, 24.45349, 24.60608, 24.75862, 24.9111, 25.06353, 
    25.2159, 25.36822, 25.52047, 25.67266, 25.82479, 25.97685, 26.12885, 
    26.28078, 26.43265, 26.58445, 26.73618, 26.88784, 27.03943, 27.19094, 
    27.34238, 27.49375, 27.64504, 27.79625, 27.94738, 28.09844, 28.24941, 
    28.4003, 28.55111, 28.70184, 28.85248, 29.00303, 29.1535, 29.30387, 
    29.45416, 29.60436, 29.75447, 29.90448, 30.0544, 30.20423, 30.35396, 
    30.50359, 30.65312, 30.80256, 30.9519, 31.10113, 31.25027, 31.3993, 
    31.54822, 31.69704, 31.84576, 31.99437, 32.14287, 32.29126, 32.43954, 
    32.58772, 32.73577, 32.88372, 33.03156, 33.17928, 33.32688, 33.47437, 
    33.62174, 33.76899, 33.91612, 34.06314, 34.21003, 34.3568, 34.50344, 
    34.64997, 34.79637, 34.94265, 35.08879, 35.23481, 35.38071, 35.52647, 
    35.67211, 35.81762, 35.96299, 36.10823, 36.25334, 36.39832, 36.54316, 
    36.68787, 36.83244, 36.97688, 37.12117, 37.26534, 37.40936, 37.55324, 
    37.69698, 37.84058, 37.98404, 38.12735, 38.27053, 38.41356, 38.55644, 
    38.69918, 38.84177, 38.98422, 39.12652, 39.26868, 39.41068, 39.55254, 
    39.69424, 39.83579, 39.9772, 40.11845, 40.25955, 40.4005, 40.54129, 
    40.68193, 40.82242, 40.96275, 41.10292, 41.24294, 41.3828, 41.52251, 
    41.66205, 41.80144, 41.94067, 42.07974, 42.21865, 42.3574, 42.49598, 
    42.63441, 42.77267, 42.91078, 43.04872, 43.18649, 43.3241,
  -19.41037, -19.28895, -19.16736, -19.04558, -18.92362, -18.80149, 
    -18.67916, -18.55667, -18.43398, -18.31112, -18.18808, -18.06486, 
    -17.94145, -17.81786, -17.6941, -17.57015, -17.44602, -17.3217, 
    -17.19721, -17.07254, -16.94768, -16.82265, -16.69743, -16.57203, 
    -16.44645, -16.32069, -16.19475, -16.06863, -15.94232, -15.81584, 
    -15.68917, -15.56233, -15.4353, -15.30809, -15.18071, -15.05314, 
    -14.92539, -14.79746, -14.66935, -14.54106, -14.41259, -14.28395, 
    -14.15512, -14.02611, -13.89692, -13.76755, -13.63801, -13.50828, 
    -13.37838, -13.24829, -13.11803, -12.98759, -12.85698, -12.72618, 
    -12.59521, -12.46406, -12.33273, -12.20122, -12.06954, -11.93768, 
    -11.80564, -11.67343, -11.54104, -11.40848, -11.27574, -11.14282, 
    -11.00973, -10.87647, -10.74303, -10.60942, -10.47563, -10.34167, 
    -10.20753, -10.07322, -9.938744, -9.80409, -9.669266, -9.534269, 
    -9.399101, -9.263762, -9.128252, -8.992572, -8.856722, -8.720701, 
    -8.584513, -8.448154, -8.311628, -8.174933, -8.038071, -7.901042, 
    -7.763845, -7.626482, -7.488954, -7.351259, -7.213399, -7.075376, 
    -6.937187, -6.798835, -6.660319, -6.521641, -6.382801, -6.243798, 
    -6.104635, -5.96531, -5.825825, -5.686181, -5.546377, -5.406415, 
    -5.266294, -5.126015, -4.985579, -4.844988, -4.70424, -4.563336, 
    -4.422278, -4.281065, -4.139699, -3.99818, -3.856509, -3.714686, 
    -3.572711, -3.430586, -3.288311, -3.145887, -3.003314, -2.860594, 
    -2.717726, -2.574711, -2.43155, -2.288244, -2.144794, -2.001199, 
    -1.857462, -1.713582, -1.569561, -1.425398, -1.281095, -1.136653, 
    -0.9920714, -0.8473522, -0.7024958, -0.5575028, -0.4123741, -0.2671105, 
    -0.1217127, 0.02381838, 0.169482, 0.3152774, 0.4612038, 0.6072602, 
    0.7534459, 0.89976, 1.046202, 1.19277, 1.339465, 1.486284, 1.633227, 
    1.780294, 1.927483, 2.074794, 2.222226, 2.369777, 2.517447, 2.665234, 
    2.813139, 2.96116, 3.109296, 3.257546, 3.405909, 3.554384, 3.702971, 
    3.851669, 4.000475, 4.14939, 4.298413, 4.447542, 4.596776, 4.746115, 
    4.895557, 5.045102, 5.194748, 5.344494, 5.49434, 5.644284, 5.794326, 
    5.944463, 6.094696, 6.245023, 6.395443, 6.545955, 6.696558, 6.847251, 
    6.998033, 7.148902, 7.299858, 7.4509, 7.602025, 7.753234, 7.904525, 
    8.055898, 8.20735, 8.358881, 8.510489, 8.662175, 8.813935, 8.965771, 
    9.117679, 9.269658, 9.421709, 9.57383, 9.726018, 9.878274, 10.0306, 
    10.18298, 10.33543, 10.48795, 10.64052, 10.79316, 10.94585, 11.0986, 
    11.25141, 11.40427, 11.55719, 11.71016, 11.86319, 12.01626, 12.16938, 
    12.32255, 12.47577, 12.62903, 12.78234, 12.93569, 13.08908, 13.24251, 
    13.39598, 13.54949, 13.70304, 13.85662, 14.01024, 14.16389, 14.31757, 
    14.47128, 14.62503, 14.7788, 14.93259, 15.08642, 15.24026, 15.39413, 
    15.54802, 15.70193, 15.85586, 16.00981, 16.16378, 16.31776, 16.47175, 
    16.62576, 16.77978, 16.93381, 17.08784, 17.24189, 17.39594, 17.55, 
    17.70406, 17.85812, 18.01219, 18.16625, 18.32031, 18.47437, 18.62843, 
    18.78248, 18.93652, 19.09056, 19.24459, 19.3986, 19.55261, 19.7066, 
    19.86058, 20.01454, 20.16849, 20.32241, 20.47632, 20.63021, 20.78408, 
    20.93792, 21.09174, 21.24553, 21.39929, 21.55303, 21.70674, 21.86042, 
    22.01406, 22.16767, 22.32125, 22.47479, 22.6283, 22.78176, 22.93519, 
    23.08857, 23.24192, 23.39522, 23.54847, 23.70168, 23.85484, 24.00796, 
    24.16102, 24.31404, 24.467, 24.61991, 24.77276, 24.92556, 25.07831, 
    25.23099, 25.38362, 25.53618, 25.68868, 25.84113, 25.9935, 26.14581, 
    26.29806, 26.45024, 26.60235, 26.75439, 26.90636, 27.05825, 27.21008, 
    27.36182, 27.5135, 27.66509, 27.81661, 27.96805, 28.11941, 28.27069, 
    28.42189, 28.573, 28.72403, 28.87497, 29.02582, 29.17659, 29.32727, 
    29.47786, 29.62836, 29.77876, 29.92908, 30.07929, 30.22941, 30.37944, 
    30.52937, 30.6792, 30.82893, 30.97856, 31.12809, 31.27752, 31.42684, 
    31.57606, 31.72517, 31.87417, 32.02307, 32.17186, 32.32054, 32.46911, 
    32.61757, 32.76591, 32.91415, 33.06226, 33.21027, 33.35815, 33.50592, 
    33.65357, 33.80111, 33.94852, 34.09581, 34.24298, 34.39003, 34.53695, 
    34.68375, 34.83042, 34.97697, 35.12339, 35.26969, 35.41585, 35.56189, 
    35.70779, 35.85357, 35.99921, 36.14472, 36.2901, 36.43534, 36.58045, 
    36.72542, 36.87025, 37.01495, 37.15951, 37.30393, 37.44821, 37.59235, 
    37.73635, 37.88021, 38.02392, 38.1675, 38.31092, 38.4542, 38.59734, 
    38.74033, 38.88318, 39.02588, 39.16843, 39.31083, 39.45308, 39.59518, 
    39.73713, 39.87893, 40.02058, 40.16207, 40.30341, 40.4446, 40.58564, 
    40.72651, 40.86724, 41.0078, 41.14822, 41.28847, 41.42857, 41.5685, 
    41.70828, 41.8479, 41.98736, 42.12666, 42.2658, 42.40477, 42.54359, 
    42.68224, 42.82073, 42.95906, 43.09722, 43.23522, 43.37305,
  -19.47595, -19.3544, -19.23267, -19.11075, -18.98866, -18.86638, -18.74392, 
    -18.62128, -18.49845, -18.37545, -18.25226, -18.12889, -18.00534, 
    -17.88161, -17.75769, -17.63359, -17.50932, -17.38486, -17.26021, 
    -17.13539, -17.01038, -16.88519, -16.75982, -16.63426, -16.50853, 
    -16.38261, -16.25651, -16.13023, -16.00377, -15.87712, -15.75029, 
    -15.62329, -15.49609, -15.36872, -15.24117, -15.11344, -14.98552, 
    -14.85742, -14.72915, -14.60069, -14.47205, -14.34323, -14.21423, 
    -14.08504, -13.95568, -13.82614, -13.69642, -13.56652, -13.43643, 
    -13.30617, -13.17573, -13.04511, -12.91431, -12.78333, -12.65218, 
    -12.52084, -12.38933, -12.25763, -12.12576, -11.99372, -11.86149, 
    -11.72909, -11.59651, -11.46375, -11.33082, -11.19771, -11.06443, 
    -10.93096, -10.79733, -10.66352, -10.52953, -10.39537, -10.26103, 
    -10.12652, -9.991841, -9.856985, -9.721956, -9.586754, -9.451379, 
    -9.315833, -9.180115, -9.044225, -8.908164, -8.771934, -8.635532, 
    -8.49896, -8.362221, -8.22531, -8.088233, -7.950986, -7.813572, -7.67599, 
    -7.538241, -7.400326, -7.262245, -7.123998, -6.985586, -6.84701, 
    -6.708269, -6.569364, -6.430296, -6.291066, -6.151672, -6.012118, 
    -5.872402, -5.732525, -5.592488, -5.452291, -5.311936, -5.171422, 
    -5.030749, -4.889919, -4.748932, -4.60779, -4.466491, -4.325037, 
    -4.183428, -4.041666, -3.89975, -3.757682, -3.615461, -3.473089, 
    -3.330566, -3.187893, -3.045071, -2.902099, -2.75898, -2.615712, 
    -2.472298, -2.328738, -2.185033, -2.041182, -1.897188, -1.75305, 
    -1.60877, -1.464347, -1.319784, -1.17508, -1.030237, -0.8852546, 
    -0.7401342, -0.5948764, -0.4494821, -0.3039519, -0.1582868, -0.01248748, 
    0.1334452, 0.2795105, 0.4257075, 0.5720356, 0.7184936, 0.865081, 
    1.011797, 1.15864, 1.30561, 1.452706, 1.599927, 1.747271, 1.894739, 
    2.04233, 2.190042, 2.337874, 2.485826, 2.633896, 2.782084, 2.930389, 
    3.07881, 3.227346, 3.375996, 3.524758, 3.673633, 3.822619, 3.971715, 
    4.12092, 4.270234, 4.419654, 4.56918, 4.718812, 4.868548, 5.018387, 
    5.168328, 5.31837, 5.468512, 5.618753, 5.769092, 5.919528, 6.070059, 
    6.220686, 6.371406, 6.522219, 6.673123, 6.824118, 6.975202, 7.126374, 
    7.277634, 7.428979, 7.58041, 7.731925, 7.883522, 8.035201, 8.18696, 
    8.338799, 8.490715, 8.642709, 8.794779, 8.946923, 9.099141, 9.251431, 
    9.403793, 9.556226, 9.708726, 9.861295, 10.01393, 10.16663, 10.3194, 
    10.47222, 10.62511, 10.77806, 10.93107, 11.08414, 11.23726, 11.39044, 
    11.54368, 11.69697, 11.85031, 12.0037, 12.15714, 12.31063, 12.46416, 
    12.61775, 12.77137, 12.92504, 13.07876, 13.23251, 13.3863, 13.54013, 
    13.694, 13.8479, 14.00184, 14.15582, 14.30982, 14.46385, 14.61792, 
    14.77201, 14.92613, 15.08028, 15.23445, 15.38864, 15.54285, 15.69709, 
    15.85134, 16.00562, 16.15991, 16.31421, 16.46853, 16.62286, 16.7772, 
    16.93156, 17.08592, 17.24029, 17.39467, 17.54905, 17.70343, 17.85782, 
    18.01221, 18.1666, 18.32099, 18.47537, 18.62975, 18.78413, 18.9385, 
    19.09286, 19.24721, 19.40155, 19.55588, 19.7102, 19.8645, 20.01879, 
    20.17306, 20.32731, 20.48154, 20.63575, 20.78994, 20.94411, 21.09825, 
    21.25237, 21.40645, 21.56051, 21.71454, 21.86854, 22.02251, 22.17644, 
    22.33034, 22.4842, 22.63803, 22.79182, 22.94556, 23.09927, 23.25293, 
    23.40655, 23.56013, 23.71366, 23.86714, 24.02057, 24.17395, 24.32728, 
    24.48056, 24.63379, 24.78696, 24.94008, 25.09314, 25.24614, 25.39908, 
    25.55196, 25.70477, 25.85753, 26.01022, 26.16284, 26.3154, 26.46789, 
    26.62031, 26.77266, 26.92494, 27.07715, 27.22928, 27.38134, 27.53332, 
    27.68522, 27.83705, 27.9888, 28.14046, 28.29205, 28.44355, 28.59497, 
    28.7463, 28.89754, 29.0487, 29.19977, 29.35075, 29.50164, 29.65244, 
    29.80315, 29.95376, 30.10427, 30.2547, 30.40502, 30.55524, 30.70537, 
    30.8554, 31.00532, 31.15515, 31.30486, 31.45448, 31.60399, 31.75339, 
    31.90269, 32.05188, 32.20095, 32.34992, 32.49878, 32.64753, 32.79616, 
    32.94468, 33.09308, 33.24136, 33.38953, 33.53759, 33.68552, 33.83333, 
    33.98103, 34.1286, 34.27604, 34.42337, 34.57057, 34.71765, 34.8646, 
    35.01142, 35.15812, 35.30468, 35.45112, 35.59743, 35.7436, 35.88965, 
    36.03556, 36.18134, 36.32698, 36.47249, 36.61786, 36.7631, 36.9082, 
    37.05316, 37.19798, 37.34266, 37.4872, 37.6316, 37.77586, 37.91998, 
    38.06395, 38.20778, 38.35146, 38.495, 38.63839, 38.78163, 38.92472, 
    39.06767, 39.21047, 39.35312, 39.49562, 39.63797, 39.78017, 39.92221, 
    40.0641, 40.20584, 40.34742, 40.48885, 40.63013, 40.77124, 40.91221, 
    41.05301, 41.19366, 41.33415, 41.47448, 41.61465, 41.75466, 41.89451, 
    42.0342, 42.17373, 42.3131, 42.4523, 42.59135, 42.73022, 42.86894, 
    43.00749, 43.14588, 43.2841, 43.42215,
  -19.5417, -19.42002, -19.29815, -19.17609, -19.05386, -18.93144, -18.80884, 
    -18.68606, -18.56309, -18.43995, -18.31661, -18.1931, -18.0694, 
    -17.94552, -17.82146, -17.69721, -17.57279, -17.44818, -17.32338, 
    -17.1984, -17.07324, -16.9479, -16.82237, -16.69666, -16.57077, -16.4447, 
    -16.31844, -16.192, -16.06538, -15.93857, -15.81158, -15.68441, 
    -15.55706, -15.42952, -15.30181, -15.17391, -15.04582, -14.91756, 
    -14.78911, -14.66048, -14.53167, -14.40268, -14.27351, -14.14415, 
    -14.01462, -13.8849, -13.755, -13.62492, -13.49466, -13.36422, -13.2336, 
    -13.1028, -12.97182, -12.84065, -12.70931, -12.57779, -12.44609, 
    -12.31421, -12.18216, -12.04992, -11.91751, -11.78491, -11.65214, 
    -11.51919, -11.38607, -11.25276, -11.11928, -10.98563, -10.85179, 
    -10.71778, -10.5836, -10.44924, -10.3147, -10.17999, -10.0451, -9.910044, 
    -9.77481, -9.639401, -9.50382, -9.368067, -9.23214, -9.096041, -8.959769, 
    -8.823327, -8.686713, -8.549929, -8.412973, -8.275848, -8.138554, 
    -8.00109, -7.863458, -7.725657, -7.587688, -7.449552, -7.311248, 
    -7.172779, -7.034142, -6.895341, -6.756374, -6.617242, -6.477947, 
    -6.338487, -6.198864, -6.059079, -5.919131, -5.779022, -5.638752, 
    -5.49832, -5.357729, -5.216979, -5.076069, -4.935, -4.793775, -4.652391, 
    -4.510851, -4.369155, -4.227304, -4.085298, -3.943137, -3.800823, 
    -3.658355, -3.515736, -3.372964, -3.230042, -3.086969, -2.943746, 
    -2.800374, -2.656854, -2.513186, -2.369371, -2.22541, -2.081302, 
    -1.93705, -1.792654, -1.648114, -1.503432, -1.358607, -1.213642, 
    -1.068535, -0.9232891, -0.777904, -0.6323807, -0.4867199, -0.3409225, 
    -0.1949892, -0.04892096, 0.09728158, 0.2436175, 0.3900861, 0.5366864, 
    0.6834176, 0.8302789, 0.9772695, 1.124388, 1.271635, 1.419008, 1.566507, 
    1.714131, 1.861878, 2.009749, 2.157742, 2.305856, 2.454091, 2.602445, 
    2.750917, 2.899508, 3.048214, 3.197037, 3.345974, 3.495025, 3.644188, 
    3.793464, 3.94285, 4.092346, 4.241951, 4.391664, 4.541484, 4.69141, 
    4.84144, 4.991574, 5.141811, 5.29215, 5.442589, 5.593128, 5.743765, 
    5.8945, 6.045332, 6.196259, 6.34728, 6.498394, 6.649601, 6.800899, 
    6.952287, 7.103763, 7.255327, 7.406978, 7.558715, 7.710536, 7.86244, 
    8.014426, 8.166493, 8.318641, 8.470867, 8.62317, 8.77555, 8.928005, 
    9.080535, 9.233137, 9.385811, 9.538555, 9.69137, 9.844252, 9.997201, 
    10.15022, 10.3033, 10.45644, 10.60964, 10.76291, 10.91624, 11.06962, 
    11.22306, 11.37656, 11.53011, 11.68372, 11.83738, 11.99109, 12.14485, 
    12.29866, 12.45252, 12.60642, 12.76037, 12.91436, 13.06839, 13.22247, 
    13.37658, 13.53073, 13.68493, 13.83915, 13.99341, 14.14771, 14.30204, 
    14.4564, 14.61078, 14.7652, 14.91965, 15.07411, 15.22861, 15.38313, 
    15.53767, 15.69223, 15.84681, 16.00141, 16.15602, 16.31065, 16.4653, 
    16.61995, 16.77462, 16.9293, 17.08399, 17.23869, 17.39339, 17.5481, 
    17.70281, 17.85752, 18.01224, 18.16695, 18.32166, 18.47638, 18.63108, 
    18.78579, 18.94048, 19.09517, 19.24985, 19.40451, 19.55917, 19.71381, 
    19.86844, 20.02305, 20.17765, 20.33222, 20.48678, 20.64132, 20.79583, 
    20.95032, 21.10479, 21.25923, 21.41364, 21.56802, 21.72238, 21.8767, 
    22.03099, 22.18525, 22.33947, 22.49365, 22.6478, 22.80191, 22.95598, 
    23.11, 23.26399, 23.41793, 23.57183, 23.72567, 23.87947, 24.03323, 
    24.18693, 24.34058, 24.49418, 24.64772, 24.80121, 24.95465, 25.10802, 
    25.26134, 25.41459, 25.56779, 25.72092, 25.87399, 26.027, 26.17994, 
    26.33281, 26.48561, 26.63834, 26.79101, 26.9436, 27.09612, 27.24856, 
    27.40093, 27.55322, 27.70543, 27.85757, 28.00962, 28.16159, 28.31349, 
    28.46529, 28.61702, 28.76865, 28.9202, 29.07167, 29.22304, 29.37432, 
    29.52552, 29.67661, 29.82762, 29.97853, 30.12935, 30.28007, 30.43069, 
    30.58121, 30.73164, 30.88196, 31.03218, 31.1823, 31.33231, 31.48222, 
    31.63202, 31.78172, 31.93131, 32.08079, 32.23016, 32.37941, 32.52856, 
    32.67759, 32.82651, 32.97532, 33.124, 33.27258, 33.42103, 33.56937, 
    33.71758, 33.86568, 34.01365, 34.1615, 34.30923, 34.45683, 34.60431, 
    34.75167, 34.89889, 35.04599, 35.19296, 35.3398, 35.48651, 35.63309, 
    35.77954, 35.92585, 36.07204, 36.21808, 36.36399, 36.50977, 36.65541, 
    36.80091, 36.94627, 37.0915, 37.23658, 37.38153, 37.52633, 37.67099, 
    37.81551, 37.95988, 38.10411, 38.24819, 38.39213, 38.53592, 38.67957, 
    38.82306, 38.96641, 39.10961, 39.25266, 39.39556, 39.53831, 39.6809, 
    39.82335, 39.96563, 40.10777, 40.24975, 40.39158, 40.53325, 40.67477, 
    40.81612, 40.95732, 41.09837, 41.23925, 41.37998, 41.52055, 41.66095, 
    41.8012, 41.94128, 42.0812, 42.22096, 42.36056, 42.49999, 42.63926, 
    42.77837, 42.91731, 43.05608, 43.19469, 43.33314, 43.47141,
  -19.60763, -19.48581, -19.3638, -19.24161, -19.11923, -18.99668, -18.87394, 
    -18.75101, -18.6279, -18.50461, -18.38114, -18.25748, -18.13364, 
    -18.00961, -17.8854, -17.76101, -17.63643, -17.51167, -17.38672, 
    -17.26159, -17.13628, -17.01078, -16.88511, -16.75924, -16.63319, 
    -16.50696, -16.38054, -16.25395, -16.12716, -16.0002, -15.87305, 
    -15.74571, -15.6182, -15.4905, -15.36261, -15.23455, -15.1063, -14.97786, 
    -14.84925, -14.72045, -14.59147, -14.46231, -14.33296, -14.20343, 
    -14.07372, -13.94383, -13.81375, -13.68349, -13.55306, -13.42244, 
    -13.29164, -13.16065, -13.02949, -12.89815, -12.76662, -12.63492, 
    -12.50303, -12.37097, -12.23872, -12.10629, -11.97369, -11.84091, 
    -11.70794, -11.5748, -11.44148, -11.30799, -11.17431, -11.04046, 
    -10.90643, -10.77222, -10.63783, -10.50327, -10.36854, -10.23362, 
    -10.09853, -9.963268, -9.827828, -9.692215, -9.556427, -9.420465, 
    -9.284328, -9.14802, -9.011538, -8.874884, -8.738057, -8.601058, 
    -8.463889, -8.326548, -8.189036, -8.051355, -7.913504, -7.775484, 
    -7.637294, -7.498936, -7.360411, -7.221717, -7.082857, -6.94383, 
    -6.804636, -6.665277, -6.525753, -6.386065, -6.246212, -6.106195, 
    -5.966015, -5.825673, -5.685168, -5.544502, -5.403675, -5.262687, 
    -5.12154, -4.980233, -4.838767, -4.697143, -4.555361, -4.413423, 
    -4.271327, -4.129077, -3.986671, -3.84411, -3.701396, -3.558528, 
    -3.415507, -3.272335, -3.12901, -2.985536, -2.841911, -2.698137, 
    -2.554214, -2.410144, -2.265926, -2.121561, -1.977051, -1.832396, 
    -1.687596, -1.542652, -1.397566, -1.252337, -1.106967, -0.9614565, 
    -0.815806, -0.6700164, -0.5240885, -0.3780231, -0.231821, -0.08548295, 
    0.06099017, 0.2075976, 0.3543384, 0.5012118, 0.6482171, 0.7953532, 
    0.9426194, 1.090015, 1.237538, 1.38519, 1.532967, 1.680871, 1.828899, 
    1.977051, 2.125326, 2.273724, 2.422242, 2.57088, 2.719638, 2.868514, 
    3.017508, 3.166618, 3.315843, 3.465183, 3.614636, 3.764203, 3.91388, 
    4.063668, 4.213566, 4.363572, 4.513686, 4.663906, 4.814232, 4.964663, 
    5.115196, 5.265832, 5.41657, 5.567408, 5.718345, 5.86938, 6.020513, 
    6.171741, 6.323064, 6.474482, 6.625992, 6.777594, 6.929286, 7.081068, 
    7.232937, 7.384895, 7.536938, 7.689067, 7.841279, 7.993574, 8.14595, 
    8.298408, 8.450944, 8.603559, 8.756249, 8.909017, 9.061858, 9.214773, 
    9.367761, 9.520819, 9.673947, 9.827145, 9.980409, 10.13374, 10.28714, 
    10.44059, 10.59412, 10.7477, 10.90134, 11.05505, 11.20881, 11.36263, 
    11.5165, 11.67042, 11.8244, 11.97843, 12.13251, 12.28664, 12.44082, 
    12.59505, 12.74932, 12.90363, 13.05799, 13.21239, 13.36682, 13.5213, 
    13.67582, 13.83037, 13.98495, 14.13957, 14.29422, 14.44891, 14.60362, 
    14.75836, 14.91313, 15.06793, 15.22275, 15.37759, 15.53246, 15.68735, 
    15.84225, 15.99718, 16.15212, 16.30708, 16.46205, 16.61703, 16.77203, 
    16.92703, 17.08205, 17.23707, 17.39211, 17.54714, 17.70218, 17.85722, 
    18.01226, 18.1673, 18.32235, 18.47738, 18.63242, 18.78745, 18.94247, 
    19.09748, 19.25249, 19.40748, 19.56247, 19.71744, 19.87239, 20.02733, 
    20.18225, 20.33716, 20.49204, 20.6469, 20.80174, 20.95656, 21.11135, 
    21.26612, 21.42085, 21.57556, 21.73024, 21.88489, 22.0395, 22.19408, 
    22.34863, 22.50314, 22.65761, 22.81204, 22.96643, 23.12078, 23.27509, 
    23.42935, 23.58357, 23.73774, 23.89186, 24.04593, 24.19996, 24.35393, 
    24.50785, 24.66171, 24.81552, 24.96927, 25.12296, 25.2766, 25.43017, 
    25.58368, 25.73713, 25.89052, 26.04384, 26.19709, 26.35028, 26.5034, 
    26.65644, 26.80942, 26.96232, 27.11515, 27.26791, 27.42059, 27.57319, 
    27.72571, 27.87816, 28.03052, 28.1828, 28.335, 28.48712, 28.63915, 
    28.79109, 28.94295, 29.09472, 29.24639, 29.39798, 29.54948, 29.70088, 
    29.85219, 30.0034, 30.15452, 30.30554, 30.45646, 30.60728, 30.758, 
    30.90862, 31.05914, 31.20955, 31.35986, 31.51007, 31.66016, 31.81015, 
    31.96003, 32.1098, 32.25946, 32.40901, 32.55845, 32.70777, 32.85698, 
    33.00607, 33.15504, 33.3039, 33.45264, 33.60126, 33.74976, 33.89814, 
    34.04639, 34.19453, 34.34253, 34.49042, 34.63818, 34.7858, 34.93331, 
    35.08068, 35.22793, 35.37505, 35.52203, 35.66888, 35.8156, 35.96219, 
    36.10864, 36.25496, 36.40114, 36.54718, 36.69309, 36.83886, 36.98448, 
    37.12997, 37.27532, 37.42052, 37.56559, 37.71051, 37.85529, 37.99992, 
    38.14441, 38.28875, 38.43294, 38.57699, 38.72089, 38.86464, 39.00824, 
    39.15169, 39.29499, 39.43814, 39.58114, 39.72398, 39.86667, 40.00921, 
    40.15159, 40.29382, 40.43589, 40.5778, 40.71955, 40.86116, 41.00259, 
    41.14388, 41.285, 41.42596, 41.56676, 41.70741, 41.84789, 41.9882, 
    42.12835, 42.26834, 42.40817, 42.54784, 42.68733, 42.82666, 42.96583, 
    43.10483, 43.24367, 43.38234, 43.52083,
  -19.67373, -19.55177, -19.42962, -19.30729, -19.18478, -19.06209, 
    -18.93921, -18.81614, -18.69289, -18.56945, -18.44584, -18.32203, 
    -18.19805, -18.07387, -17.94951, -17.82497, -17.70025, -17.57533, 
    -17.45024, -17.32496, -17.19949, -17.07384, -16.94801, -16.82199, 
    -16.69578, -16.5694, -16.44282, -16.31606, -16.18912, -16.06199, 
    -15.93468, -15.80719, -15.67951, -15.55164, -15.42359, -15.29536, 
    -15.16694, -15.03834, -14.90956, -14.78059, -14.65144, -14.5221, 
    -14.39258, -14.26288, -14.133, -14.00293, -13.87268, -13.74224, 
    -13.61163, -13.48083, -13.34984, -13.21868, -13.08734, -12.95581, 
    -12.8241, -12.69221, -12.56014, -12.42789, -12.29545, -12.16284, 
    -12.03004, -11.89707, -11.76392, -11.63058, -11.49707, -11.36338, 
    -11.2295, -11.09546, -10.96123, -10.82682, -10.69224, -10.55747, 
    -10.42254, -10.28742, -10.15213, -10.01666, -9.881014, -9.745194, 
    -9.609199, -9.473028, -9.336683, -9.200164, -9.063471, -8.926604, 
    -8.789564, -8.652351, -8.514967, -8.37741, -8.239681, -8.101782, 
    -7.963712, -7.825471, -7.687061, -7.548481, -7.409732, -7.270815, 
    -7.13173, -6.992477, -6.853057, -6.71347, -6.573717, -6.433799, 
    -6.293715, -6.153467, -6.013054, -5.872478, -5.731739, -5.590837, 
    -5.449774, -5.308548, -5.167162, -5.025616, -4.88391, -4.742045, 
    -4.600021, -4.457839, -4.3155, -4.173004, -4.030352, -3.887545, 
    -3.744582, -3.601465, -3.458195, -3.314772, -3.171196, -3.027469, 
    -2.883591, -2.739563, -2.595384, -2.451057, -2.306582, -2.16196, 
    -2.01719, -1.872275, -1.727215, -1.582009, -1.43666, -1.291168, 
    -1.145534, -0.999758, -0.8538413, -0.7077847, -0.5615889, -0.4152547, 
    -0.2687829, -0.1221744, 0.02457009, 0.1714497, 0.3184636, 0.465611, 
    0.612891, 0.7603027, 0.9078454, 1.055518, 1.20332, 1.35125, 1.499308, 
    1.647492, 1.795801, 1.944236, 2.092794, 2.241475, 2.390277, 2.539201, 
    2.688245, 2.837408, 2.98669, 3.136088, 3.285603, 3.435232, 3.584976, 
    3.734834, 3.884804, 4.034885, 4.185076, 4.335377, 4.485785, 4.636302, 
    4.786924, 4.937652, 5.088483, 5.239418, 5.390455, 5.541593, 5.69283, 
    5.844167, 5.995601, 6.147132, 6.298759, 6.45048, 6.602294, 6.754201, 
    6.906199, 7.058287, 7.210464, 7.362729, 7.51508, 7.667517, 7.820039, 
    7.972643, 8.12533, 8.278098, 8.430945, 8.583872, 8.736876, 8.889956, 
    9.043111, 9.196341, 9.349642, 9.503016, 9.656459, 9.809972, 9.963552, 
    10.1172, 10.27091, 10.42469, 10.57853, 10.73243, 10.8864, 11.04042, 
    11.1945, 11.34864, 11.50283, 11.65708, 11.81138, 11.96573, 12.12013, 
    12.27458, 12.42909, 12.58363, 12.73823, 12.89286, 13.04754, 13.20227, 
    13.35703, 13.51183, 13.66667, 13.82155, 13.97646, 14.1314, 14.28638, 
    14.44139, 14.59643, 14.7515, 14.9066, 15.06172, 15.21687, 15.37204, 
    15.52723, 15.68245, 15.83768, 15.99293, 16.1482, 16.30349, 16.45879, 
    16.6141, 16.76943, 16.92476, 17.0801, 17.23546, 17.39082, 17.54618, 
    17.70155, 17.85692, 18.01229, 18.16766, 18.32303, 18.4784, 18.63376, 
    18.78912, 18.94447, 19.09981, 19.25514, 19.41047, 19.56578, 19.72108, 
    19.87636, 20.03163, 20.18688, 20.34211, 20.49732, 20.65251, 20.80768, 
    20.96282, 21.11794, 21.27303, 21.42809, 21.58313, 21.73813, 21.89311, 
    22.04805, 22.20296, 22.35783, 22.51266, 22.66746, 22.82221, 22.97693, 
    23.1316, 23.28623, 23.44082, 23.59536, 23.74985, 23.90429, 24.05869, 
    24.21303, 24.36733, 24.52157, 24.67575, 24.82988, 24.98395, 25.13796, 
    25.29192, 25.44581, 25.59964, 25.75341, 25.90711, 26.06075, 26.21432, 
    26.36782, 26.52125, 26.67461, 26.8279, 26.98112, 27.13426, 27.28733, 
    27.44032, 27.59324, 27.74607, 27.89883, 28.0515, 28.20409, 28.3566, 
    28.50903, 28.66136, 28.81361, 28.96578, 29.11785, 29.26983, 29.42173, 
    29.57353, 29.72523, 29.87684, 30.02836, 30.17978, 30.3311, 30.48232, 
    30.63344, 30.78446, 30.93538, 31.0862, 31.23691, 31.38751, 31.53801, 
    31.68841, 31.83869, 31.98886, 32.13893, 32.28888, 32.43872, 32.58844, 
    32.73806, 32.88755, 33.03693, 33.1862, 33.33534, 33.48436, 33.63327, 
    33.78205, 33.93071, 34.07925, 34.22767, 34.37596, 34.52412, 34.67216, 
    34.82007, 34.96785, 35.1155, 35.26302, 35.41042, 35.55767, 35.7048, 
    35.8518, 35.99865, 36.14537, 36.29196, 36.43841, 36.58472, 36.7309, 
    36.87693, 37.02283, 37.16858, 37.31419, 37.45966, 37.60499, 37.75017, 
    37.89521, 38.0401, 38.18484, 38.32944, 38.4739, 38.6182, 38.76236, 
    38.90636, 39.05021, 39.19392, 39.33747, 39.48087, 39.62411, 39.76721, 
    39.91014, 40.05293, 40.19556, 40.33803, 40.48034, 40.6225, 40.7645, 
    40.90634, 41.04802, 41.18954, 41.3309, 41.4721, 41.61314, 41.75401, 
    41.89473, 42.03527, 42.17566, 42.31588, 42.45594, 42.59584, 42.73556, 
    42.87512, 43.01451, 43.15374, 43.2928, 43.43169, 43.57042,
  -19.74, -19.6179, -19.49562, -19.37316, -19.2505, -19.12767, -19.00465, 
    -18.88144, -18.75805, -18.63447, -18.51071, -18.38676, -18.26263, 
    -18.13831, -18.0138, -17.88911, -17.76424, -17.63918, -17.51393, 
    -17.3885, -17.26288, -17.13708, -17.01109, -16.88491, -16.75855, 
    -16.63201, -16.50527, -16.37836, -16.25126, -16.12397, -15.99649, 
    -15.86884, -15.74099, -15.61296, -15.48475, -15.35635, -15.22777, 
    -15.099, -14.97004, -14.84091, -14.71158, -14.58208, -14.45238, 
    -14.32251, -14.19245, -14.0622, -13.93178, -13.80116, -13.67037, 
    -13.53939, -13.40823, -13.27688, -13.14536, -13.01364, -12.88175, 
    -12.74968, -12.61742, -12.48498, -12.35236, -12.21955, -12.08657, 
    -11.9534, -11.82006, -11.68653, -11.55282, -11.41894, -11.28487, 
    -11.15062, -11.0162, -10.88159, -10.74681, -10.61185, -10.47671, 
    -10.34139, -10.20589, -10.07022, -9.934367, -9.79834, -9.662137, 
    -9.525758, -9.389203, -9.252474, -9.115569, -8.97849, -8.841236, 
    -8.703809, -8.566209, -8.428435, -8.29049, -8.152371, -8.014082, 
    -7.875621, -7.736989, -7.598187, -7.459215, -7.320074, -7.180763, 
    -7.041284, -6.901636, -6.761821, -6.62184, -6.48169, -6.341376, 
    -6.200895, -6.06025, -5.919439, -5.778465, -5.637328, -5.496027, 
    -5.354564, -5.212939, -5.071153, -4.929206, -4.787099, -4.644832, 
    -4.502407, -4.359823, -4.217081, -4.074183, -3.931128, -3.787917, 
    -3.64455, -3.50103, -3.357355, -3.213527, -3.069547, -2.925415, 
    -2.781131, -2.636697, -2.492113, -2.34738, -2.202499, -2.05747, 
    -1.912294, -1.766972, -1.621504, -1.475892, -1.330136, -1.184236, 
    -1.038194, -0.8920108, -0.7456864, -0.5992219, -0.4526182, -0.305876, 
    -0.1589962, -0.01197959, 0.135173, 0.2824608, 0.4298829, 0.5774385, 
    0.7251267, 0.8729466, 1.020897, 1.168978, 1.317188, 1.465526, 1.613992, 
    1.762584, 1.911301, 2.060143, 2.209109, 2.358197, 2.507407, 2.656738, 
    2.806189, 2.955759, 3.105446, 3.255251, 3.405172, 3.555208, 3.705358, 
    3.855621, 4.005995, 4.156481, 4.307077, 4.457782, 4.608595, 4.759515, 
    4.910541, 5.061671, 5.212905, 5.364243, 5.515681, 5.667221, 5.81886, 
    5.970597, 6.122431, 6.274362, 6.426388, 6.578508, 6.730721, 6.883026, 
    7.035421, 7.187906, 7.340479, 7.49314, 7.645886, 7.798718, 7.951634, 
    8.104632, 8.257712, 8.410872, 8.564112, 8.717429, 8.870823, 9.024293, 
    9.177837, 9.331454, 9.485144, 9.638905, 9.792734, 9.946632, 10.1006, 
    10.25463, 10.40873, 10.56289, 10.71711, 10.87139, 11.02573, 11.18013, 
    11.33459, 11.48911, 11.64368, 11.7983, 11.95298, 12.1077, 12.26248, 
    12.4173, 12.57218, 12.72709, 12.88205, 13.03706, 13.19211, 13.3472, 
    13.50232, 13.65749, 13.81269, 13.96793, 14.1232, 14.27851, 14.43385, 
    14.58921, 14.74461, 14.90004, 15.05549, 15.21096, 15.36646, 15.52199, 
    15.67753, 15.83309, 15.98867, 16.14427, 16.29989, 16.45551, 16.61116, 
    16.76681, 16.92248, 17.07815, 17.23383, 17.38952, 17.54522, 17.70091, 
    17.85661, 18.01231, 18.16802, 18.32372, 18.47941, 18.63511, 18.79079, 
    18.94647, 19.10215, 19.25781, 19.41346, 19.5691, 19.72473, 19.88034, 
    20.03594, 20.19152, 20.34708, 20.50262, 20.65814, 20.81363, 20.9691, 
    21.12455, 21.27997, 21.43536, 21.59073, 21.74606, 21.90136, 22.05663, 
    22.21186, 22.36706, 22.52222, 22.67734, 22.83242, 22.98746, 23.14246, 
    23.29742, 23.45233, 23.60719, 23.76201, 23.91678, 24.0715, 24.22616, 
    24.38078, 24.53534, 24.68984, 24.84429, 24.99869, 25.15302, 25.30729, 
    25.4615, 25.61565, 25.76974, 25.92376, 26.07772, 26.2316, 26.38542, 
    26.53917, 26.69285, 26.84646, 26.99999, 27.15345, 27.30683, 27.46013, 
    27.61336, 27.76651, 27.91957, 28.07256, 28.22546, 28.37828, 28.53102, 
    28.68366, 28.83622, 28.98869, 29.14107, 29.29336, 29.44556, 29.59767, 
    29.74968, 29.90159, 30.05341, 30.20513, 30.35676, 30.50828, 30.6597, 
    30.81102, 30.96224, 31.11336, 31.26436, 31.41527, 31.56606, 31.71675, 
    31.86733, 32.0178, 32.16816, 32.3184, 32.46853, 32.61855, 32.76845, 
    32.91824, 33.06791, 33.21746, 33.36689, 33.5162, 33.66539, 33.81446, 
    33.96341, 34.11223, 34.26093, 34.4095, 34.55795, 34.70626, 34.85445, 
    35.00251, 35.15044, 35.29824, 35.44591, 35.59344, 35.74085, 35.88811, 
    36.03524, 36.18224, 36.3291, 36.47582, 36.6224, 36.76884, 36.91515, 
    37.06131, 37.20732, 37.3532, 37.49894, 37.64452, 37.78997, 37.93527, 
    38.08042, 38.22543, 38.37029, 38.515, 38.65955, 38.80396, 38.94822, 
    39.09233, 39.23629, 39.38009, 39.52374, 39.66724, 39.81058, 39.95377, 
    40.0968, 40.23967, 40.38239, 40.52495, 40.66735, 40.80959, 40.95167, 
    41.09359, 41.23535, 41.37695, 41.51839, 41.65966, 41.80078, 41.94172, 
    42.08251, 42.22313, 42.36358, 42.50387, 42.64399, 42.78395, 42.92374, 
    43.06336, 43.20281, 43.34209, 43.48121, 43.62016,
  -19.80644, -19.68421, -19.56179, -19.43919, -19.3164, -19.19343, -19.07026, 
    -18.94692, -18.82338, -18.69966, -18.57576, -18.45166, -18.32738, 
    -18.20292, -18.07827, -17.95343, -17.82841, -17.70319, -17.5778, 
    -17.45221, -17.32644, -17.20049, -17.07434, -16.94801, -16.8215, 
    -16.69479, -16.5679, -16.44083, -16.31356, -16.18612, -16.05848, 
    -15.93066, -15.80265, -15.67446, -15.54608, -15.41751, -15.28876, 
    -15.15983, -15.0307, -14.90139, -14.7719, -14.64222, -14.51236, 
    -14.38231, -14.25207, -14.12165, -13.99105, -13.86026, -13.72929, 
    -13.59813, -13.46678, -13.33526, -13.20355, -13.07165, -12.93958, 
    -12.80732, -12.67487, -12.54224, -12.40944, -12.27644, -12.14327, 
    -12.00991, -11.87637, -11.74265, -11.60875, -11.47467, -11.34041, 
    -11.20596, -11.07134, -10.93653, -10.80155, -10.66639, -10.53104, 
    -10.39552, -10.25982, -10.12394, -9.987888, -9.851654, -9.715243, 
    -9.578655, -9.441891, -9.30495, -9.167833, -9.030541, -8.893074, 
    -8.755432, -8.617616, -8.479626, -8.341462, -8.203126, -8.064616, 
    -7.925934, -7.787081, -7.648056, -7.50886, -7.369493, -7.229957, 
    -7.090251, -6.950376, -6.810332, -6.670121, -6.529741, -6.389195, 
    -6.248482, -6.107603, -5.966558, -5.825348, -5.683974, -5.542436, 
    -5.400734, -5.25887, -5.116843, -4.974655, -4.832305, -4.689795, 
    -4.547125, -4.404296, -4.261309, -4.118163, -3.974859, -3.831399, 
    -3.687783, -3.544012, -3.400085, -3.256004, -3.11177, -2.967383, 
    -2.822844, -2.678153, -2.533312, -2.38832, -2.24318, -2.09789, -1.952453, 
    -1.806869, -1.661138, -1.515262, -1.369241, -1.223075, -1.076767, 
    -0.9303154, -0.7837225, -0.6369886, -0.4901146, -0.3431013, -0.1959494, 
    -0.04865981, 0.09876664, 0.2463291, 0.3940268, 0.5418587, 0.6898242, 
    0.8379222, 0.9861519, 1.134513, 1.283003, 1.431623, 1.58037, 1.729245, 
    1.878247, 2.027373, 2.176625, 2.325999, 2.475497, 2.625115, 2.774855, 
    2.924714, 3.074692, 3.224788, 3.375001, 3.525329, 3.675773, 3.826329, 
    3.976999, 4.127781, 4.278673, 4.429675, 4.580786, 4.732004, 4.883329, 
    5.03476, 5.186295, 5.337933, 5.489674, 5.641515, 5.793458, 5.945498, 
    6.097638, 6.249874, 6.402206, 6.554632, 6.707152, 6.859765, 7.012469, 
    7.165263, 7.318146, 7.471117, 7.624174, 7.777317, 7.930545, 8.083856, 
    8.237248, 8.390722, 8.544276, 8.697907, 8.851617, 9.005403, 9.159264, 
    9.313197, 9.467204, 9.621283, 9.775431, 9.929647, 10.08393, 10.23828, 
    10.3927, 10.54718, 10.70172, 10.85633, 11.01099, 11.16572, 11.3205, 
    11.47534, 11.63023, 11.78517, 11.94017, 12.09522, 12.25033, 12.40548, 
    12.56067, 12.71592, 12.8712, 13.02654, 13.18191, 13.33733, 13.49278, 
    13.64827, 13.8038, 13.95937, 14.11497, 14.27061, 14.42627, 14.58197, 
    14.73769, 14.89345, 15.04923, 15.20504, 15.36086, 15.51672, 15.67259, 
    15.82848, 15.9844, 16.14033, 16.29627, 16.45223, 16.6082, 16.76419, 
    16.92019, 17.07619, 17.2322, 17.38822, 17.54425, 17.70028, 17.85631, 
    18.01234, 18.16837, 18.3244, 18.48043, 18.63646, 18.79248, 18.94849, 
    19.10449, 19.26049, 19.41647, 19.57244, 19.7284, 19.88434, 20.04027, 
    20.19618, 20.35207, 20.50794, 20.66379, 20.81961, 20.97541, 21.13119, 
    21.28694, 21.44266, 21.59835, 21.75401, 21.90964, 22.06524, 22.2208, 
    22.37633, 22.53181, 22.68726, 22.84267, 22.99804, 23.15336, 23.30865, 
    23.46388, 23.61907, 23.77421, 23.92931, 24.08435, 24.23934, 24.39428, 
    24.54916, 24.70399, 24.85876, 25.01348, 25.16813, 25.32273, 25.47726, 
    25.63173, 25.78614, 25.94048, 26.09475, 26.24896, 26.4031, 26.55716, 
    26.71116, 26.86508, 27.01893, 27.1727, 27.3264, 27.48002, 27.63356, 
    27.78702, 27.9404, 28.0937, 28.24691, 28.40004, 28.55309, 28.70604, 
    28.85891, 29.01169, 29.16438, 29.31698, 29.46949, 29.6219, 29.77421, 
    29.92644, 30.07856, 30.23058, 30.38251, 30.53434, 30.68606, 30.83768, 
    30.9892, 31.14062, 31.29192, 31.44312, 31.59422, 31.7452, 31.89608, 
    32.04684, 32.19749, 32.34803, 32.49846, 32.64877, 32.79896, 32.94904, 
    33.099, 33.24884, 33.39856, 33.54816, 33.69764, 33.84699, 33.99622, 
    34.14533, 34.29431, 34.44317, 34.5919, 34.74049, 34.88897, 35.0373, 
    35.18551, 35.33359, 35.48153, 35.62934, 35.77702, 35.92456, 36.07197, 
    36.21923, 36.36637, 36.51336, 36.66021, 36.80692, 36.95349, 37.09992, 
    37.2462, 37.39235, 37.53835, 37.6842, 37.82991, 37.97547, 38.12088, 
    38.26615, 38.41127, 38.55623, 38.70105, 38.84572, 38.99023, 39.1346, 
    39.2788, 39.42286, 39.56676, 39.71051, 39.8541, 39.99754, 40.14082, 
    40.28394, 40.4269, 40.56971, 40.71235, 40.85483, 40.99716, 41.13932, 
    41.28132, 41.42316, 41.56483, 41.70635, 41.84769, 41.98888, 42.1299, 
    42.27075, 42.41144, 42.55196, 42.69231, 42.8325, 42.97252, 43.11236, 
    43.25204, 43.39155, 43.53089, 43.67006,
  -19.87307, -19.7507, -19.62814, -19.5054, -19.38247, -19.25936, -19.13606, 
    -19.01257, -18.88889, -18.76503, -18.64098, -18.51674, -18.39232, 
    -18.26771, -18.14291, -18.01792, -17.89275, -17.76739, -17.64184, 
    -17.5161, -17.39018, -17.26407, -17.13777, -17.01129, -16.88461, 
    -16.75775, -16.63071, -16.50347, -16.37605, -16.24844, -16.12064, 
    -15.99266, -15.86449, -15.73613, -15.60759, -15.47886, -15.34994, 
    -15.22083, -15.09154, -14.96206, -14.8324, -14.70255, -14.57251, 
    -14.44228, -14.31187, -14.18128, -14.0505, -13.91953, -13.78838, 
    -13.65704, -13.52552, -13.39381, -13.26192, -13.12984, -12.99758, 
    -12.86513, -12.7325, -12.59968, -12.46669, -12.3335, -12.20014, 
    -12.06659, -11.93286, -11.79895, -11.66485, -11.53057, -11.39612, 
    -11.26147, -11.12665, -10.99165, -10.85646, -10.7211, -10.58555, 
    -10.44983, -10.31392, -10.17784, -10.04158, -9.905138, -9.768518, 
    -9.631721, -9.494746, -9.357594, -9.220265, -9.082761, -8.945079, 
    -8.807222, -8.669189, -8.530982, -8.3926, -8.254045, -8.115314, 
    -7.976412, -7.837336, -7.698088, -7.558668, -7.419076, -7.279314, 
    -7.13938, -6.999277, -6.859004, -6.718563, -6.577952, -6.437173, 
    -6.296227, -6.155114, -6.013834, -5.872388, -5.730777, -5.589001, 
    -5.44706, -5.304956, -5.162688, -5.020258, -4.877666, -4.734912, 
    -4.591997, -4.448922, -4.305687, -4.162294, -4.018742, -3.875032, 
    -3.731165, -3.587142, -3.442963, -3.298629, -3.15414, -3.009497, 
    -2.864702, -2.719754, -2.574654, -2.429404, -2.284003, -2.138453, 
    -1.992753, -1.846906, -1.700912, -1.55477, -1.408484, -1.262052, 
    -1.115476, -0.9687562, -0.821894, -0.6748899, -0.5277448, -0.3804595, 
    -0.2330348, -0.08547149, 0.06222956, 0.2100675, 0.3580415, 0.5061507, 
    0.6543942, 0.8027712, 0.9512807, 1.099922, 1.248694, 1.397596, 1.546627, 
    1.695786, 1.845072, 1.994484, 2.144022, 2.293684, 2.443469, 2.593377, 
    2.743406, 2.893556, 3.043825, 3.194213, 3.344718, 3.495341, 3.646078, 
    3.79693, 3.947896, 4.098974, 4.250164, 4.401464, 4.552873, 4.704391, 
    4.856016, 5.007747, 5.159584, 5.311524, 5.463568, 5.615714, 5.76796, 
    5.920306, 6.072751, 6.225294, 6.377933, 6.530666, 6.683495, 6.836416, 
    6.989429, 7.142534, 7.295727, 7.449009, 7.602379, 7.755835, 7.909376, 
    8.063, 8.216707, 8.370496, 8.524364, 8.678312, 8.832338, 8.986441, 
    9.140618, 9.29487, 9.449196, 9.603593, 9.75806, 9.912598, 10.0672, 
    10.22187, 10.37661, 10.53141, 10.68628, 10.84121, 10.99619, 11.15124, 
    11.30635, 11.46151, 11.61673, 11.772, 11.92732, 12.0827, 12.23813, 
    12.3936, 12.54913, 12.7047, 12.86031, 13.01597, 13.17167, 13.32742, 
    13.4832, 13.63902, 13.79488, 13.95078, 14.10671, 14.26267, 14.41867, 
    14.5747, 14.73075, 14.88684, 15.04295, 15.19908, 15.35524, 15.51143, 
    15.66763, 15.82386, 15.9801, 16.13636, 16.29264, 16.44893, 16.60524, 
    16.76156, 16.91788, 17.07422, 17.23057, 17.38692, 17.54328, 17.69964, 
    17.856, 18.01237, 18.16873, 18.3251, 18.48146, 18.63781, 18.79416, 
    18.95051, 19.10685, 19.26317, 19.41949, 19.57579, 19.73208, 19.88836, 
    20.04461, 20.20086, 20.35708, 20.51328, 20.66946, 20.82562, 20.98175, 
    21.13786, 21.29394, 21.44999, 21.60601, 21.762, 21.91796, 22.07388, 
    22.22977, 22.38563, 22.54144, 22.69722, 22.85296, 23.00866, 23.16431, 
    23.31992, 23.47548, 23.63099, 23.78646, 23.94188, 24.09725, 24.25257, 
    24.40783, 24.56304, 24.71819, 24.87329, 25.02833, 25.18331, 25.33822, 
    25.49308, 25.64787, 25.8026, 25.95726, 26.11185, 26.26638, 26.42084, 
    26.57522, 26.72953, 26.88378, 27.03794, 27.19203, 27.34604, 27.49998, 
    27.65384, 27.80761, 27.96131, 28.11492, 28.26845, 28.42189, 28.57524, 
    28.72851, 28.88169, 29.03478, 29.18778, 29.34069, 29.4935, 29.64622, 
    29.79884, 29.95137, 30.1038, 30.25613, 30.40836, 30.56049, 30.71252, 
    30.86444, 31.01626, 31.16798, 31.31958, 31.47108, 31.62248, 31.77376, 
    31.92493, 32.07599, 32.22694, 32.37777, 32.52849, 32.6791, 32.82958, 
    32.97995, 33.1302, 33.28033, 33.43034, 33.58023, 33.73, 33.87964, 
    34.02916, 34.17855, 34.32782, 34.47696, 34.62597, 34.77485, 34.9236, 
    35.07222, 35.22071, 35.36906, 35.51729, 35.66537, 35.81333, 35.96114, 
    36.10882, 36.25636, 36.40377, 36.55103, 36.69815, 36.84513, 36.99197, 
    37.13867, 37.28522, 37.43163, 37.5779, 37.72401, 37.86999, 38.01581, 
    38.16149, 38.30701, 38.45239, 38.59762, 38.74269, 38.88762, 39.03239, 
    39.17701, 39.32147, 39.46578, 39.60994, 39.75393, 39.89777, 40.04146, 
    40.18499, 40.32835, 40.47157, 40.61462, 40.7575, 40.90023, 41.0428, 
    41.1852, 41.32745, 41.46952, 41.61144, 41.75319, 41.89478, 42.03619, 
    42.17745, 42.31853, 42.45945, 42.6002, 42.74079, 42.88121, 43.02145, 
    43.16153, 43.30143, 43.44117, 43.58073, 43.72013,
  -19.93986, -19.81736, -19.69467, -19.57179, -19.44872, -19.32547, 
    -19.20203, -19.0784, -18.95458, -18.83057, -18.70638, -18.582, -18.45743, 
    -18.33267, -18.20773, -18.08259, -17.95727, -17.83176, -17.70606, 
    -17.58017, -17.4541, -17.32783, -17.20138, -17.07474, -16.94791, 
    -16.82089, -16.69369, -16.5663, -16.43871, -16.31094, -16.18299, 
    -16.05484, -15.9265, -15.79798, -15.66927, -15.54037, -15.41129, 
    -15.28201, -15.15255, -15.0229, -14.89307, -14.76305, -14.63283, 
    -14.50244, -14.37185, -14.24108, -14.11012, -13.97898, -13.84765, 
    -13.71613, -13.58442, -13.45253, -13.32046, -13.1882, -13.05575, 
    -12.92312, -12.7903, -12.6573, -12.52411, -12.39074, -12.25719, 
    -12.12345, -11.98952, -11.85542, -11.72113, -11.58665, -11.452, 
    -11.31716, -11.18214, -11.04693, -10.91155, -10.77598, -10.64023, 
    -10.50431, -10.3682, -10.23191, -10.09544, -9.958792, -9.821963, 
    -9.684957, -9.547771, -9.410408, -9.272866, -9.135148, -8.997252, 
    -8.859179, -8.72093, -8.582505, -8.443905, -8.305129, -8.166179, 
    -8.027055, -7.887756, -7.748284, -7.60864, -7.468822, -7.328834, 
    -7.188673, -7.048341, -6.907838, -6.767166, -6.626324, -6.485312, 
    -6.344133, -6.202785, -6.061269, -5.919587, -5.777738, -5.635724, 
    -5.493543, -5.351198, -5.208689, -5.066017, -4.923181, -4.780182, 
    -4.637022, -4.493701, -4.350219, -4.206577, -4.062776, -3.918816, 
    -3.774698, -3.630422, -3.48599, -3.341401, -3.196657, -3.051759, 
    -2.906706, -2.7615, -2.616142, -2.470631, -2.32497, -2.179158, -2.033196, 
    -1.887085, -1.740826, -1.594419, -1.447866, -1.301167, -1.154323, 
    -1.007334, -0.8602018, -0.7129268, -0.5655099, -0.4179518, -0.2702534, 
    -0.1224156, 0.02556087, 0.1736751, 0.3219263, 0.4703135, 0.6188359, 
    0.7674927, 0.9162828, 1.065206, 1.21426, 1.363445, 1.51276, 1.662204, 
    1.811776, 1.961475, 2.1113, 2.26125, 2.411324, 2.561522, 2.711841, 
    2.862283, 3.012844, 3.163525, 3.314324, 3.46524, 3.616273, 3.767421, 
    3.918684, 4.070059, 4.221547, 4.373147, 4.524856, 4.676674, 4.8286, 
    4.980634, 5.132772, 5.285017, 5.437364, 5.589815, 5.742366, 5.895019, 
    6.047771, 6.20062, 6.353567, 6.50661, 6.659748, 6.812979, 6.966303, 
    7.119719, 7.273224, 7.426818, 7.580501, 7.734271, 7.888125, 8.042065, 
    8.196087, 8.350191, 8.504377, 8.658642, 8.812985, 8.967405, 9.121902, 
    9.276474, 9.431118, 9.585835, 9.740623, 9.895482, 10.05041, 10.2054, 
    10.36046, 10.51559, 10.67078, 10.82603, 10.98134, 11.13671, 11.29214, 
    11.44763, 11.60317, 11.75877, 11.91442, 12.07012, 12.22588, 12.38168, 
    12.53753, 12.69343, 12.84938, 13.00536, 13.1614, 13.31747, 13.47358, 
    13.62973, 13.78592, 13.94215, 14.09841, 14.25471, 14.41103, 14.56739, 
    14.72378, 14.8802, 15.03664, 15.19311, 15.3496, 15.50612, 15.66266, 
    15.81921, 15.97579, 16.13239, 16.289, 16.44562, 16.60226, 16.75891, 
    16.91557, 17.07224, 17.22892, 17.38561, 17.5423, 17.699, 17.85569, 
    18.01239, 18.16909, 18.32579, 18.48248, 18.63918, 18.79586, 18.95254, 
    19.10921, 19.26587, 19.42252, 19.57915, 19.73578, 19.89239, 20.04898, 
    20.20555, 20.36211, 20.51864, 20.67515, 20.83164, 20.98811, 21.14455, 
    21.30096, 21.45734, 21.6137, 21.77002, 21.92631, 22.08256, 22.23878, 
    22.39497, 22.55112, 22.70722, 22.86329, 23.01931, 23.17529, 23.33123, 
    23.48712, 23.64297, 23.79876, 23.95451, 24.1102, 24.26585, 24.42144, 
    24.57697, 24.73245, 24.88787, 25.04323, 25.19854, 25.35378, 25.50896, 
    25.66407, 25.81912, 25.9741, 26.12902, 26.28387, 26.43864, 26.59335, 
    26.74798, 26.90254, 27.05703, 27.21144, 27.36577, 27.52002, 27.67419, 
    27.82828, 27.98229, 28.13622, 28.29006, 28.44382, 28.59748, 28.75106, 
    28.90456, 29.05796, 29.21127, 29.36448, 29.5176, 29.67063, 29.82356, 
    29.9764, 30.12914, 30.28177, 30.43431, 30.58674, 30.73907, 30.8913, 
    31.04342, 31.19544, 31.34735, 31.49915, 31.65084, 31.80242, 31.95389, 
    32.10525, 32.2565, 32.40763, 32.55864, 32.70954, 32.86032, 33.01098, 
    33.16152, 33.31194, 33.46225, 33.61242, 33.76248, 33.91241, 34.06221, 
    34.21189, 34.36144, 34.51087, 34.66016, 34.80933, 34.95836, 35.10726, 
    35.25603, 35.40467, 35.55317, 35.70153, 35.84976, 35.99786, 36.14581, 
    36.29362, 36.4413, 36.58884, 36.73623, 36.88348, 37.03059, 37.17756, 
    37.32438, 37.47106, 37.61759, 37.76397, 37.91021, 38.05629, 38.20223, 
    38.34802, 38.49366, 38.63914, 38.78448, 38.92966, 39.07469, 39.21956, 
    39.36428, 39.50885, 39.65326, 39.7975, 39.9416, 40.08553, 40.22931, 
    40.37292, 40.51638, 40.65968, 40.80281, 40.94579, 41.0886, 41.23124, 
    41.37373, 41.51604, 41.6582, 41.80019, 41.94201, 42.08367, 42.22515, 
    42.36648, 42.50763, 42.64861, 42.78943, 42.93008, 43.07055, 43.21085, 
    43.35099, 43.49095, 43.63074, 43.77036,
  -20.00684, -19.8842, -19.76137, -19.63835, -19.51515, -19.39176, -19.26818, 
    -19.1444, -19.02044, -18.8963, -18.77196, -18.64743, -18.52272, 
    -18.39782, -18.27272, -18.14744, -18.02197, -17.89631, -17.77046, 
    -17.64442, -17.51819, -17.39178, -17.26517, -17.13837, -17.01139, 
    -16.88421, -16.75685, -16.6293, -16.50156, -16.37362, -16.2455, -16.1172, 
    -15.9887, -15.86001, -15.73114, -15.60207, -15.47282, -15.34338, 
    -15.21375, -15.08393, -14.95392, -14.82372, -14.69334, -14.56277, 
    -14.43201, -14.30106, -14.16992, -14.0386, -13.90709, -13.77539, 
    -13.64351, -13.51144, -13.37918, -13.24673, -13.1141, -12.98128, 
    -12.84828, -12.71509, -12.58172, -12.44815, -12.31441, -12.18048, 
    -12.04636, -11.91206, -11.77757, -11.64291, -11.50805, -11.37302, 
    -11.2378, -11.10239, -10.96681, -10.83104, -10.69509, -10.55896, 
    -10.42264, -10.28615, -10.14947, -10.01262, -9.87558, -9.738363, 
    -9.600967, -9.463392, -9.325638, -9.187705, -9.049594, -8.911305, 
    -8.77284, -8.634196, -8.495378, -8.356381, -8.217211, -8.077864, 
    -7.938343, -7.798647, -7.658777, -7.518734, -7.378518, -7.238129, 
    -7.097568, -6.956835, -6.815932, -6.674858, -6.533613, -6.3922, 
    -6.250617, -6.108865, -5.966946, -5.824859, -5.682605, -5.540184, 
    -5.397599, -5.254848, -5.111932, -4.968852, -4.825608, -4.682202, 
    -4.538634, -4.394904, -4.251013, -4.106962, -3.962751, -3.818381, 
    -3.673852, -3.529166, -3.384323, -3.239324, -3.094168, -2.948858, 
    -2.803394, -2.657775, -2.512004, -2.366081, -2.220007, -2.073781, 
    -1.927406, -1.780882, -1.634209, -1.487389, -1.340422, -1.193308, 
    -1.04605, -0.8986469, -0.7511002, -0.6034106, -0.455579, -0.3076063, 
    -0.1594931, -0.01124041, 0.1371509, 0.2856801, 0.4343462, 0.5831484, 
    0.7320858, 0.8811574, 1.030362, 1.1797, 1.329169, 1.478769, 1.628499, 
    1.778357, 1.928343, 2.078457, 2.228696, 2.37906, 2.529548, 2.68016, 
    2.830893, 2.981748, 3.132722, 3.283816, 3.435028, 3.586357, 3.737803, 
    3.889363, 4.041037, 4.192824, 4.344723, 4.496733, 4.648853, 4.801082, 
    4.953418, 5.105861, 5.258409, 5.411062, 5.563818, 5.716676, 5.869636, 
    6.022695, 6.175853, 6.329109, 6.482462, 6.63591, 6.789453, 6.943089, 
    7.096816, 7.250635, 7.404543, 7.558539, 7.712624, 7.866794, 8.021049, 
    8.175388, 8.329809, 8.484312, 8.638896, 8.793558, 8.948298, 9.103114, 
    9.258005, 9.412971, 9.568009, 9.72312, 9.8783, 10.03355, 10.18887, 
    10.34425, 10.4997, 10.65521, 10.81079, 10.96642, 11.12212, 11.27788, 
    11.43369, 11.58956, 11.74549, 11.90147, 12.0575, 12.21358, 12.36971, 
    12.5259, 12.68212, 12.8384, 12.99472, 13.15108, 13.30748, 13.46393, 
    13.62041, 13.77693, 13.93349, 14.09008, 14.24671, 14.40337, 14.56006, 
    14.71678, 14.87353, 15.03031, 15.18711, 15.34394, 15.50079, 15.65766, 
    15.81455, 15.97146, 16.12839, 16.28534, 16.4423, 16.59927, 16.75626, 
    16.91325, 17.07026, 17.22728, 17.3843, 17.54132, 17.69835, 17.85539, 
    18.01242, 18.16945, 18.32649, 18.48352, 18.64054, 18.79756, 18.95458, 
    19.11158, 19.26858, 19.42556, 19.58253, 19.73949, 19.89643, 20.05336, 
    20.21027, 20.36716, 20.52402, 20.68087, 20.83769, 20.99449, 21.15126, 
    21.30801, 21.46473, 21.62141, 21.77807, 21.93469, 22.09128, 22.24783, 
    22.40434, 22.56082, 22.71726, 22.87366, 23.03001, 23.18633, 23.34259, 
    23.49881, 23.65499, 23.81111, 23.96719, 24.12321, 24.27918, 24.4351, 
    24.59096, 24.74676, 24.90251, 25.0582, 25.21383, 25.36939, 25.52489, 
    25.68033, 25.83571, 25.99101, 26.14625, 26.30142, 26.45652, 26.61155, 
    26.7665, 26.92138, 27.07619, 27.23091, 27.38556, 27.54013, 27.69462, 
    27.84903, 28.00336, 28.1576, 28.31176, 28.46583, 28.61981, 28.7737, 
    28.92751, 29.08122, 29.23484, 29.38837, 29.5418, 29.69514, 29.84838, 
    30.00152, 30.15457, 30.30751, 30.46035, 30.61309, 30.76573, 30.91826, 
    31.07069, 31.22301, 31.37522, 31.52732, 31.67931, 31.83119, 31.98296, 
    32.13462, 32.28616, 32.43759, 32.5889, 32.74009, 32.89117, 33.04212, 
    33.19296, 33.34367, 33.49427, 33.64473, 33.79508, 33.9453, 34.09539, 
    34.24536, 34.3952, 34.5449, 34.69448, 34.84393, 34.99325, 35.14243, 
    35.29148, 35.4404, 35.58918, 35.73782, 35.88633, 36.0347, 36.18293, 
    36.33102, 36.47897, 36.62678, 36.77445, 36.92197, 37.06936, 37.21659, 
    37.36368, 37.51062, 37.65742, 37.80407, 37.95057, 38.09692, 38.24312, 
    38.38918, 38.53507, 38.68082, 38.82641, 38.97186, 39.11714, 39.26227, 
    39.40725, 39.55206, 39.69672, 39.84123, 39.98557, 40.12976, 40.27378, 
    40.41765, 40.56136, 40.7049, 40.84828, 40.9915, 41.13455, 41.27744, 
    41.42017, 41.56273, 41.70512, 41.84735, 41.98941, 42.1313, 42.27303, 
    42.41458, 42.55597, 42.69719, 42.83823, 42.97911, 43.11982, 43.26035, 
    43.40071, 43.5409, 43.68091, 43.82076,
  -20.07399, -19.95122, -19.82825, -19.7051, -19.58175, -19.45822, -19.3345, 
    -19.21059, -19.08649, -18.9622, -18.83772, -18.71305, -18.58819, 
    -18.46314, -18.3379, -18.21247, -18.08685, -17.96104, -17.83504, 
    -17.70885, -17.58247, -17.4559, -17.32914, -17.20218, -17.07504, 
    -16.94771, -16.82019, -16.69248, -16.56458, -16.43649, -16.3082, 
    -16.17973, -16.05107, -15.92222, -15.79318, -15.66395, -15.53453, 
    -15.40492, -15.27512, -15.14513, -15.01495, -14.88458, -14.75402, 
    -14.62328, -14.49234, -14.36122, -14.22991, -14.09841, -13.96672, 
    -13.83484, -13.70277, -13.57052, -13.43808, -13.30545, -13.17263, 
    -13.03963, -12.90644, -12.77306, -12.63949, -12.50574, -12.37181, 
    -12.23768, -12.10337, -11.96888, -11.8342, -11.69933, -11.56428, 
    -11.42905, -11.29363, -11.15803, -11.02224, -10.88627, -10.75012, 
    -10.61378, -10.47726, -10.34056, -10.20368, -10.06662, -9.929369, 
    -9.791942, -9.654335, -9.516547, -9.378579, -9.240433, -9.102106, 
    -8.963601, -8.824918, -8.686057, -8.547018, -8.407803, -8.26841, 
    -8.12884, -7.989096, -7.849176, -7.709081, -7.568811, -7.428367, 
    -7.28775, -7.14696, -7.005997, -6.864861, -6.723555, -6.582077, 
    -6.440429, -6.29861, -6.156622, -6.014465, -5.872139, -5.729646, 
    -5.586985, -5.444158, -5.301164, -5.158004, -5.01468, -4.871191, 
    -4.727538, -4.583722, -4.439744, -4.295603, -4.151301, -4.006839, 
    -3.862216, -3.717435, -3.572494, -3.427395, -3.282139, -3.136727, 
    -2.991158, -2.845434, -2.699556, -2.553524, -2.407338, -2.261001, 
    -2.114511, -1.967871, -1.821081, -1.674141, -1.527053, -1.379817, 
    -1.232434, -1.084905, -0.9372303, -0.7894111, -0.6414481, -0.4933422, 
    -0.3450942, -0.1967049, -0.04817522, 0.100494, 0.249302, 0.3982478, 
    0.5473306, 0.6965494, 0.8459034, 0.9953917, 1.145013, 1.294767, 1.444653, 
    1.594669, 1.744815, 1.89509, 2.045492, 2.196021, 2.346677, 2.497456, 
    2.64836, 2.799387, 2.950536, 3.101805, 3.253195, 3.404703, 3.556329, 
    3.708073, 3.859932, 4.011905, 4.163993, 4.316193, 4.468505, 4.620927, 
    4.773459, 4.926099, 5.078847, 5.2317, 5.384659, 5.537723, 5.690888, 
    5.844156, 5.997524, 6.150992, 6.304558, 6.458222, 6.611982, 6.765836, 
    6.919785, 7.073826, 7.227959, 7.382182, 7.536493, 7.690894, 7.84538, 
    7.999952, 8.154609, 8.309349, 8.46417, 8.619073, 8.774055, 8.929115, 
    9.084252, 9.239466, 9.394753, 9.550115, 9.705547, 9.861051, 10.01662, 
    10.17227, 10.32797, 10.48375, 10.63959, 10.79549, 10.95145, 11.10748, 
    11.26356, 11.4197, 11.5759, 11.73216, 11.88847, 12.04483, 12.20124, 
    12.3577, 12.51421, 12.67077, 12.82738, 12.98403, 13.14072, 13.29746, 
    13.45423, 13.61105, 13.76791, 13.9248, 14.08172, 14.23868, 14.39568, 
    14.5527, 14.70976, 14.86684, 15.02395, 15.18109, 15.33825, 15.49544, 
    15.65265, 15.80987, 15.96712, 16.12438, 16.28167, 16.43896, 16.59627, 
    16.75359, 16.91093, 17.06827, 17.22562, 17.38298, 17.54034, 17.69771, 
    17.85508, 18.01245, 18.16982, 18.32719, 18.48455, 18.64191, 18.79927, 
    18.95662, 19.11396, 19.27129, 19.42861, 19.58592, 19.74322, 19.90049, 
    20.05776, 20.215, 20.37222, 20.52943, 20.68661, 20.84377, 21.0009, 
    21.15801, 21.31509, 21.47214, 21.62916, 21.78615, 21.9431, 22.10002, 
    22.25691, 22.41376, 22.57057, 22.72734, 22.88407, 23.04075, 23.1974, 
    23.354, 23.51055, 23.66705, 23.82351, 23.97991, 24.13626, 24.29256, 
    24.44881, 24.605, 24.76113, 24.91721, 25.07322, 25.22918, 25.38507, 
    25.5409, 25.69666, 25.85236, 26.00799, 26.16355, 26.31904, 26.47447, 
    26.62982, 26.78509, 26.94029, 27.09542, 27.25047, 27.40544, 27.56033, 
    27.71513, 27.86986, 28.0245, 28.17906, 28.33354, 28.48792, 28.64222, 
    28.79643, 28.95055, 29.10457, 29.25851, 29.41235, 29.56609, 29.71974, 
    29.87329, 30.02674, 30.1801, 30.33335, 30.4865, 30.63954, 30.79249, 
    30.94532, 31.09805, 31.25068, 31.40319, 31.5556, 31.70789, 31.86007, 
    32.01214, 32.1641, 32.31594, 32.46766, 32.61927, 32.77076, 32.92213, 
    33.07338, 33.22451, 33.37552, 33.5264, 33.67716, 33.8278, 33.97831, 
    34.12869, 34.27895, 34.42907, 34.57906, 34.72893, 34.87866, 35.02826, 
    35.17773, 35.32706, 35.47626, 35.62532, 35.77425, 35.92303, 36.07168, 
    36.22019, 36.36855, 36.51678, 36.66486, 36.81281, 36.9606, 37.10825, 
    37.25576, 37.40312, 37.55033, 37.6974, 37.84431, 37.99108, 38.1377, 
    38.28416, 38.43047, 38.57663, 38.72264, 38.8685, 39.01419, 39.15974, 
    39.30513, 39.45036, 39.59543, 39.74035, 39.88511, 40.0297, 40.17414, 
    40.31842, 40.46253, 40.60648, 40.75027, 40.8939, 41.03736, 41.18066, 
    41.3238, 41.46676, 41.60956, 41.7522, 41.89466, 42.03696, 42.17909, 
    42.32106, 42.46284, 42.60447, 42.74592, 42.8872, 43.02831, 43.16924, 
    43.31001, 43.4506, 43.59101, 43.73125, 43.87132,
  -20.14132, -20.01841, -19.89531, -19.77202, -19.64854, -19.52487, 
    -19.40101, -19.27696, -19.15271, -19.02828, -18.90366, -18.77884, 
    -18.65384, -18.52864, -18.40326, -18.27768, -18.15191, -18.02595, 
    -17.8998, -17.77346, -17.64692, -17.5202, -17.39329, -17.26618, 
    -17.13888, -17.01139, -16.88371, -16.75584, -16.62778, -16.49953, 
    -16.37109, -16.24245, -16.11363, -15.98461, -15.8554, -15.72601, 
    -15.59642, -15.46664, -15.33667, -15.20651, -15.07616, -14.94562, 
    -14.81489, -14.68397, -14.55286, -14.42156, -14.29007, -14.15839, 
    -14.02652, -13.89446, -13.76222, -13.62978, -13.49716, -13.36434, 
    -13.23134, -13.09815, -12.96477, -12.83121, -12.69745, -12.56351, 
    -12.42938, -12.29507, -12.16057, -12.02588, -11.891, -11.75594, 
    -11.62069, -11.48526, -11.34964, -11.21384, -11.07785, -10.94168, 
    -10.80532, -10.66878, -10.53206, -10.39515, -10.25806, -10.12079, 
    -9.983331, -9.845694, -9.707874, -9.569875, -9.431693, -9.293332, 
    -9.15479, -9.016068, -8.877168, -8.738088, -8.598829, -8.459393, 
    -8.319778, -8.179987, -8.040018, -7.899873, -7.759552, -7.619055, 
    -7.478384, -7.337537, -7.196517, -7.055323, -6.913956, -6.772416, 
    -6.630704, -6.488821, -6.346766, -6.204541, -6.062146, -5.919581, 
    -5.776848, -5.633946, -5.490876, -5.347639, -5.204236, -5.060666, 
    -4.916931, -4.773031, -4.628967, -4.484739, -4.340349, -4.195796, 
    -4.051081, -3.906205, -3.761169, -3.615974, -3.470619, -3.325106, 
    -3.179435, -3.033608, -2.887624, -2.741485, -2.59519, -2.448742, 
    -2.302141, -2.155386, -2.008481, -1.861424, -1.714216, -1.566859, 
    -1.419354, -1.271701, -1.1239, -0.975953, -0.8278605, -0.6796234, 
    -0.5312424, -0.3827183, -0.2340521, -0.08524454, 0.06370348, 0.2127911, 
    0.3620175, 0.5113816, 0.6608828, 0.81052, 0.9602923, 1.110199, 1.260239, 
    1.410411, 1.560715, 1.711149, 1.861713, 2.012406, 2.163226, 2.314173, 
    2.465245, 2.616442, 2.767763, 2.919207, 3.070772, 3.222459, 3.374264, 
    3.526189, 3.678231, 3.83039, 3.982664, 4.135053, 4.287555, 4.44017, 
    4.592896, 4.745732, 4.898677, 5.05173, 5.204891, 5.358157, 5.511528, 
    5.665002, 5.818579, 5.972257, 6.126036, 6.279913, 6.433889, 6.587961, 
    6.742129, 6.896392, 7.050747, 7.205195, 7.359734, 7.514362, 7.66908, 
    7.823884, 7.978775, 8.13375, 8.288809, 8.443951, 8.599174, 8.754477, 
    8.909859, 9.065318, 9.220854, 9.376465, 9.532149, 9.687906, 9.843735, 
    9.999634, 10.1556, 10.31164, 10.46774, 10.6239, 10.78013, 10.93642, 
    11.09278, 11.24919, 11.40566, 11.56219, 11.71877, 11.87541, 12.0321, 
    12.18885, 12.34564, 12.50248, 12.65938, 12.81631, 12.9733, 13.13032, 
    13.28739, 13.4445, 13.60165, 13.75884, 13.91607, 14.07333, 14.23063, 
    14.38795, 14.54531, 14.70271, 14.86012, 15.01757, 15.17505, 15.33254, 
    15.49007, 15.64761, 15.80517, 15.96276, 16.12036, 16.27798, 16.43561, 
    16.59326, 16.75092, 16.90859, 17.06627, 17.22396, 17.38165, 17.53935, 
    17.69706, 17.85476, 18.01247, 18.17018, 18.32789, 18.48559, 18.64329, 
    18.80099, 18.95868, 19.11635, 19.27402, 19.43168, 19.58932, 19.74696, 
    19.90457, 20.06217, 20.21975, 20.37731, 20.53485, 20.69237, 20.84986, 
    21.00734, 21.16478, 21.32219, 21.47958, 21.63694, 21.79426, 21.95155, 
    22.10881, 22.26603, 22.42321, 22.58035, 22.73746, 22.89452, 23.05154, 
    23.20852, 23.36545, 23.52233, 23.67916, 23.83595, 23.99269, 24.14937, 
    24.306, 24.46257, 24.61909, 24.77556, 24.93196, 25.0883, 25.24459, 
    25.4008, 25.55696, 25.71305, 25.86908, 26.02503, 26.18092, 26.33674, 
    26.49248, 26.64816, 26.80375, 26.95928, 27.11473, 27.27009, 27.42538, 
    27.5806, 27.73572, 27.89077, 28.04573, 28.20061, 28.3554, 28.5101, 
    28.66472, 28.81924, 28.97367, 29.12802, 29.28226, 29.43642, 29.59047, 
    29.74443, 29.8983, 30.05206, 30.20572, 30.35928, 30.51274, 30.66609, 
    30.81934, 30.97249, 31.12552, 31.27845, 31.43127, 31.58398, 31.73658, 
    31.88906, 32.04143, 32.19369, 32.34583, 32.49785, 32.64976, 32.80154, 
    32.95321, 33.10476, 33.25618, 33.40748, 33.55866, 33.70971, 33.86064, 
    34.01144, 34.16211, 34.31266, 34.46307, 34.61335, 34.7635, 34.91352, 
    35.06341, 35.21316, 35.36277, 35.51225, 35.6616, 35.8108, 35.95987, 
    36.10879, 36.25758, 36.40622, 36.55472, 36.70308, 36.8513, 36.99937, 
    37.14729, 37.29507, 37.4427, 37.59018, 37.73751, 37.8847, 38.03173, 
    38.17861, 38.32534, 38.47192, 38.61834, 38.76461, 38.91073, 39.05669, 
    39.20249, 39.34813, 39.49362, 39.63895, 39.78412, 39.92913, 40.07398, 
    40.21867, 40.3632, 40.50756, 40.65177, 40.7958, 40.93968, 41.08339, 
    41.22693, 41.37031, 41.51352, 41.65656, 41.79944, 41.94214, 42.08468, 
    42.22705, 42.36925, 42.51128, 42.65313, 42.79482, 42.93633, 43.07767, 
    43.21884, 43.35983, 43.50065, 43.64129, 43.78176, 43.92205,
  -20.20883, -20.08579, -19.96255, -19.83912, -19.71551, -19.5917, -19.4677, 
    -19.3435, -19.21912, -19.09455, -18.96978, -18.84482, -18.71967, 
    -18.59433, -18.46879, -18.34307, -18.21715, -18.09104, -17.96474, 
    -17.83825, -17.71156, -17.58468, -17.45761, -17.33035, -17.2029, 
    -17.07526, -16.94742, -16.81939, -16.69117, -16.56276, -16.43415, 
    -16.30535, -16.17636, -16.04718, -15.91781, -15.78825, -15.65849, 
    -15.52854, -15.3984, -15.26807, -15.13755, -15.00684, -14.87594, 
    -14.74484, -14.61356, -14.48208, -14.35041, -14.21856, -14.08651, 
    -13.95427, -13.82184, -13.68922, -13.55641, -13.42342, -13.29023, 
    -13.15685, -13.02329, -12.88953, -12.75559, -12.62146, -12.48714, 
    -12.35263, -12.21794, -12.08305, -11.94798, -11.81272, -11.67728, 
    -11.54165, -11.40583, -11.26983, -11.13364, -10.99726, -10.8607, 
    -10.72396, -10.58703, -10.44991, -10.31261, -10.17513, -10.03747, 
    -9.899619, -9.761589, -9.623376, -9.484981, -9.346404, -9.207646, 
    -9.068707, -8.929589, -8.79029, -8.650811, -8.511153, -8.371317, 
    -8.231302, -8.091109, -7.950739, -7.810192, -7.669468, -7.528568, 
    -7.387492, -7.246242, -7.104816, -6.963216, -6.821443, -6.679497, 
    -6.537378, -6.395087, -6.252624, -6.10999, -5.967186, -5.824212, 
    -5.681068, -5.537755, -5.394275, -5.250627, -5.106812, -4.96283, 
    -4.818682, -4.674369, -4.529891, -4.38525, -4.240446, -4.095478, 
    -3.950349, -3.805058, -3.659607, -3.513995, -3.368224, -3.222295, 
    -3.076208, -2.929963, -2.783562, -2.637006, -2.490294, -2.343428, 
    -2.196408, -2.049236, -1.901911, -1.754436, -1.606809, -1.459033, 
    -1.311109, -1.163036, -1.014816, -0.8664495, -0.7179374, -0.5692804, 
    -0.4204796, -0.2715356, -0.1224494, 0.02677824, 0.1761463, 0.3256541, 
    0.4753006, 0.6250849, 0.7750062, 0.9250635, 1.075256, 1.225582, 1.376042, 
    1.526635, 1.677358, 1.828212, 1.979196, 2.130308, 2.281547, 2.432913, 
    2.584405, 2.736021, 2.887761, 3.039623, 3.191607, 3.343711, 3.495935, 
    3.648277, 3.800736, 3.953312, 4.106003, 4.258809, 4.411727, 4.564758, 
    4.717899, 4.87115, 5.024511, 5.177979, 5.331553, 5.485233, 5.639017, 
    5.792904, 5.946894, 6.100984, 6.255174, 6.409462, 6.563848, 6.718331, 
    6.872909, 7.02758, 7.182344, 7.3372, 7.492146, 7.647182, 7.802304, 
    7.957514, 8.11281, 8.268189, 8.423653, 8.579197, 8.734822, 8.890527, 
    9.04631, 9.202169, 9.358105, 9.514114, 9.670197, 9.826351, 9.982576, 
    10.13887, 10.29523, 10.45166, 10.60816, 10.76471, 10.92134, 11.07802, 
    11.23476, 11.39156, 11.54842, 11.70534, 11.86231, 12.01933, 12.17641, 
    12.33353, 12.49071, 12.64793, 12.80521, 12.96252, 13.11988, 13.27729, 
    13.43473, 13.59222, 13.74974, 13.9073, 14.0649, 14.22253, 14.3802, 
    14.5379, 14.69562, 14.85338, 15.01117, 15.16898, 15.32681, 15.48467, 
    15.64255, 15.80046, 15.95838, 16.11632, 16.27427, 16.43225, 16.59023, 
    16.74823, 16.90624, 17.06426, 17.22229, 17.38032, 17.53836, 17.69641, 
    17.85445, 18.0125, 18.17055, 18.32859, 18.48664, 18.64468, 18.80271, 
    18.96074, 19.11875, 19.27676, 19.43476, 19.59274, 19.75071, 19.90867, 
    20.0666, 20.22452, 20.38242, 20.5403, 20.69816, 20.85599, 21.0138, 
    21.17158, 21.32933, 21.48705, 21.64474, 21.8024, 21.96003, 22.11762, 
    22.27518, 22.4327, 22.59018, 22.74761, 22.90501, 23.06237, 23.21968, 
    23.37694, 23.53416, 23.69133, 23.84844, 24.00551, 24.16253, 24.31949, 
    24.47639, 24.63325, 24.79004, 24.94677, 25.10344, 25.26006, 25.4166, 
    25.57309, 25.72951, 25.88586, 26.04214, 26.19835, 26.3545, 26.51057, 
    26.66657, 26.82249, 26.97834, 27.13411, 27.2898, 27.44541, 27.60094, 
    27.7564, 27.91176, 28.06704, 28.22224, 28.37735, 28.53237, 28.6873, 
    28.84214, 28.99689, 29.15155, 29.30611, 29.46058, 29.61495, 29.76922, 
    29.9234, 30.07747, 30.23145, 30.38532, 30.53908, 30.69275, 30.8463, 
    30.99976, 31.1531, 31.30633, 31.45946, 31.61247, 31.76537, 31.91816, 
    32.07083, 32.22339, 32.37583, 32.52815, 32.68036, 32.83244, 32.98441, 
    33.13625, 33.28797, 33.43957, 33.59104, 33.74239, 33.8936, 34.0447, 
    34.19566, 34.34649, 34.4972, 34.64777, 34.79821, 34.94851, 35.09868, 
    35.24872, 35.39862, 35.54838, 35.69801, 35.84749, 35.99684, 36.14604, 
    36.2951, 36.44403, 36.5928, 36.74144, 36.88993, 37.03827, 37.18647, 
    37.33452, 37.48242, 37.63017, 37.77777, 37.92522, 38.07253, 38.21967, 
    38.36667, 38.51351, 38.6602, 38.80673, 38.95311, 39.09933, 39.24539, 
    39.39129, 39.53704, 39.68262, 39.82805, 39.97332, 40.11842, 40.26336, 
    40.40814, 40.55276, 40.69721, 40.8415, 40.98561, 41.12957, 41.27336, 
    41.41698, 41.56044, 41.70372, 41.84684, 41.98979, 42.13256, 42.27517, 
    42.41761, 42.55987, 42.70196, 42.84388, 42.98563, 43.1272, 43.2686, 
    43.40982, 43.55087, 43.69174, 43.83244, 43.97295,
  -20.27653, -20.15335, -20.02998, -19.90641, -19.78266, -19.65871, 
    -19.53457, -19.41023, -19.28571, -19.16099, -19.03608, -18.91098, 
    -18.78568, -18.6602, -18.53452, -18.40864, -18.28258, -18.15632, 
    -18.02987, -17.90322, -17.77638, -17.64935, -17.52213, -17.39471, 
    -17.2671, -17.1393, -17.01131, -16.88312, -16.75474, -16.62616, -16.4974, 
    -16.36844, -16.23928, -16.10994, -15.9804, -15.85067, -15.72075, 
    -15.59063, -15.46032, -15.32982, -15.19913, -15.06824, -14.93717, 
    -14.8059, -14.67444, -14.54278, -14.41094, -14.2789, -14.14668, 
    -14.01426, -13.88165, -13.74885, -13.61585, -13.48267, -13.3493, 
    -13.21574, -13.08198, -12.94804, -12.81391, -12.67959, -12.54508, 
    -12.41037, -12.27549, -12.14041, -12.00514, -11.86969, -11.73404, 
    -11.59821, -11.4622, -11.32599, -11.1896, -11.05302, -10.91626, 
    -10.77931, -10.64217, -10.50485, -10.36735, -10.22966, -10.09178, 
    -9.953721, -9.815477, -9.677052, -9.538443, -9.399651, -9.260676, 
    -9.12152, -8.982183, -8.842665, -8.702966, -8.563087, -8.423027, 
    -8.282788, -8.142371, -8.001776, -7.861001, -7.72005, -7.578921, 
    -7.437615, -7.296134, -7.154477, -7.012644, -6.870637, -6.728456, 
    -6.5861, -6.443572, -6.300871, -6.157999, -6.014954, -5.871738, 
    -5.728353, -5.584797, -5.441072, -5.297179, -5.153117, -5.008888, 
    -4.864492, -4.71993, -4.575202, -4.430309, -4.285252, -4.140031, 
    -3.994648, -3.849102, -3.703394, -3.557525, -3.411496, -3.265307, 
    -3.118959, -2.972454, -2.82579, -2.67897, -2.531994, -2.384863, 
    -2.237577, -2.090137, -1.942545, -1.7948, -1.646904, -1.498857, -1.35066, 
    -1.202314, -1.05382, -0.905179, -0.756391, -0.6074574, -0.4583789, 
    -0.3091564, -0.1597907, -0.01028264, 0.1393668, 0.2891568, 0.4390864, 
    0.5891547, 0.7393609, 0.8897041, 1.040183, 1.190797, 1.341546, 1.492427, 
    1.643441, 1.794586, 1.945862, 2.097266, 2.2488, 2.40046, 2.552247, 
    2.704159, 2.856196, 3.008356, 3.160638, 3.313042, 3.465566, 3.618209, 
    3.77097, 3.923849, 4.076843, 4.229953, 4.383176, 4.536512, 4.68996, 
    4.843519, 4.997187, 5.150963, 5.304847, 5.458837, 5.612932, 5.76713, 
    5.921432, 6.075835, 6.230339, 6.384942, 6.539643, 6.694441, 6.849335, 
    7.004323, 7.159404, 7.314579, 7.469843, 7.625198, 7.780641, 7.936172, 
    8.091788, 8.24749, 8.403275, 8.559142, 8.715092, 8.87112, 9.027227, 
    9.183413, 9.339673, 9.496009, 9.652418, 9.8089, 9.965452, 10.12208, 
    10.27877, 10.43552, 10.59235, 10.74924, 10.90619, 11.0632, 11.22027, 
    11.37741, 11.5346, 11.69185, 11.84915, 12.00651, 12.16392, 12.32138, 
    12.47889, 12.63645, 12.79405, 12.95171, 13.1094, 13.26714, 13.42492, 
    13.58275, 13.74061, 13.89851, 14.05644, 14.21441, 14.37241, 14.53045, 
    14.68851, 14.84661, 15.00473, 15.16288, 15.32106, 15.47926, 15.63748, 
    15.79572, 15.95398, 16.11226, 16.27056, 16.42887, 16.5872, 16.74553, 
    16.90388, 17.06224, 17.22061, 17.37899, 17.53737, 17.69575, 17.85414, 
    18.01253, 18.17092, 18.3293, 18.48769, 18.64606, 18.80444, 18.96281, 
    19.12116, 19.27951, 19.43785, 19.59617, 19.75448, 19.91278, 20.07105, 
    20.22931, 20.38755, 20.54577, 20.70396, 20.86213, 21.02028, 21.1784, 
    21.33649, 21.49455, 21.65258, 21.81058, 21.96854, 22.12647, 22.28437, 
    22.44222, 22.60004, 22.75781, 22.91555, 23.07323, 23.23088, 23.38848, 
    23.54603, 23.70354, 23.86099, 24.01839, 24.17574, 24.33303, 24.49027, 
    24.64745, 24.80458, 24.96164, 25.11864, 25.27559, 25.43246, 25.58928, 
    25.74603, 25.9027, 26.05932, 26.21586, 26.37233, 26.52873, 26.68505, 
    26.8413, 26.99747, 27.15357, 27.30958, 27.46552, 27.62137, 27.77715, 
    27.93283, 28.08844, 28.24395, 28.39938, 28.55472, 28.70997, 28.86513, 
    29.0202, 29.17517, 29.33005, 29.48483, 29.63952, 29.79411, 29.9486, 
    30.10298, 30.25727, 30.41145, 30.56553, 30.7195, 30.87337, 31.02713, 
    31.18078, 31.33432, 31.48775, 31.64107, 31.79427, 31.94736, 32.10034, 
    32.2532, 32.40594, 32.55857, 32.71107, 32.86346, 33.01572, 33.16786, 
    33.31988, 33.47177, 33.62354, 33.77518, 33.92669, 34.07808, 34.22933, 
    34.38046, 34.53145, 34.68231, 34.83303, 34.98363, 35.13409, 35.28441, 
    35.43459, 35.58464, 35.73455, 35.88432, 36.03394, 36.18343, 36.33277, 
    36.48197, 36.63103, 36.77994, 36.9287, 37.07732, 37.22579, 37.37411, 
    37.52229, 37.67031, 37.81818, 37.9659, 38.11347, 38.26089, 38.40815, 
    38.55525, 38.70221, 38.849, 38.99564, 39.14212, 39.28844, 39.4346, 
    39.58061, 39.72645, 39.87214, 40.01765, 40.16301, 40.30821, 40.45324, 
    40.59811, 40.74281, 40.88734, 41.03172, 41.17591, 41.31995, 41.46382, 
    41.60752, 41.75105, 41.89441, 42.03759, 42.18061, 42.32346, 42.46613, 
    42.60863, 42.75096, 42.89311, 43.03509, 43.1769, 43.31853, 43.45998, 
    43.60126, 43.74236, 43.88328, 44.02403,
  -20.3444, -20.22109, -20.09758, -19.97388, -19.84999, -19.7259, -19.60162, 
    -19.47715, -19.35248, -19.22762, -19.10257, -18.97732, -18.85188, 
    -18.72625, -18.60042, -18.4744, -18.34819, -18.22178, -18.09517, 
    -17.96838, -17.84139, -17.71421, -17.58683, -17.45926, -17.33149, 
    -17.20353, -17.07538, -16.94703, -16.81849, -16.68976, -16.56083, 
    -16.4317, -16.30239, -16.17288, -16.04317, -15.91328, -15.78319, 
    -15.6529, -15.52242, -15.39175, -15.26089, -15.12983, -14.99858, 
    -14.86714, -14.7355, -14.60367, -14.47165, -14.33943, -14.20703, 
    -14.07443, -13.94164, -13.80865, -13.67548, -13.54211, -13.40855, 
    -13.2748, -13.14086, -13.00673, -12.87241, -12.7379, -12.60319, -12.4683, 
    -12.33322, -12.19794, -12.06248, -11.92683, -11.79099, -11.65496, 
    -11.51874, -11.38234, -11.24574, -11.10896, -10.972, -10.83484, -10.6975, 
    -10.55997, -10.42225, -10.28436, -10.14627, -10.008, -9.869543, 
    -9.730904, -9.592079, -9.453072, -9.313881, -9.174507, -9.034951, 
    -8.895213, -8.755293, -8.615192, -8.47491, -8.334448, -8.193805, 
    -8.052983, -7.911982, -7.770802, -7.629444, -7.487908, -7.346195, 
    -7.204306, -7.06224, -6.919998, -6.777581, -6.63499, -6.492224, 
    -6.349284, -6.206172, -6.062887, -5.91943, -5.775801, -5.632001, 
    -5.488032, -5.343893, -5.199584, -5.055107, -4.910462, -4.76565, 
    -4.620671, -4.475527, -4.330217, -4.184742, -4.039103, -3.893301, 
    -3.747336, -3.601209, -3.454921, -3.308472, -3.161864, -3.015096, 
    -2.868169, -2.721085, -2.573844, -2.426447, -2.278894, -2.131186, 
    -1.983325, -1.83531, -1.687143, -1.538825, -1.390355, -1.241736, 
    -1.092967, -0.94405, -0.7949855, -0.6457744, -0.4964174, -0.3469155, 
    -0.1972694, -0.04748015, 0.1024515, 0.2525245, 0.4027381, 0.5530914, 
    0.7035834, 0.8542133, 1.00498, 1.155883, 1.306921, 1.458092, 1.609397, 
    1.760834, 1.912403, 2.064101, 2.215929, 2.367885, 2.519968, 2.672177, 
    2.824512, 2.976971, 3.129553, 3.282257, 3.435082, 3.588027, 3.741091, 
    3.894273, 4.047572, 4.200987, 4.354516, 4.508159, 4.661914, 4.815781, 
    4.969758, 5.123844, 5.278039, 5.432339, 5.586746, 5.741258, 5.895873, 
    6.05059, 6.205408, 6.360326, 6.515343, 6.670458, 6.825669, 6.980975, 
    7.136375, 7.291869, 7.447453, 7.603128, 7.758893, 7.914745, 8.070684, 
    8.226708, 8.382817, 8.539009, 8.695283, 8.851637, 9.00807, 9.164581, 
    9.321169, 9.477832, 9.634569, 9.791379, 9.94826, 10.10521, 10.26223, 
    10.41932, 10.57648, 10.7337, 10.89098, 11.04832, 11.20573, 11.3632, 
    11.52072, 11.6783, 11.83594, 11.99363, 12.15138, 12.30917, 12.46702, 
    12.62491, 12.78286, 12.94085, 13.09888, 13.25696, 13.41508, 13.57324, 
    13.73143, 13.88967, 14.04795, 14.20625, 14.3646, 14.52297, 14.68138, 
    14.83981, 14.99828, 15.15677, 15.31528, 15.47382, 15.63238, 15.79097, 
    15.94957, 16.10819, 16.26683, 16.42548, 16.58415, 16.74283, 16.90152, 
    17.06022, 17.21893, 17.37765, 17.53637, 17.6951, 17.85382, 18.01255, 
    18.17128, 18.33001, 18.48874, 18.64746, 18.80618, 18.96488, 19.12358, 
    19.28227, 19.44095, 19.59962, 19.75827, 19.9169, 20.07552, 20.23412, 
    20.3927, 20.55126, 20.70979, 20.86831, 21.02679, 21.18525, 21.34368, 
    21.50208, 21.66045, 21.81879, 21.97709, 22.13536, 22.29359, 22.45179, 
    22.60994, 22.76805, 22.92612, 23.08415, 23.24213, 23.40007, 23.55795, 
    23.71579, 23.87358, 24.03132, 24.189, 24.34663, 24.5042, 24.66172, 
    24.81917, 24.97657, 25.13391, 25.29118, 25.44839, 25.60553, 25.76261, 
    25.91962, 26.07656, 26.23343, 26.39023, 26.54696, 26.70361, 26.86018, 
    27.01668, 27.1731, 27.32944, 27.4857, 27.64188, 27.79798, 27.95399, 
    28.10991, 28.26575, 28.4215, 28.57716, 28.73273, 28.88821, 29.0436, 
    29.19889, 29.35409, 29.50918, 29.66419, 29.81909, 29.97389, 30.12859, 
    30.28319, 30.43769, 30.59208, 30.74636, 30.90054, 31.05461, 31.20856, 
    31.36242, 31.51615, 31.66978, 31.82329, 31.97668, 32.12997, 32.28313, 
    32.43617, 32.5891, 32.74191, 32.89459, 33.04715, 33.19959, 33.35191, 
    33.5041, 33.65616, 33.8081, 33.9599, 34.11158, 34.26313, 34.41455, 
    34.56583, 34.71698, 34.868, 35.01888, 35.16962, 35.32023, 35.4707, 
    35.62103, 35.77122, 35.92128, 36.07118, 36.22095, 36.37057, 36.52005, 
    36.66939, 36.81858, 36.96762, 37.11651, 37.26525, 37.41385, 37.5623, 
    37.71059, 37.85873, 38.00673, 38.15456, 38.30225, 38.44977, 38.59715, 
    38.74436, 38.89142, 39.03832, 39.18507, 39.33165, 39.47807, 39.62434, 
    39.77044, 39.91637, 40.06215, 40.20776, 40.35321, 40.4985, 40.64362, 
    40.78857, 40.93335, 41.07797, 41.22242, 41.3667, 41.51082, 41.65476, 
    41.79853, 41.94213, 42.08556, 42.22882, 42.37191, 42.51482, 42.65756, 
    42.80012, 42.94251, 43.08472, 43.22676, 43.36863, 43.51031, 43.65182, 
    43.79315, 43.9343, 44.07527,
  -20.41247, -20.28901, -20.16537, -20.04153, -19.9175, -19.79328, -19.66886, 
    -19.54424, -19.41944, -19.29444, -19.16924, -19.04385, -18.91826, 
    -18.79248, -18.66651, -18.54034, -18.41398, -18.28742, -18.16067, 
    -18.03372, -17.90658, -17.77924, -17.65171, -17.52398, -17.39606, 
    -17.26795, -17.13964, -17.01113, -16.88243, -16.75353, -16.62444, 
    -16.49516, -16.36568, -16.236, -16.10613, -15.97607, -15.84581, 
    -15.71536, -15.58471, -15.45387, -15.32283, -15.1916, -15.06018, 
    -14.92856, -14.79675, -14.66474, -14.53254, -14.40015, -14.26756, 
    -14.13478, -14.00181, -13.86864, -13.73528, -13.60173, -13.46799, 
    -13.33405, -13.19992, -13.0656, -12.93109, -12.79639, -12.66149, 
    -12.52641, -12.39113, -12.25566, -12.12, -11.98415, -11.84812, -11.71189, 
    -11.57547, -11.43886, -11.30207, -11.16508, -11.02791, -10.89055, 
    -10.753, -10.61527, -10.47734, -10.33923, -10.20094, -10.06245, 
    -9.923785, -9.784932, -9.645893, -9.50667, -9.367262, -9.227671, 
    -9.087895, -8.947937, -8.807796, -8.667472, -8.526967, -8.38628, 
    -8.245412, -8.104363, -7.963134, -7.821726, -7.680139, -7.538372, 
    -7.396427, -7.254305, -7.112005, -6.969528, -6.826876, -6.684047, 
    -6.541043, -6.397864, -6.254512, -6.110985, -5.967286, -5.823414, 
    -5.67937, -5.535155, -5.390769, -5.246214, -5.101488, -4.956594, 
    -4.811532, -4.666301, -4.520904, -4.37534, -4.229611, -4.083716, 
    -3.937657, -3.791435, -3.645049, -3.498502, -3.351792, -3.204922, 
    -3.057891, -2.910701, -2.763352, -2.615845, -2.468181, -2.320361, 
    -2.172385, -2.024253, -1.875968, -1.727529, -1.578938, -1.430195, 
    -1.281301, -1.132257, -0.9830636, -0.8337218, -0.6842323, -0.534596, 
    -0.3848138, -0.2348867, -0.08481531, 0.06539932, 0.2157563, 0.3662548, 
    0.5168939, 0.6676726, 0.81859, 0.9696453, 1.120837, 1.272165, 1.423628, 
    1.575225, 1.726956, 1.878818, 2.030811, 2.182934, 2.335186, 2.487567, 
    2.640074, 2.792708, 2.945466, 3.098349, 3.251354, 3.404482, 3.55773, 
    3.711098, 3.864585, 4.018189, 4.17191, 4.325746, 4.479697, 4.63376, 
    4.787937, 4.942224, 5.096621, 5.251126, 5.405739, 5.560459, 5.715284, 
    5.870214, 6.025246, 6.18038, 6.335615, 6.490949, 6.646381, 6.801911, 
    6.957537, 7.113256, 7.26907, 7.424976, 7.580973, 7.73706, 7.893235, 
    8.049498, 8.205846, 8.36228, 8.518797, 8.675396, 8.832077, 8.988836, 
    9.145676, 9.302591, 9.459583, 9.61665, 9.773788, 9.931001, 10.08828, 
    10.24564, 10.40306, 10.56054, 10.71809, 10.87571, 11.03339, 11.19113, 
    11.34893, 11.50679, 11.66471, 11.82268, 11.98071, 12.13879, 12.29692, 
    12.4551, 12.61334, 12.77162, 12.92994, 13.08832, 13.24673, 13.40519, 
    13.56369, 13.72223, 13.8808, 14.03942, 14.19807, 14.35675, 14.51546, 
    14.67421, 14.83299, 14.99179, 15.15062, 15.30948, 15.46836, 15.62727, 
    15.78619, 15.94514, 16.1041, 16.26308, 16.42208, 16.58109, 16.74011, 
    16.89914, 17.05819, 17.21724, 17.3763, 17.53537, 17.69444, 17.85351, 
    18.01258, 18.17166, 18.33073, 18.4898, 18.64886, 18.80792, 18.96697, 
    19.12601, 19.28505, 19.44407, 19.60308, 19.76207, 19.92105, 20.08001, 
    20.23895, 20.39787, 20.55677, 20.71565, 20.8745, 21.03333, 21.19213, 
    21.3509, 21.50965, 21.66835, 21.82703, 21.98568, 22.14428, 22.30285, 
    22.46139, 22.61988, 22.77833, 22.93674, 23.09511, 23.25343, 23.4117, 
    23.56992, 23.7281, 23.88622, 24.04429, 24.20231, 24.36028, 24.51819, 
    24.67603, 24.83383, 24.99156, 25.14923, 25.30683, 25.46437, 25.62185, 
    25.77926, 25.9366, 26.09387, 26.25107, 26.4082, 26.56526, 26.72223, 
    26.87914, 27.03596, 27.19271, 27.34938, 27.50597, 27.66247, 27.81889, 
    27.97523, 28.13148, 28.28764, 28.44371, 28.59969, 28.75558, 28.91138, 
    29.06709, 29.2227, 29.37821, 29.53363, 29.68895, 29.84417, 29.99928, 
    30.1543, 30.30921, 30.46402, 30.61872, 30.77332, 30.92781, 31.08219, 
    31.23646, 31.39062, 31.54466, 31.6986, 31.85242, 32.00611, 32.1597, 
    32.31317, 32.46652, 32.61975, 32.77286, 32.92584, 33.0787, 33.23145, 
    33.38406, 33.53654, 33.68891, 33.84114, 33.99324, 34.14521, 34.29705, 
    34.44876, 34.60034, 34.75178, 34.90309, 35.05426, 35.20529, 35.35619, 
    35.50694, 35.65756, 35.80804, 35.95837, 36.10856, 36.25861, 36.40852, 
    36.55828, 36.70789, 36.85736, 37.00667, 37.15584, 37.30486, 37.45374, 
    37.60245, 37.75102, 37.89943, 38.0477, 38.1958, 38.34375, 38.49155, 
    38.63919, 38.78667, 38.93399, 39.08116, 39.22816, 39.37501, 39.52169, 
    39.66822, 39.81458, 39.96077, 40.1068, 40.25267, 40.39838, 40.54391, 
    40.68929, 40.83449, 40.97953, 41.12439, 41.26909, 41.41362, 41.55798, 
    41.70217, 41.84618, 41.99003, 42.1337, 42.2772, 42.42052, 42.56367, 
    42.70665, 42.84945, 42.99208, 43.13453, 43.2768, 43.41889, 43.56081, 
    43.70255, 43.8441, 43.98549, 44.12669,
  -20.48071, -20.35712, -20.23335, -20.10937, -19.9852, -19.86084, -19.73628, 
    -19.61153, -19.48658, -19.36143, -19.2361, -19.11056, -18.98483, 
    -18.85891, -18.73279, -18.60647, -18.47996, -18.35325, -18.22635, 
    -18.09925, -17.97196, -17.84447, -17.71678, -17.5889, -17.46082, 
    -17.33255, -17.20408, -17.07542, -16.94655, -16.8175, -16.68825, 
    -16.5588, -16.42915, -16.29931, -16.16928, -16.03905, -15.90862, -15.778, 
    -15.64718, -15.51617, -15.38496, -15.25356, -15.12196, -14.99017, 
    -14.85818, -14.726, -14.59362, -14.46105, -14.32828, -14.19532, 
    -14.06217, -13.92882, -13.79528, -13.66154, -13.52761, -13.39349, 
    -13.25917, -13.12466, -12.98996, -12.85506, -12.71998, -12.5847, 
    -12.44923, -12.31356, -12.17771, -12.04166, -11.90543, -11.769, 
    -11.63238, -11.49557, -11.35857, -11.22139, -11.08401, -10.94644, 
    -10.80869, -10.67074, -10.53261, -10.39429, -10.25578, -10.11709, 
    -9.978207, -9.839139, -9.699885, -9.560446, -9.42082, -9.28101, 
    -9.141015, -9.000836, -8.860474, -8.719927, -8.579198, -8.438287, 
    -8.297193, -8.155917, -8.014461, -7.872823, -7.731005, -7.589007, 
    -7.446831, -7.304475, -7.161941, -7.019228, -6.876339, -6.733273, 
    -6.590031, -6.446612, -6.303019, -6.159251, -6.015309, -5.871193, 
    -5.726905, -5.582444, -5.437811, -5.293007, -5.148033, -5.002888, 
    -4.857574, -4.712092, -4.566442, -4.420624, -4.274639, -4.128488, 
    -3.982172, -3.835691, -3.689046, -3.542238, -3.395267, -3.248134, 
    -3.10084, -2.953386, -2.805772, -2.657999, -2.510067, -2.361978, 
    -2.213732, -2.065331, -1.916774, -1.768063, -1.619199, -1.470181, 
    -1.321012, -1.171692, -1.022221, -0.8726008, -0.7228322, -0.5729158, 
    -0.4228526, -0.2726434, -0.1222891, 0.0282094, 0.1788512, 0.3296354, 
    0.4805612, 0.6316274, 0.7828334, 0.9341781, 1.08566, 1.23728, 1.389035, 
    1.540925, 1.692949, 1.845106, 1.997394, 2.149814, 2.302364, 2.455043, 
    2.607849, 2.760782, 2.913842, 3.067026, 3.220334, 3.373765, 3.527317, 
    3.68099, 3.834782, 3.988693, 4.142721, 4.296865, 4.451125, 4.605498, 
    4.759984, 4.914583, 5.069292, 5.22411, 5.379036, 5.53407, 5.68921, 
    5.844455, 5.999804, 6.155254, 6.310807, 6.466459, 6.622211, 6.77806, 
    6.934006, 7.090047, 7.246182, 7.402411, 7.558731, 7.715141, 7.87164, 
    8.028228, 8.184901, 8.34166, 8.498505, 8.655431, 8.812439, 8.969527, 
    9.126695, 9.28394, 9.441261, 9.598659, 9.756129, 9.913672, 10.07129, 
    10.22897, 10.38672, 10.54454, 10.70243, 10.86038, 11.01839, 11.17647, 
    11.33461, 11.4928, 11.65105, 11.80936, 11.96773, 12.12615, 12.28462, 
    12.44314, 12.60171, 12.76033, 12.919, 13.07771, 13.23646, 13.39526, 
    13.5541, 13.71298, 13.8719, 14.03085, 14.18984, 14.34887, 14.50793, 
    14.66702, 14.82613, 14.98528, 15.14446, 15.30366, 15.46288, 15.62213, 
    15.7814, 15.94069, 16.09999, 16.25932, 16.41866, 16.57801, 16.73738, 
    16.89676, 17.05615, 17.21555, 17.37495, 17.53436, 17.69377, 17.85319, 
    18.01261, 18.17203, 18.33144, 18.49086, 18.65027, 18.80967, 18.96906, 
    19.12845, 19.28783, 19.4472, 19.60655, 19.76589, 19.92521, 20.08451, 
    20.2438, 20.40306, 20.56231, 20.72153, 20.88072, 21.03989, 21.19904, 
    21.35815, 21.51724, 21.67629, 21.83531, 21.99429, 22.15324, 22.31215, 
    22.47103, 22.62986, 22.78865, 22.9474, 23.10611, 23.26476, 23.42338, 
    23.58194, 23.74045, 23.89892, 24.05733, 24.21568, 24.37398, 24.53223, 
    24.69041, 24.84854, 25.00661, 25.16461, 25.32255, 25.48042, 25.63824, 
    25.79598, 25.95365, 26.11125, 26.26879, 26.42624, 26.58363, 26.74094, 
    26.89817, 27.05533, 27.2124, 27.3694, 27.52631, 27.68314, 27.83989, 
    27.99655, 28.15312, 28.30961, 28.466, 28.62231, 28.77852, 28.93464, 
    29.09067, 29.2466, 29.40243, 29.55817, 29.71381, 29.86934, 30.02478, 
    30.18011, 30.33534, 30.49046, 30.64548, 30.80039, 30.95519, 31.10988, 
    31.26446, 31.41893, 31.57328, 31.72753, 31.88165, 32.03566, 32.18955, 
    32.34333, 32.49698, 32.65051, 32.80392, 32.95721, 33.11038, 33.26342, 
    33.41633, 33.56912, 33.72178, 33.87431, 34.0267, 34.17897, 34.33111, 
    34.48311, 34.63498, 34.78671, 34.93831, 35.08977, 35.24109, 35.39228, 
    35.54332, 35.69423, 35.84499, 35.99561, 36.14608, 36.29641, 36.4466, 
    36.59664, 36.74653, 36.89628, 37.04588, 37.19532, 37.34462, 37.49376, 
    37.64276, 37.7916, 37.94028, 38.08882, 38.23719, 38.38541, 38.53348, 
    38.68139, 38.82913, 38.97672, 39.12415, 39.27142, 39.41853, 39.56547, 
    39.71225, 39.85887, 40.00533, 40.15162, 40.29774, 40.4437, 40.58949, 
    40.73512, 40.88057, 41.02586, 41.17097, 41.31593, 41.4607, 41.60531, 
    41.74974, 41.894, 42.03809, 42.182, 42.32574, 42.46931, 42.6127, 
    42.75592, 42.89895, 43.04182, 43.1845, 43.327, 43.46933, 43.61148, 
    43.75345, 43.89524, 44.03685, 44.17828,
  -20.54914, -20.42542, -20.30151, -20.17739, -20.05309, -19.92859, 
    -19.80389, -19.679, -19.55391, -19.42862, -19.30314, -19.17746, 
    -19.05159, -18.92552, -18.79925, -18.67279, -18.54613, -18.41927, 
    -18.29222, -18.16497, -18.03752, -17.90988, -17.78204, -17.654, 
    -17.52577, -17.39734, -17.26871, -17.13989, -17.01087, -16.88165, 
    -16.75224, -16.62263, -16.49282, -16.36281, -16.23261, -16.10221, 
    -15.97162, -15.84083, -15.70984, -15.57866, -15.44728, -15.31571, 
    -15.18393, -15.05197, -14.9198, -14.78744, -14.65489, -14.52214, 
    -14.38919, -14.25605, -14.12271, -13.98918, -13.85545, -13.72153, 
    -13.58742, -13.45311, -13.3186, -13.1839, -13.04901, -12.91392, 
    -12.77864, -12.64317, -12.50751, -12.37165, -12.2356, -12.09935, 
    -11.96292, -11.82629, -11.68947, -11.55246, -11.41526, -11.27787, 
    -11.14029, -11.00251, -10.86455, -10.7264, -10.58806, -10.44953, 
    -10.31081, -10.1719, -10.03281, -9.893525, -9.754056, -9.6144, -9.474557, 
    -9.334528, -9.194313, -9.053913, -8.913328, -8.772559, -8.631606, 
    -8.490469, -8.349149, -8.207645, -8.065961, -7.924094, -7.782045, 
    -7.639816, -7.497406, -7.354817, -7.212048, -7.0691, -6.925974, -6.78267, 
    -6.639188, -6.49553, -6.351695, -6.207685, -6.063499, -5.919139, 
    -5.774605, -5.629898, -5.485018, -5.339965, -5.194741, -5.049346, 
    -4.90378, -4.758045, -4.612141, -4.466068, -4.319828, -4.17342, 
    -4.026846, -3.880106, -3.733201, -3.586132, -3.438899, -3.291503, 
    -3.143945, -2.996226, -2.848345, -2.700305, -2.552105, -2.403747, 
    -2.255231, -2.106559, -1.95773, -1.808746, -1.659607, -1.510314, 
    -1.360869, -1.211272, -1.061523, -0.9116237, -0.7615751, -0.6113778, 
    -0.4610327, -0.3105406, -0.1599026, -0.009119328, 0.1418082, 0.292879, 
    0.4440923, 0.5954471, 0.7469424, 0.8985773, 1.050351, 1.202262, 1.354311, 
    1.506494, 1.658813, 1.811266, 1.963851, 2.116568, 2.269416, 2.422394, 
    2.575501, 2.728735, 2.882096, 3.035583, 3.189194, 3.342929, 3.496787, 
    3.650765, 3.804864, 3.959083, 4.113419, 4.267873, 4.422442, 4.577126, 
    4.731924, 4.886834, 5.041856, 5.196988, 5.352229, 5.507578, 5.663034, 
    5.818595, 5.974261, 6.130031, 6.285902, 6.441874, 6.597946, 6.754116, 
    6.910383, 7.066746, 7.223205, 7.379756, 7.5364, 7.693135, 7.84996, 
    8.006873, 8.163874, 8.32096, 8.478131, 8.635386, 8.792724, 8.950142, 
    9.107639, 9.265215, 9.422868, 9.580596, 9.738399, 9.896275, 10.05422, 
    10.21224, 10.37033, 10.52848, 10.6867, 10.84499, 11.00334, 11.16175, 
    11.32022, 11.47876, 11.63735, 11.79599, 11.9547, 12.11345, 12.27227, 
    12.43113, 12.59004, 12.749, 12.908, 13.06706, 13.22615, 13.38529, 
    13.54448, 13.7037, 13.86296, 14.02226, 14.18159, 14.34096, 14.50036, 
    14.65979, 14.81925, 14.97875, 15.13826, 15.29781, 15.45738, 15.61697, 
    15.77658, 15.93622, 16.09587, 16.25554, 16.41523, 16.57493, 16.73464, 
    16.89437, 17.0541, 17.21384, 17.37359, 17.53335, 17.69311, 17.85287, 
    18.01264, 18.1724, 18.33216, 18.49192, 18.65168, 18.81143, 18.97117, 
    19.1309, 19.29062, 19.45034, 19.61003, 19.76972, 19.92938, 20.08904, 
    20.24866, 20.40828, 20.56787, 20.72743, 20.88697, 21.04649, 21.20597, 
    21.36543, 21.52486, 21.68425, 21.84362, 22.00294, 22.16224, 22.32149, 
    22.48071, 22.63988, 22.79902, 22.95811, 23.11715, 23.27615, 23.4351, 
    23.59401, 23.75286, 23.91166, 24.07041, 24.2291, 24.38774, 24.54633, 
    24.70485, 24.86331, 25.02171, 25.18005, 25.33833, 25.49654, 25.65468, 
    25.81276, 25.97077, 26.1287, 26.28657, 26.44436, 26.60208, 26.75972, 
    26.91728, 27.07476, 27.23217, 27.38949, 27.54674, 27.70389, 27.86097, 
    28.01795, 28.17485, 28.33166, 28.48838, 28.64501, 28.80155, 28.95799, 
    29.11434, 29.27059, 29.42675, 29.58281, 29.73876, 29.89462, 30.05037, 
    30.20602, 30.36156, 30.517, 30.67233, 30.82756, 30.98267, 31.13768, 
    31.29257, 31.44735, 31.60202, 31.75657, 31.911, 32.06532, 32.21952, 
    32.3736, 32.52756, 32.6814, 32.83511, 32.9887, 33.14217, 33.29551, 
    33.44873, 33.60181, 33.75477, 33.9076, 34.0603, 34.21286, 34.36529, 
    34.51759, 34.66975, 34.82178, 34.97367, 35.12542, 35.27703, 35.4285, 
    35.57984, 35.73103, 35.88208, 36.03298, 36.18374, 36.33435, 36.48483, 
    36.63515, 36.78532, 36.93534, 37.08522, 37.23495, 37.38452, 37.53394, 
    37.68321, 37.83232, 37.98128, 38.13008, 38.27874, 38.42723, 38.57556, 
    38.72373, 38.87175, 39.0196, 39.1673, 39.31483, 39.4622, 39.60941, 
    39.75645, 39.90333, 40.05004, 40.19659, 40.34297, 40.48919, 40.63523, 
    40.78111, 40.92682, 41.07236, 41.21772, 41.36292, 41.50795, 41.6528, 
    41.79748, 41.94199, 42.08632, 42.23048, 42.37446, 42.51826, 42.6619, 
    42.80535, 42.94863, 43.09172, 43.23464, 43.37738, 43.51995, 43.66233, 
    43.80453, 43.94655, 44.08839, 44.23004,
  -20.61776, -20.4939, -20.36985, -20.24561, -20.12116, -19.99652, -19.87169, 
    -19.74665, -19.62142, -19.496, -19.37037, -19.24455, -19.11853, 
    -18.99232, -18.8659, -18.73929, -18.61248, -18.48548, -18.35828, 
    -18.23088, -18.10328, -17.97548, -17.84749, -17.7193, -17.59091, 
    -17.46232, -17.33353, -17.20455, -17.07537, -16.94599, -16.81642, 
    -16.68664, -16.55667, -16.4265, -16.29613, -16.16557, -16.03481, 
    -15.90385, -15.77269, -15.64134, -15.50979, -15.37804, -15.24609, 
    -15.11395, -14.98161, -14.84907, -14.71634, -14.58341, -14.45029, 
    -14.31696, -14.18344, -14.04973, -13.91582, -13.78171, -13.64741, 
    -13.51291, -13.37822, -13.24333, -13.10825, -12.97297, -12.8375, 
    -12.70183, -12.56597, -12.42992, -12.29367, -12.15723, -12.0206, 
    -11.88377, -11.74675, -11.60954, -11.47213, -11.33454, -11.19675, 
    -11.05877, -10.9206, -10.78224, -10.64369, -10.50495, -10.36602, 
    -10.2269, -10.08759, -9.948092, -9.808407, -9.668533, -9.528473, 
    -9.388225, -9.247789, -9.107168, -8.966361, -8.825369, -8.684191, 
    -8.542829, -8.401281, -8.259551, -8.117637, -7.97554, -7.833261, 
    -7.690799, -7.548156, -7.405333, -7.262328, -7.119144, -6.97578, 
    -6.832238, -6.688517, -6.544618, -6.400541, -6.256288, -6.111859, 
    -5.967254, -5.822474, -5.677519, -5.532391, -5.387089, -5.241615, 
    -5.095969, -4.950151, -4.804163, -4.658004, -4.511675, -4.365178, 
    -4.218513, -4.071681, -3.924681, -3.777515, -3.630184, -3.482689, 
    -3.335029, -3.187206, -3.039221, -2.891073, -2.742765, -2.594297, 
    -2.445669, -2.296882, -2.147938, -1.998836, -1.849578, -1.700164, 
    -1.550596, -1.400873, -1.250998, -1.100971, -0.9507915, -0.8004621, 
    -0.649983, -0.4993552, -0.3485795, -0.1976567, -0.04658788, 0.1046262, 
    0.2559845, 0.4074862, 0.5591304, 0.710916, 0.8628422, 1.014908, 1.167112, 
    1.319455, 1.471933, 1.624548, 1.777297, 1.93018, 2.083196, 2.236343, 
    2.389621, 2.543029, 2.696565, 2.850229, 3.004019, 3.157935, 3.311975, 
    3.466139, 3.620424, 3.774831, 3.929358, 4.084004, 4.238768, 4.393648, 
    4.548644, 4.703754, 4.858978, 5.014314, 5.169761, 5.325317, 5.480983, 
    5.636755, 5.792635, 5.948619, 6.104708, 6.260899, 6.417192, 6.573585, 
    6.730077, 6.886667, 7.043354, 7.200136, 7.357012, 7.513981, 7.671042, 
    7.828194, 7.985434, 8.142762, 8.300178, 8.457678, 8.615262, 8.772929, 
    8.930678, 9.088507, 9.246415, 9.4044, 9.562461, 9.720597, 9.878807, 
    10.03709, 10.19544, 10.35386, 10.51236, 10.67091, 10.82954, 10.98822, 
    11.14697, 11.30578, 11.46465, 11.62358, 11.78257, 11.94162, 12.10071, 
    12.25986, 12.41907, 12.57832, 12.73762, 12.89697, 13.05636, 13.2158, 
    13.37529, 13.53481, 13.69438, 13.85398, 14.01362, 14.1733, 14.33301, 
    14.49276, 14.65254, 14.81235, 14.97218, 15.13205, 15.29194, 15.45185, 
    15.61179, 15.77175, 15.93173, 16.09173, 16.25175, 16.41178, 16.57183, 
    16.73189, 16.89196, 17.05204, 17.21213, 17.37223, 17.53233, 17.69244, 
    17.85255, 18.01266, 18.17278, 18.33289, 18.49299, 18.6531, 18.81319, 
    18.97328, 19.13336, 19.29343, 19.45349, 19.61353, 19.77357, 19.93358, 
    20.09357, 20.25355, 20.41351, 20.57344, 20.73336, 20.89324, 21.0531, 
    21.21294, 21.37274, 21.53251, 21.69225, 21.85196, 22.01163, 22.17127, 
    22.33087, 22.49043, 22.64994, 22.80942, 22.96885, 23.12824, 23.28758, 
    23.44688, 23.60612, 23.76532, 23.92446, 24.08355, 24.24258, 24.40156, 
    24.56048, 24.71934, 24.87814, 25.03688, 25.19556, 25.35417, 25.51272, 
    25.6712, 25.82961, 25.98795, 26.14622, 26.30442, 26.46255, 26.6206, 
    26.77857, 26.93646, 27.09428, 27.25202, 27.40967, 27.56724, 27.72473, 
    27.88213, 28.03944, 28.19667, 28.35381, 28.51085, 28.66781, 28.82467, 
    28.98144, 29.13811, 29.29469, 29.45116, 29.60754, 29.76381, 29.91999, 
    30.07606, 30.23203, 30.38789, 30.54365, 30.6993, 30.85484, 31.01027, 
    31.16558, 31.32079, 31.47588, 31.63086, 31.78572, 31.94047, 32.09509, 
    32.2496, 32.40399, 32.55825, 32.7124, 32.86642, 33.02032, 33.17409, 
    33.32773, 33.48125, 33.63463, 33.78789, 33.94102, 34.09401, 34.24688, 
    34.3996, 34.5522, 34.70465, 34.85697, 35.00916, 35.1612, 35.3131, 
    35.46487, 35.61649, 35.76797, 35.9193, 36.0705, 36.22154, 36.37244, 
    36.52319, 36.6738, 36.82425, 36.97456, 37.12471, 37.27472, 37.42457, 
    37.57426, 37.72381, 37.8732, 38.02243, 38.17151, 38.32043, 38.46919, 
    38.61779, 38.76624, 38.91452, 39.06264, 39.2106, 39.3584, 39.50603, 
    39.6535, 39.8008, 39.94794, 40.09492, 40.24173, 40.38836, 40.53483, 
    40.68113, 40.82727, 40.97323, 41.11902, 41.26464, 41.41008, 41.55536, 
    41.70046, 41.84539, 41.99014, 42.13472, 42.27912, 42.42334, 42.56739, 
    42.71126, 42.85496, 42.99847, 43.1418, 43.28496, 43.42794, 43.57073, 
    43.71334, 43.85578, 43.99803, 44.1401, 44.28198,
  -20.68656, -20.56257, -20.43839, -20.314, -20.18942, -20.06465, -19.93967, 
    -19.8145, -19.68913, -19.56356, -19.43779, -19.31183, -19.18567, 
    -19.0593, -18.93274, -18.80599, -18.67903, -18.55188, -18.42452, 
    -18.29697, -18.16922, -18.04127, -17.91312, -17.78478, -17.65623, 
    -17.52749, -17.39854, -17.2694, -17.14006, -17.01052, -16.88079, 
    -16.75085, -16.62071, -16.49038, -16.35985, -16.22912, -16.09819, 
    -15.96706, -15.83573, -15.70421, -15.57248, -15.44056, -15.30844, 
    -15.17613, -15.04361, -14.9109, -14.77799, -14.64488, -14.51157, 
    -14.37807, -14.24437, -14.11047, -13.97637, -13.84208, -13.70759, 
    -13.57291, -13.43803, -13.30295, -13.16768, -13.03221, -12.89654, 
    -12.76068, -12.62463, -12.48838, -12.35193, -12.21529, -12.07846, 
    -11.94143, -11.80421, -11.6668, -11.52919, -11.39139, -11.2534, 
    -11.11521, -10.97683, -10.83826, -10.6995, -10.56055, -10.42141, 
    -10.28208, -10.14255, -10.00284, -9.86294, -9.722849, -9.58257, 
    -9.442102, -9.301447, -9.160604, -9.019573, -8.878357, -8.736954, 
    -8.595366, -8.453591, -8.311633, -8.16949, -8.027163, -7.884652, 
    -7.741958, -7.599081, -7.456023, -7.312783, -7.169362, -7.02576, 
    -6.881979, -6.738017, -6.593877, -6.449558, -6.305062, -6.160388, 
    -6.015538, -5.870512, -5.725309, -5.579932, -5.434381, -5.288656, 
    -5.142757, -4.996686, -4.850444, -4.704031, -4.557446, -4.410692, 
    -4.263768, -4.116676, -3.969417, -3.82199, -3.674396, -3.526637, 
    -3.378713, -3.230625, -3.082373, -2.933958, -2.785381, -2.636643, 
    -2.487744, -2.338686, -2.189469, -2.040093, -1.89056, -1.740871, 
    -1.591026, -1.441026, -1.290872, -1.140565, -0.9901053, -0.8394943, 
    -0.6887326, -0.5378212, -0.3867609, -0.2355526, -0.08419731, 0.06730418, 
    0.2189509, 0.3707419, 0.5226763, 0.6747532, 0.8269715, 0.9793304, 
    1.131829, 1.284466, 1.43724, 1.590152, 1.743199, 1.89638, 2.049695, 
    2.203143, 2.356722, 2.510432, 2.664271, 2.818238, 2.972334, 3.126555, 
    3.280901, 3.435372, 3.589966, 3.744681, 3.899518, 4.054474, 4.209549, 
    4.364742, 4.520051, 4.675475, 4.831013, 4.986664, 5.142426, 5.2983, 
    5.454283, 5.610374, 5.766572, 5.922876, 6.079285, 6.235797, 6.392412, 
    6.549127, 6.705943, 6.862856, 7.019868, 7.176975, 7.334177, 7.491473, 
    7.648861, 7.806341, 7.96391, 8.121567, 8.279312, 8.437142, 8.595057, 
    8.753057, 8.911137, 9.069299, 9.227539, 9.385859, 9.544253, 9.702724, 
    9.86127, 10.01989, 10.17858, 10.33734, 10.49616, 10.65506, 10.81402, 
    10.97305, 11.13214, 11.29129, 11.4505, 11.60977, 11.7691, 11.92848, 
    12.08792, 12.24741, 12.40696, 12.56655, 12.7262, 12.88589, 13.04563, 
    13.20541, 13.36524, 13.52511, 13.68502, 13.84497, 14.00496, 14.16498, 
    14.32504, 14.48513, 14.64525, 14.80541, 14.96559, 15.1258, 15.28604, 
    15.44631, 15.60659, 15.7669, 15.92723, 16.08758, 16.24794, 16.40832, 
    16.56872, 16.72913, 16.88955, 17.04998, 17.21042, 17.37086, 17.53131, 
    17.69177, 17.85223, 18.01269, 18.17315, 18.33361, 18.49407, 18.65452, 
    18.81496, 18.9754, 19.13583, 19.29625, 19.45666, 19.61705, 19.77743, 
    19.93779, 20.09813, 20.25846, 20.41876, 20.57905, 20.73931, 20.89954, 
    21.05975, 21.21993, 21.38008, 21.5402, 21.70028, 21.86034, 22.02036, 
    22.18034, 22.34028, 22.50018, 22.66005, 22.81987, 22.97964, 23.13938, 
    23.29906, 23.4587, 23.61828, 23.77782, 23.93731, 24.09674, 24.25611, 
    24.41543, 24.57469, 24.73389, 24.89303, 25.05211, 25.21113, 25.37008, 
    25.52896, 25.68778, 25.84653, 26.00521, 26.16381, 26.32235, 26.48081, 
    26.63919, 26.7975, 26.95572, 27.11387, 27.27194, 27.42993, 27.58783, 
    27.74565, 27.90338, 28.06102, 28.21858, 28.37604, 28.53341, 28.6907, 
    28.84788, 29.00498, 29.16197, 29.31887, 29.47567, 29.63237, 29.78897, 
    29.94546, 30.10186, 30.25814, 30.41432, 30.5704, 30.72636, 30.88222, 
    31.03797, 31.1936, 31.34912, 31.50452, 31.65981, 31.81499, 31.97005, 
    32.12498, 32.2798, 32.4345, 32.58907, 32.74352, 32.89785, 33.05205, 
    33.20612, 33.36007, 33.51389, 33.66758, 33.82114, 33.97457, 34.12786, 
    34.28102, 34.43404, 34.58694, 34.73969, 34.8923, 35.04478, 35.19712, 
    35.34931, 35.50137, 35.65328, 35.80505, 35.95667, 36.10815, 36.25948, 
    36.41067, 36.5617, 36.71259, 36.86333, 37.01392, 37.16435, 37.31464, 
    37.46476, 37.61474, 37.76456, 37.91422, 38.06373, 38.21308, 38.36227, 
    38.51131, 38.66018, 38.8089, 38.95745, 39.10583, 39.25406, 39.40212, 
    39.55002, 39.69775, 39.84532, 39.99272, 40.13995, 40.28702, 40.43392, 
    40.58065, 40.7272, 40.87359, 41.01981, 41.16585, 41.31172, 41.45742, 
    41.60294, 41.74829, 41.89346, 42.03846, 42.18328, 42.32793, 42.4724, 
    42.61669, 42.7608, 42.90474, 43.04849, 43.19206, 43.33545, 43.47866, 
    43.62169, 43.76454, 43.90721, 44.04969, 44.19199, 44.3341,
  -20.75556, -20.63143, -20.50711, -20.38259, -20.25788, -20.13296, 
    -20.00785, -19.88253, -19.75702, -19.63131, -19.5054, -19.3793, 
    -19.25299, -19.12648, -18.99978, -18.87287, -18.74577, -18.61846, 
    -18.49096, -18.36326, -18.23536, -18.10725, -17.97895, -17.85045, 
    -17.72175, -17.59285, -17.46375, -17.33445, -17.20495, -17.07525, 
    -16.94535, -16.81525, -16.68495, -16.55445, -16.42375, -16.29285, 
    -16.16176, -16.03046, -15.89896, -15.76727, -15.63537, -15.50328, 
    -15.37098, -15.23849, -15.1058, -14.97291, -14.83982, -14.70653, 
    -14.57304, -14.43936, -14.30548, -14.1714, -14.03712, -13.90264, 
    -13.76796, -13.63309, -13.49802, -13.36275, -13.22729, -13.09163, 
    -12.95577, -12.81972, -12.68347, -12.54702, -12.41038, -12.27354, 
    -12.13651, -11.99928, -11.86186, -11.72424, -11.58643, -11.44843, 
    -11.31023, -11.17184, -11.03325, -10.89447, -10.7555, -10.61634, 
    -10.47698, -10.33744, -10.1977, -10.05777, -9.917655, -9.777347, 
    -9.636848, -9.496161, -9.355285, -9.214219, -9.072967, -8.931525, 
    -8.789897, -8.648083, -8.506081, -8.363894, -8.22152, -8.078962, 
    -7.93622, -7.793293, -7.650182, -7.506889, -7.363412, -7.219754, 
    -7.075914, -6.931893, -6.787691, -6.643309, -6.498748, -6.354007, 
    -6.209089, -6.063993, -5.918719, -5.773269, -5.627642, -5.481841, 
    -5.335864, -5.189713, -5.043389, -4.896892, -4.750222, -4.603381, 
    -4.456369, -4.309187, -4.161835, -4.014314, -3.866625, -3.718769, 
    -3.570746, -3.422556, -3.274202, -3.125682, -2.977, -2.828153, -2.679145, 
    -2.529975, -2.380644, -2.231153, -2.081503, -1.931695, -1.781729, 
    -1.631607, -1.481328, -1.330895, -1.180307, -1.029566, -0.8786727, 
    -0.7276275, -0.5764316, -0.425086, -0.2735913, -0.1219486, 0.02984118, 
    0.1817772, 0.3338584, 0.486084, 0.638453, 0.7909644, 0.9436173, 1.096411, 
    1.249344, 1.402415, 1.555624, 1.708969, 1.86245, 2.016066, 2.169815, 
    2.323696, 2.477709, 2.631852, 2.786124, 2.940525, 3.095053, 3.249707, 
    3.404486, 3.559389, 3.714414, 3.869561, 4.024829, 4.180217, 4.335722, 
    4.491345, 4.647084, 4.802938, 4.958905, 5.114985, 5.271176, 5.427477, 
    5.583888, 5.740407, 5.897031, 6.053761, 6.210596, 6.367534, 6.524573, 
    6.681713, 6.838952, 6.996289, 7.153722, 7.311252, 7.468875, 7.626592, 
    7.7844, 7.942299, 8.100286, 8.258363, 8.416525, 8.574772, 8.733104, 
    8.891518, 9.050013, 9.208588, 9.367242, 9.525972, 9.68478, 9.843661, 
    10.00262, 10.16164, 10.32074, 10.47991, 10.63914, 10.79844, 10.95781, 
    11.11724, 11.27673, 11.43628, 11.59589, 11.75556, 11.91529, 12.07507, 
    12.23491, 12.3948, 12.55474, 12.71473, 12.87476, 13.03485, 13.19498, 
    13.35515, 13.51536, 13.67562, 13.83592, 13.99625, 14.15662, 14.31703, 
    14.47747, 14.63794, 14.79844, 14.95898, 15.11954, 15.28012, 15.44073, 
    15.60137, 15.76203, 15.92271, 16.0834, 16.24412, 16.40485, 16.56559, 
    16.72635, 16.88712, 17.0479, 17.20869, 17.36949, 17.53029, 17.6911, 
    17.85191, 18.01272, 18.17353, 18.33434, 18.49515, 18.65595, 18.81674, 
    18.97753, 19.13831, 19.29908, 19.45984, 19.62058, 19.78131, 19.94202, 
    20.10271, 20.26339, 20.42404, 20.58467, 20.74528, 20.90586, 21.06642, 
    21.22695, 21.38745, 21.54791, 21.70835, 21.86875, 22.02911, 22.18944, 
    22.34973, 22.50998, 22.67019, 22.83036, 22.99048, 23.15055, 23.31059, 
    23.47057, 23.6305, 23.79038, 23.9502, 24.10998, 24.2697, 24.42936, 
    24.58896, 24.7485, 24.90799, 25.06741, 25.22676, 25.38605, 25.54527, 
    25.70443, 25.86352, 26.02253, 26.18148, 26.34035, 26.49914, 26.65786, 
    26.8165, 26.97506, 27.13355, 27.29195, 27.45027, 27.6085, 27.76665, 
    27.92471, 28.08268, 28.24057, 28.39836, 28.55606, 28.71367, 28.87119, 
    29.02861, 29.18593, 29.34315, 29.50027, 29.6573, 29.81422, 29.97104, 
    30.12775, 30.28436, 30.44086, 30.59725, 30.75354, 30.90971, 31.06577, 
    31.22172, 31.37756, 31.53328, 31.68888, 31.84437, 31.99974, 32.15499, 
    32.31012, 32.46512, 32.62001, 32.77477, 32.9294, 33.08391, 33.23829, 
    33.39254, 33.54666, 33.70065, 33.85452, 34.00824, 34.16184, 34.3153, 
    34.46862, 34.62181, 34.77486, 34.92777, 35.08054, 35.23317, 35.38566, 
    35.53801, 35.69021, 35.84227, 35.99418, 36.14595, 36.29757, 36.44904, 
    36.60036, 36.75153, 36.90255, 37.05342, 37.20414, 37.3547, 37.50511, 
    37.65536, 37.80546, 37.9554, 38.10519, 38.25481, 38.40428, 38.55358, 
    38.70273, 38.85171, 39.00053, 39.14919, 39.29768, 39.44601, 39.59417, 
    39.74217, 39.89, 40.03766, 40.18515, 40.33248, 40.47964, 40.62662, 
    40.77343, 40.92008, 41.06655, 41.21284, 41.35897, 41.50492, 41.65069, 
    41.79629, 41.94171, 42.08696, 42.23203, 42.37691, 42.52163, 42.66616, 
    42.81051, 42.95469, 43.09868, 43.24249, 43.38612, 43.52957, 43.67283, 
    43.81591, 43.95881, 44.10152, 44.24405, 44.3864,
  -20.82474, -20.70048, -20.57603, -20.45137, -20.32652, -20.20147, 
    -20.07621, -19.95076, -19.82511, -19.69926, -19.57321, -19.44695, 
    -19.3205, -19.19385, -19.067, -18.93995, -18.81269, -18.68524, -18.55759, 
    -18.42974, -18.30168, -18.17343, -18.04497, -17.91632, -17.78746, 
    -17.6584, -17.52914, -17.39968, -17.27002, -17.14016, -17.0101, 
    -16.87984, -16.74937, -16.61871, -16.48785, -16.35678, -16.22552, 
    -16.09405, -15.96239, -15.83052, -15.69845, -15.56618, -15.43372, 
    -15.30105, -15.16818, -15.03511, -14.90184, -14.76838, -14.63471, 
    -14.50084, -14.36678, -14.23251, -14.09805, -13.96339, -13.82853, 
    -13.69347, -13.55821, -13.42275, -13.2871, -13.15124, -13.01519, 
    -12.87894, -12.7425, -12.60586, -12.46902, -12.33198, -12.19475, 
    -12.05732, -11.9197, -11.78188, -11.64386, -11.50565, -11.36725, 
    -11.22865, -11.08986, -10.95087, -10.81169, -10.67231, -10.53275, 
    -10.39299, -10.25303, -10.11289, -9.972554, -9.832028, -9.691311, 
    -9.550403, -9.409305, -9.268018, -9.126541, -8.984876, -8.843021, 
    -8.700979, -8.55875, -8.416334, -8.27373, -8.130941, -7.987966, 
    -7.844806, -7.701461, -7.557932, -7.414218, -7.270322, -7.126243, 
    -6.981982, -6.837539, -6.692915, -6.54811, -6.403126, -6.257962, 
    -6.112619, -5.967097, -5.821398, -5.675522, -5.529469, -5.383241, 
    -5.236837, -5.090259, -4.943507, -4.796581, -4.649482, -4.502212, 
    -4.35477, -4.207158, -4.059375, -3.911423, -3.763303, -3.615015, 
    -3.46656, -3.317939, -3.169151, -3.020199, -2.871083, -2.721803, 
    -2.572361, -2.422757, -2.272993, -2.123067, -1.972983, -1.82274, 
    -1.672339, -1.521781, -1.371068, -1.220199, -1.069175, -0.9179983, 
    -0.7666689, -0.6151877, -0.4635557, -0.3117738, -0.1598429, -0.007763894, 
    0.1444623, 0.2968347, 0.4493524, 0.6020144, 0.7548198, 0.9077676, 
    1.060857, 1.214087, 1.367456, 1.520963, 1.674608, 1.82839, 1.982307, 
    2.136358, 2.290543, 2.44486, 2.599308, 2.753886, 2.908593, 3.063429, 
    3.218391, 3.373479, 3.528692, 3.684029, 3.839488, 3.995068, 4.150769, 
    4.306589, 4.462527, 4.618581, 4.774752, 4.931036, 5.087435, 5.243945, 
    5.400566, 5.557297, 5.714137, 5.871084, 6.028137, 6.185295, 6.342556, 
    6.499921, 6.657386, 6.814951, 6.972615, 7.130377, 7.288235, 7.446187, 
    7.604233, 7.762372, 7.920601, 8.078921, 8.237329, 8.395823, 8.554404, 
    8.71307, 8.871819, 9.030649, 9.18956, 9.34855, 9.507618, 9.666762, 
    9.825982, 9.985275, 10.14464, 10.30408, 10.46358, 10.62316, 10.7828, 
    10.94251, 11.10228, 11.26211, 11.42201, 11.58196, 11.74198, 11.90205, 
    12.06217, 12.22235, 12.38259, 12.54287, 12.70321, 12.86359, 13.02402, 
    13.1845, 13.34502, 13.50558, 13.66619, 13.82683, 13.98751, 14.14823, 
    14.30899, 14.46978, 14.6306, 14.79145, 14.95233, 15.11324, 15.27418, 
    15.43514, 15.59613, 15.75714, 15.91816, 16.07921, 16.24028, 16.40136, 
    16.56246, 16.72357, 16.88469, 17.04582, 17.20696, 17.36811, 17.52926, 
    17.69042, 17.85158, 18.01275, 18.17391, 18.33507, 18.49623, 18.65738, 
    18.81853, 18.97967, 19.1408, 19.30192, 19.46303, 19.62412, 19.7852, 
    19.94626, 20.10731, 20.26834, 20.42934, 20.59032, 20.75128, 20.91221, 
    21.07312, 21.234, 21.39484, 21.55566, 21.71644, 21.87719, 22.03791, 
    22.19858, 22.35922, 22.51982, 22.68038, 22.84089, 23.00136, 23.16178, 
    23.32216, 23.48248, 23.64276, 23.80299, 23.96316, 24.12328, 24.28334, 
    24.44334, 24.60329, 24.76317, 24.923, 25.08276, 25.24246, 25.40209, 
    25.56165, 25.72115, 25.88057, 26.03993, 26.19921, 26.35842, 26.51755, 
    26.67661, 26.83558, 26.99448, 27.1533, 27.31203, 27.47069, 27.62925, 
    27.78773, 27.94613, 28.10443, 28.26265, 28.42077, 28.5788, 28.73674, 
    28.89458, 29.05233, 29.20998, 29.36753, 29.52498, 29.68233, 29.83957, 
    29.99671, 30.15375, 30.31068, 30.4675, 30.62422, 30.78082, 30.93731, 
    31.09369, 31.24996, 31.40611, 31.56215, 31.71807, 31.87387, 32.02955, 
    32.18511, 32.34055, 32.49587, 32.65106, 32.80613, 32.96107, 33.11589, 
    33.27058, 33.42513, 33.57956, 33.73386, 33.88802, 34.04205, 34.19595, 
    34.3497, 34.50333, 34.65681, 34.81016, 34.96337, 35.11644, 35.26936, 
    35.42214, 35.57478, 35.72728, 35.87963, 36.03183, 36.18389, 36.33579, 
    36.48755, 36.63916, 36.79062, 36.94192, 37.09307, 37.24408, 37.39492, 
    37.54561, 37.69614, 37.84652, 37.99673, 38.14679, 38.29669, 38.44643, 
    38.59601, 38.74543, 38.89468, 39.04377, 39.1927, 39.34146, 39.49006, 
    39.63848, 39.78674, 39.93484, 40.08276, 40.23052, 40.37811, 40.52552, 
    40.67276, 40.81983, 40.96673, 41.11346, 41.26001, 41.40638, 41.55259, 
    41.69861, 41.84446, 41.99013, 42.13562, 42.28094, 42.42607, 42.57103, 
    42.71581, 42.8604, 43.00481, 43.14905, 43.2931, 43.43696, 43.58065, 
    43.72415, 43.86746, 44.01059, 44.15354, 44.2963, 44.43887,
  -20.89411, -20.76972, -20.64513, -20.52034, -20.39535, -20.27016, 
    -20.14477, -20.01918, -19.89339, -19.7674, -19.6412, -19.51481, 
    -19.38821, -19.26141, -19.13442, -19.00722, -18.87982, -18.75221, 
    -18.62441, -18.49641, -18.3682, -18.23979, -18.11118, -17.98237, 
    -17.85336, -17.72415, -17.59473, -17.46511, -17.33529, -17.20527, 
    -17.07505, -16.94462, -16.814, -16.68317, -16.55214, -16.42091, 
    -16.28947, -16.15784, -16.026, -15.89396, -15.76172, -15.62928, 
    -15.49664, -15.3638, -15.23075, -15.09751, -14.96406, -14.83042, 
    -14.69657, -14.56252, -14.42827, -14.29383, -14.15918, -14.02433, 
    -13.88928, -13.75403, -13.61858, -13.48294, -13.34709, -13.21105, 
    -13.0748, -12.93836, -12.80172, -12.66488, -12.52785, -12.39061, 
    -12.25318, -12.11555, -11.97772, -11.8397, -11.70148, -11.56307, 
    -11.42446, -11.28565, -11.14665, -11.00745, -10.86806, -10.72847, 
    -10.58869, -10.44872, -10.30855, -10.16819, -10.02764, -9.886894, 
    -9.745957, -9.604829, -9.46351, -9.321999, -9.180299, -9.038408, 
    -8.896328, -8.754059, -8.611601, -8.468955, -8.326121, -8.183101, 
    -8.039892, -7.896498, -7.752918, -7.609153, -7.465202, -7.321068, 
    -7.17675, -7.032248, -6.887563, -6.742696, -6.597648, -6.452418, 
    -6.307008, -6.161418, -6.015648, -5.8697, -5.723574, -5.57727, -5.430789, 
    -5.284131, -5.137298, -4.99029, -4.843107, -4.69575, -4.548221, 
    -4.400519, -4.252645, -4.1046, -3.956385, -3.808001, -3.659447, 
    -3.510725, -3.361836, -3.21278, -3.063559, -2.914172, -2.76462, 
    -2.614905, -2.465027, -2.314987, -2.164786, -2.014425, -1.863904, 
    -1.713224, -1.562386, -1.411391, -1.26024, -1.108933, -0.9574723, 
    -0.8058577, -0.6540904, -0.5021713, -0.3501012, -0.1978812, -0.04551208, 
    0.1070052, 0.2596696, 0.4124803, 0.5654363, 0.7185367, 0.8717803, 
    1.025166, 1.178694, 1.332362, 1.486169, 1.640115, 1.794198, 1.948417, 
    2.102771, 2.25726, 2.411882, 2.566636, 2.721521, 2.876537, 3.031681, 
    3.186952, 3.342351, 3.497875, 3.653524, 3.809296, 3.96519, 4.121205, 
    4.27734, 4.433595, 4.589966, 4.746454, 4.903058, 5.059775, 5.216606, 
    5.373548, 5.530601, 5.687763, 5.845033, 6.00241, 6.159893, 6.31748, 
    6.47517, 6.632962, 6.790855, 6.948847, 7.106937, 7.265125, 7.423408, 
    7.581785, 7.740255, 7.898817, 8.057468, 8.21621, 8.375039, 8.533955, 
    8.692955, 8.852039, 9.011207, 9.170455, 9.329782, 9.489188, 9.648672, 
    9.80823, 9.967864, 10.12757, 10.28735, 10.4472, 10.60711, 10.7671, 
    10.92715, 11.08726, 11.24744, 11.40768, 11.56798, 11.72834, 11.88875, 
    12.04922, 12.20975, 12.37033, 12.53096, 12.69164, 12.85238, 13.01315, 
    13.17398, 13.33485, 13.49576, 13.65671, 13.81771, 13.97874, 14.13981, 
    14.30091, 14.46205, 14.62322, 14.78443, 14.94566, 15.10692, 15.26821, 
    15.42953, 15.59086, 15.75222, 15.9136, 16.075, 16.23642, 16.39786, 
    16.55931, 16.72077, 16.88224, 17.04373, 17.20522, 17.36672, 17.52823, 
    17.68974, 17.85126, 18.01278, 18.17429, 18.3358, 18.49732, 18.65882, 
    18.82032, 18.98182, 19.1433, 19.30477, 19.46623, 19.62768, 19.78911, 
    19.95053, 20.11193, 20.2733, 20.43466, 20.59599, 20.7573, 20.91859, 
    21.07985, 21.24107, 21.40227, 21.56344, 21.72458, 21.88567, 22.04674, 
    22.20776, 22.36875, 22.5297, 22.6906, 22.85147, 23.01228, 23.17305, 
    23.33378, 23.49445, 23.65508, 23.81565, 23.97616, 24.13663, 24.29704, 
    24.45738, 24.61767, 24.7779, 24.93807, 25.09818, 25.25822, 25.41819, 
    25.57809, 25.73793, 25.8977, 26.05739, 26.21701, 26.37656, 26.53603, 
    26.69543, 26.85474, 27.01398, 27.17313, 27.3322, 27.49119, 27.65009, 
    27.80891, 27.96763, 28.12627, 28.28482, 28.44327, 28.60164, 28.7599, 
    28.91808, 29.07615, 29.23413, 29.392, 29.54978, 29.70745, 29.86503, 
    30.02249, 30.17985, 30.3371, 30.49425, 30.65129, 30.80821, 30.96502, 
    31.12172, 31.27831, 31.43478, 31.59113, 31.74737, 31.90348, 32.05948, 
    32.21535, 32.37111, 32.52673, 32.68224, 32.83762, 32.99287, 33.14799, 
    33.30299, 33.45785, 33.61259, 33.76719, 33.92165, 34.07599, 34.23019, 
    34.38425, 34.53817, 34.69196, 34.8456, 34.99911, 35.15247, 35.30569, 
    35.45877, 35.6117, 35.76449, 35.91713, 36.06963, 36.22197, 36.37416, 
    36.52621, 36.67811, 36.82985, 36.98144, 37.13288, 37.28416, 37.43529, 
    37.58626, 37.73707, 37.88773, 38.03822, 38.18856, 38.33873, 38.48875, 
    38.6386, 38.78829, 38.93781, 39.08717, 39.23637, 39.3854, 39.53426, 
    39.68296, 39.83149, 39.97984, 40.12803, 40.27605, 40.42389, 40.57157, 
    40.71907, 40.8664, 41.01356, 41.16054, 41.30734, 41.45397, 41.60043, 
    41.7467, 41.8928, 42.03872, 42.18446, 42.33002, 42.4754, 42.62061, 
    42.76562, 42.91046, 43.05512, 43.19959, 43.34388, 43.48798, 43.63191, 
    43.77564, 43.91919, 44.06256, 44.20574, 44.34873, 44.49153,
  -20.96368, -20.83916, -20.71443, -20.58951, -20.46438, -20.33905, 
    -20.21352, -20.08779, -19.96186, -19.83572, -19.70939, -19.58285, 
    -19.45611, -19.32917, -19.20203, -19.07468, -18.94713, -18.81938, 
    -18.69143, -18.56327, -18.43492, -18.30635, -18.17759, -18.04863, 
    -17.91946, -17.79009, -17.66051, -17.53074, -17.40075, -17.27057, 
    -17.14019, -17.0096, -16.87881, -16.74782, -16.61662, -16.48522, 
    -16.35362, -16.22182, -16.08981, -15.9576, -15.82519, -15.69258, 
    -15.55976, -15.42674, -15.29352, -15.1601, -15.02648, -14.89265, 
    -14.75862, -14.62439, -14.48996, -14.35533, -14.2205, -14.08546, 
    -13.95023, -13.81479, -13.67916, -13.54332, -13.40728, -13.27104, 
    -13.13461, -12.99797, -12.86113, -12.7241, -12.58686, -12.44943, 
    -12.3118, -12.17397, -12.03594, -11.89771, -11.75929, -11.62067, 
    -11.48185, -11.34284, -11.20363, -11.06422, -10.92462, -10.78482, 
    -10.64483, -10.50464, -10.36426, -10.22368, -10.08291, -9.941946, 
    -9.80079, -9.65944, -9.517899, -9.376165, -9.234241, -9.092124, 
    -8.949818, -8.807321, -8.664634, -8.521758, -8.378694, -8.23544, 
    -8.091999, -7.948371, -7.804555, -7.660553, -7.516366, -7.371992, 
    -7.227434, -7.082691, -6.937764, -6.792654, -6.647361, -6.501886, 
    -6.356229, -6.210392, -6.064373, -5.918175, -5.771798, -5.625241, 
    -5.478507, -5.331595, -5.184507, -5.037242, -4.889802, -4.742187, 
    -4.594398, -4.446434, -4.298299, -4.149992, -4.001513, -3.852863, 
    -3.704043, -3.555054, -3.405896, -3.256571, -3.107079, -2.95742, 
    -2.807596, -2.657607, -2.507455, -2.357139, -2.206661, -2.056022, 
    -1.905222, -1.754262, -1.603143, -1.451866, -1.300432, -1.148842, 
    -0.9970958, -0.8451952, -0.6931409, -0.5409337, -0.3885746, -0.2360646, 
    -0.08340447, 0.06940477, 0.2223622, 0.3754668, 0.5287178, 0.6821139, 
    0.8356545, 0.9893383, 1.143165, 1.297132, 1.45124, 1.605487, 1.759873, 
    1.914395, 2.069054, 2.223848, 2.378776, 2.533837, 2.68903, 2.844354, 
    2.999808, 3.155391, 3.3111, 3.466937, 3.622899, 3.778985, 3.935194, 
    4.091525, 4.247976, 4.404548, 4.561238, 4.718045, 4.874968, 5.032006, 
    5.189157, 5.346422, 5.503798, 5.661283, 5.818878, 5.97658, 6.134388, 
    6.292302, 6.45032, 6.60844, 6.766662, 6.924983, 7.083404, 7.241922, 
    7.400536, 7.559246, 7.718049, 7.876944, 8.03593, 8.195006, 8.354171, 
    8.513422, 8.672759, 8.832181, 8.991686, 9.151272, 9.310939, 9.470684, 
    9.630507, 9.790406, 9.95038, 10.11043, 10.27055, 10.43074, 10.591, 
    10.75133, 10.91172, 11.07218, 11.2327, 11.39329, 11.55393, 11.71464, 
    11.8754, 12.03622, 12.19709, 12.35802, 12.519, 12.68003, 12.84111, 
    13.00224, 13.16341, 13.32463, 13.48589, 13.6472, 13.80854, 13.96993, 
    14.13135, 14.2928, 14.4543, 14.61582, 14.77738, 14.93896, 15.10058, 
    15.26222, 15.42389, 15.58558, 15.74729, 15.90902, 16.07078, 16.23255, 
    16.39434, 16.55614, 16.71796, 16.87979, 17.04163, 17.20348, 17.36533, 
    17.5272, 17.68906, 17.85093, 18.0128, 18.17467, 18.33654, 18.49841, 
    18.66027, 18.82212, 18.98397, 19.14581, 19.30764, 19.46945, 19.63125, 
    19.79304, 19.95481, 20.11656, 20.27829, 20.44, 20.60169, 20.76335, 
    20.92499, 21.0866, 21.24818, 21.40973, 21.57125, 21.73274, 21.89419, 
    22.0556, 22.21698, 22.37832, 22.53962, 22.70087, 22.86209, 23.02325, 
    23.18437, 23.34544, 23.50647, 23.66744, 23.82836, 23.98922, 24.15003, 
    24.31079, 24.47148, 24.63212, 24.7927, 24.95321, 25.11366, 25.27404, 
    25.43436, 25.59461, 25.75479, 25.91489, 26.07493, 26.23489, 26.39478, 
    26.55459, 26.71432, 26.87398, 27.03355, 27.19304, 27.35245, 27.51177, 
    27.67101, 27.83016, 27.98923, 28.1482, 28.30708, 28.46587, 28.62456, 
    28.78316, 28.94166, 29.10007, 29.25837, 29.41658, 29.57468, 29.73269, 
    29.89058, 30.04837, 30.20606, 30.36364, 30.5211, 30.67846, 30.83571, 
    30.99284, 31.14986, 31.30677, 31.46356, 31.62023, 31.77678, 31.93321, 
    32.08952, 32.24571, 32.40178, 32.55772, 32.71354, 32.86923, 33.02479, 
    33.18023, 33.33553, 33.4907, 33.64574, 33.80065, 33.95542, 34.11006, 
    34.26456, 34.41892, 34.57315, 34.72723, 34.88118, 35.03498, 35.18864, 
    35.34216, 35.49553, 35.64876, 35.80184, 35.95478, 36.10756, 36.2602, 
    36.41269, 36.56502, 36.71721, 36.86923, 37.02111, 37.17283, 37.3244, 
    37.47581, 37.62706, 37.77815, 37.92909, 38.07986, 38.23048, 38.38093, 
    38.53122, 38.68134, 38.83131, 38.98111, 39.13074, 39.2802, 39.4295, 
    39.57863, 39.7276, 39.87639, 40.02501, 40.17346, 40.32174, 40.46985, 
    40.61779, 40.76555, 40.91314, 41.06055, 41.20779, 41.35485, 41.50173, 
    41.64844, 41.79496, 41.94131, 42.08748, 42.23347, 42.37928, 42.52491, 
    42.67036, 42.81562, 42.9607, 43.1056, 43.25031, 43.39484, 43.53918, 
    43.68335, 43.82732, 43.9711, 44.1147, 44.25811, 44.40134, 44.54437,
  -21.03344, -20.90878, -20.78392, -20.65886, -20.5336, -20.40813, -20.28247, 
    -20.1566, -20.03053, -19.90425, -19.77777, -19.65109, -19.52421, 
    -19.39712, -19.26983, -19.14234, -19.01464, -18.88674, -18.75864, 
    -18.63033, -18.50183, -18.37311, -18.24419, -18.11507, -17.98575, 
    -17.85622, -17.72649, -17.59656, -17.46642, -17.33607, -17.20553, 
    -17.07478, -16.94382, -16.81266, -16.6813, -16.54974, -16.41797, 
    -16.28599, -16.15382, -16.02144, -15.88885, -15.75607, -15.62308, 
    -15.48988, -15.35649, -15.22289, -15.08909, -14.95508, -14.82087, 
    -14.68646, -14.55185, -14.41703, -14.28201, -14.14679, -14.01137, 
    -13.87575, -13.73992, -13.60389, -13.46766, -13.33123, -13.1946, 
    -13.05777, -12.92074, -12.78351, -12.64608, -12.50844, -12.37061, 
    -12.23258, -12.09435, -11.95592, -11.81729, -11.67847, -11.53944, 
    -11.40022, -11.2608, -11.12118, -10.98137, -10.84136, -10.70115, 
    -10.56075, -10.42015, -10.27936, -10.13837, -9.997186, -9.855809, 
    -9.714238, -9.572474, -9.430517, -9.288367, -9.146026, -9.003492, 
    -8.860767, -8.717852, -8.574745, -8.431449, -8.287963, -8.144288, 
    -8.000425, -7.856374, -7.712135, -7.567708, -7.423096, -7.278297, 
    -7.133313, -6.988143, -6.84279, -6.697252, -6.551531, -6.405627, 
    -6.259541, -6.113273, -5.966825, -5.820195, -5.673387, -5.526398, 
    -5.379232, -5.231887, -5.084365, -4.936667, -4.788793, -4.640743, 
    -4.492518, -4.344121, -4.195549, -4.046805, -3.89789, -3.748803, 
    -3.599546, -3.450119, -3.300524, -3.15076, -3.000829, -2.850732, 
    -2.700469, -2.550041, -2.399449, -2.248693, -2.097775, -1.946696, 
    -1.795455, -1.644055, -1.492495, -1.340777, -1.188902, -1.03687, 
    -0.8846824, -0.7323402, -0.5798441, -0.4271951, -0.2743941, -0.1214421, 
    0.03166004, 0.1849113, 0.3383109, 0.4918576, 0.6455507, 0.7993889, 
    0.9533716, 1.107497, 1.261766, 1.416175, 1.570725, 1.725414, 1.880241, 
    2.035205, 2.190305, 2.345541, 2.50091, 2.656412, 2.812046, 2.96781, 
    3.123704, 3.279727, 3.435877, 3.592153, 3.748554, 3.905079, 4.061727, 
    4.218496, 4.375386, 4.532395, 4.689522, 4.846766, 5.004126, 5.1616, 
    5.319188, 5.476887, 5.634697, 5.792618, 5.950646, 6.108782, 6.267024, 
    6.425369, 6.583819, 6.742371, 6.901023, 7.059775, 7.218625, 7.377572, 
    7.536615, 7.695752, 7.854982, 8.014303, 8.173716, 8.333217, 8.492805, 
    8.652481, 8.812241, 8.972084, 9.13201, 9.292017, 9.452104, 9.612268, 
    9.77251, 9.932826, 10.09322, 10.25368, 10.41421, 10.57482, 10.73549, 
    10.89623, 11.05704, 11.2179, 11.37884, 11.53983, 11.70088, 11.86199, 
    12.02316, 12.18438, 12.34566, 12.50699, 12.66837, 12.8298, 12.99128, 
    13.15281, 13.31438, 13.47599, 13.63765, 13.79934, 13.96108, 14.12285, 
    14.28466, 14.44651, 14.60839, 14.7703, 14.93224, 15.0942, 15.2562, 
    15.41822, 15.58027, 15.74234, 15.90443, 16.06654, 16.22866, 16.39081, 
    16.55297, 16.71514, 16.87733, 17.03952, 17.20173, 17.36394, 17.52616, 
    17.68838, 17.8506, 18.01283, 18.17506, 18.33728, 18.4995, 18.66172, 
    18.82393, 18.98614, 19.14833, 19.31051, 19.47268, 19.63484, 19.79698, 
    19.95911, 20.12122, 20.2833, 20.44537, 20.60741, 20.76943, 20.93142, 
    21.09338, 21.25532, 21.41722, 21.5791, 21.74094, 21.90274, 22.06451, 
    22.22624, 22.38793, 22.54958, 22.71119, 22.87275, 23.03427, 23.19574, 
    23.35716, 23.51853, 23.67985, 23.84112, 24.00234, 24.1635, 24.3246, 
    24.48564, 24.64663, 24.80755, 24.9684, 25.1292, 25.28993, 25.45059, 
    25.61119, 25.77171, 25.93216, 26.09254, 26.25284, 26.41307, 26.57323, 
    26.7333, 26.89329, 27.05321, 27.21304, 27.37278, 27.53244, 27.69202, 
    27.85151, 28.0109, 28.17021, 28.32943, 28.48855, 28.64758, 28.80651, 
    28.96534, 29.12408, 29.28272, 29.44125, 29.59969, 29.75801, 29.91624, 
    30.07436, 30.23237, 30.39027, 30.54807, 30.70575, 30.86332, 31.02077, 
    31.17812, 31.33534, 31.49245, 31.64944, 31.80631, 31.96306, 32.11969, 
    32.2762, 32.43258, 32.58883, 32.74496, 32.90096, 33.05684, 33.21258, 
    33.36819, 33.52368, 33.67902, 33.83424, 33.98932, 34.14426, 34.29906, 
    34.45373, 34.60826, 34.76265, 34.91689, 35.071, 35.22496, 35.37877, 
    35.53244, 35.68596, 35.83934, 35.99257, 36.14565, 36.29858, 36.45135, 
    36.60398, 36.75645, 36.90877, 37.06093, 37.21294, 37.36479, 37.51648, 
    37.66801, 37.81939, 37.9706, 38.12166, 38.27255, 38.42328, 38.57385, 
    38.72425, 38.87449, 39.02456, 39.17446, 39.3242, 39.47377, 39.62317, 
    39.7724, 39.92146, 40.07035, 40.21906, 40.36761, 40.51598, 40.66417, 
    40.81219, 40.96004, 41.10771, 41.25521, 41.40252, 41.54966, 41.69662, 
    41.8434, 41.99, 42.13642, 42.28266, 42.42872, 42.57459, 42.72029, 
    42.8658, 43.01112, 43.15626, 43.30122, 43.44598, 43.59057, 43.73496, 
    43.87917, 44.02319, 44.16703, 44.31067, 44.45413, 44.5974,
  -21.1034, -20.97861, -20.85361, -20.72841, -20.60302, -20.47741, -20.35161, 
    -20.2256, -20.09939, -19.97297, -19.84635, -19.71953, -19.5925, 
    -19.46527, -19.33783, -19.21019, -19.08235, -18.9543, -18.82605, 
    -18.69759, -18.56893, -18.44007, -18.311, -18.18172, -18.05224, 
    -17.92256, -17.79267, -17.66257, -17.53227, -17.40177, -17.27106, 
    -17.14015, -17.00903, -16.87771, -16.74618, -16.61445, -16.48251, 
    -16.35037, -16.21802, -16.08547, -15.95271, -15.81975, -15.68659, 
    -15.55322, -15.41965, -15.28587, -15.15189, -15.0177, -14.88332, 
    -14.74872, -14.61393, -14.47893, -14.34372, -14.20832, -14.07271, 
    -13.9369, -13.80088, -13.66466, -13.52824, -13.39162, -13.2548, 
    -13.11777, -12.98054, -12.84311, -12.70548, -12.56765, -12.42962, 
    -12.29138, -12.15295, -12.01432, -11.87549, -11.73645, -11.59722, 
    -11.45779, -11.31816, -11.17833, -11.03831, -10.89809, -10.75767, 
    -10.61705, -10.47623, -10.33522, -10.19402, -10.05261, -9.911016, 
    -9.769224, -9.627237, -9.485056, -9.342681, -9.200113, -9.057352, 
    -8.914399, -8.771254, -8.627916, -8.484388, -8.34067, -8.196761, 
    -8.052662, -7.908374, -7.763898, -7.619233, -7.47438, -7.329341, 
    -7.184114, -7.038702, -6.893104, -6.747321, -6.601353, -6.455202, 
    -6.308867, -6.162349, -6.015649, -5.868768, -5.721706, -5.574463, 
    -5.427041, -5.27944, -5.13166, -4.983703, -4.835569, -4.687258, 
    -4.538772, -4.39011, -4.241275, -4.092266, -3.943083, -3.793729, 
    -3.644203, -3.494507, -3.34464, -3.194605, -3.044401, -2.89403, 
    -2.743491, -2.592787, -2.441918, -2.290884, -2.139686, -1.988326, 
    -1.836804, -1.685121, -1.533278, -1.381275, -1.229114, -1.076796, 
    -0.9243203, -0.7716894, -0.6189035, -0.4659637, -0.3128709, -0.1596261, 
    -0.006230134, 0.147316, 0.3010113, 0.4548549, 0.6088457, 0.7629827, 
    0.9172651, 1.071692, 1.226261, 1.380974, 1.535827, 1.69082, 1.845953, 
    2.001223, 2.156631, 2.312174, 2.467853, 2.623665, 2.77961, 2.935686, 
    3.091893, 3.248229, 3.404693, 3.561285, 3.718002, 3.874844, 4.031809, 
    4.188898, 4.346107, 4.503437, 4.660885, 4.818451, 4.976134, 5.133932, 
    5.291843, 5.449869, 5.608005, 5.766252, 5.924608, 6.083072, 6.241642, 
    6.400318, 6.559098, 6.717981, 6.876966, 7.03605, 7.195233, 7.354515, 
    7.513892, 7.673365, 7.832931, 7.992589, 8.152338, 8.312178, 8.472105, 
    8.632119, 8.792219, 8.952403, 9.11267, 9.273019, 9.433447, 9.593954, 
    9.754539, 9.915199, 10.07593, 10.23674, 10.39762, 10.55857, 10.71959, 
    10.88068, 11.04183, 11.20305, 11.36433, 11.52567, 11.68707, 11.84853, 
    12.01005, 12.17162, 12.33325, 12.49493, 12.65666, 12.81844, 12.98028, 
    13.14215, 13.30408, 13.46604, 13.62805, 13.7901, 13.95219, 14.11432, 
    14.27649, 14.43869, 14.60092, 14.76318, 14.92548, 15.0878, 15.25016, 
    15.41253, 15.57494, 15.73736, 15.89981, 16.06227, 16.22476, 16.38726, 
    16.54978, 16.71231, 16.87485, 17.0374, 17.19997, 17.36254, 17.52511, 
    17.68769, 17.85028, 18.01286, 18.17544, 18.33803, 18.50061, 18.66318, 
    18.82575, 18.98831, 19.15086, 19.3134, 19.47593, 19.63844, 19.80094, 
    19.96342, 20.12589, 20.28833, 20.45075, 20.61315, 20.77553, 20.93787, 
    21.10019, 21.26249, 21.42475, 21.58697, 21.74917, 21.91133, 22.07345, 
    22.23553, 22.39758, 22.55958, 22.72154, 22.88346, 23.04533, 23.20715, 
    23.36893, 23.53065, 23.69232, 23.85394, 24.0155, 24.17701, 24.33846, 
    24.49986, 24.66119, 24.82246, 24.98367, 25.14481, 25.30588, 25.46689, 
    25.62783, 25.7887, 25.9495, 26.11022, 26.27087, 26.43144, 26.59194, 
    26.75235, 26.91269, 27.07294, 27.23311, 27.3932, 27.5532, 27.71311, 
    27.87294, 28.03267, 28.19232, 28.35187, 28.51133, 28.67069, 28.82995, 
    28.98912, 29.14819, 29.30716, 29.46602, 29.62479, 29.78345, 29.942, 
    30.10045, 30.25879, 30.41702, 30.57514, 30.73314, 30.89104, 31.04882, 
    31.20648, 31.36403, 31.52146, 31.67877, 31.83596, 31.99303, 32.14997, 
    32.3068, 32.46349, 32.62006, 32.77651, 32.93283, 33.08901, 33.24507, 
    33.40099, 33.55678, 33.71244, 33.86796, 34.02335, 34.1786, 34.33371, 
    34.48868, 34.64351, 34.7982, 34.95275, 35.10715, 35.26141, 35.41552, 
    35.56949, 35.72331, 35.87698, 36.03051, 36.18388, 36.3371, 36.49017, 
    36.64308, 36.79585, 36.94845, 37.1009, 37.25319, 37.40533, 37.55731, 
    37.70913, 37.86078, 38.01228, 38.16362, 38.31479, 38.46579, 38.61664, 
    38.76731, 38.91783, 39.06817, 39.21835, 39.36836, 39.5182, 39.66787, 
    39.81737, 39.96669, 40.11585, 40.26483, 40.41364, 40.56227, 40.71073, 
    40.85901, 41.00712, 41.15505, 41.3028, 41.45037, 41.59777, 41.74498, 
    41.89201, 42.03887, 42.18554, 42.33203, 42.47833, 42.62445, 42.77039, 
    42.91615, 43.06172, 43.2071, 43.35229, 43.49731, 43.64213, 43.78677, 
    43.93121, 44.07547, 44.21954, 44.36341, 44.50711, 44.6506,
  -21.17355, -21.04862, -20.92349, -20.79816, -20.67263, -20.54689, 
    -20.42094, -20.2948, -20.16844, -20.04189, -19.91513, -19.78816, 
    -19.66099, -19.53361, -19.40603, -19.27825, -19.15026, -19.02206, 
    -18.89366, -18.76505, -18.63624, -18.50722, -18.37799, -18.24856, 
    -18.11893, -17.98909, -17.85904, -17.72879, -17.59833, -17.46766, 
    -17.33679, -17.20572, -17.07444, -16.94295, -16.81125, -16.67936, 
    -16.54725, -16.41494, -16.28242, -16.1497, -16.01677, -15.88364, 
    -15.7503, -15.61676, -15.48301, -15.34905, -15.21489, -15.08053, 
    -14.94596, -14.81118, -14.6762, -14.54102, -14.40563, -14.27004, 
    -14.13424, -13.99824, -13.86204, -13.72563, -13.58902, -13.4522, 
    -13.31518, -13.17796, -13.04054, -12.90291, -12.76508, -12.62705, 
    -12.48882, -12.35038, -12.21175, -12.07291, -11.93387, -11.79463, 
    -11.65519, -11.51556, -11.37572, -11.23568, -11.09544, -10.95501, 
    -10.81437, -10.67354, -10.53251, -10.39128, -10.24985, -10.10823, 
    -9.966413, -9.824399, -9.682189, -9.539783, -9.397183, -9.254389, 
    -9.1114, -8.968218, -8.824842, -8.681274, -8.537514, -8.393561, 
    -8.249418, -8.105083, -7.960559, -7.815844, -7.67094, -7.525847, 
    -7.380566, -7.235097, -7.089441, -6.943598, -6.797569, -6.651354, 
    -6.504954, -6.35837, -6.211602, -6.064651, -5.917517, -5.770201, 
    -5.622704, -5.475025, -5.327167, -5.179129, -5.030912, -4.882517, 
    -4.733945, -4.585196, -4.43627, -4.287169, -4.137894, -3.988445, 
    -3.838822, -3.689027, -3.53906, -3.388922, -3.238614, -3.088136, 
    -2.93749, -2.786676, -2.635694, -2.484547, -2.333234, -2.181756, 
    -2.030115, -1.87831, -1.726344, -1.574216, -1.421928, -1.26948, 
    -1.116874, -0.9641103, -0.8111897, -0.6581131, -0.5048816, -0.3514961, 
    -0.1979575, -0.04426682, 0.1095751, 0.2635671, 0.4177084, 0.5719979, 
    0.7264347, 0.8810177, 1.035746, 1.190619, 1.345634, 1.500792, 1.656091, 
    1.81153, 1.967108, 2.122824, 2.278677, 2.434665, 2.590788, 2.747045, 
    2.903434, 3.059955, 3.216606, 3.373385, 3.530293, 3.687328, 3.844488, 
    4.001773, 4.159181, 4.316711, 4.474362, 4.632133, 4.790022, 4.948029, 
    5.106152, 5.26439, 5.422741, 5.581204, 5.739779, 5.898464, 6.057258, 
    6.216158, 6.375165, 6.534277, 6.693492, 6.85281, 7.012228, 7.171747, 
    7.331363, 7.491076, 7.650886, 7.810789, 7.970786, 8.130874, 8.291052, 
    8.451319, 8.611674, 8.772115, 8.932641, 9.09325, 9.253942, 9.414714, 
    9.575565, 9.736494, 9.8975, 10.05858, 10.21974, 10.38096, 10.54226, 
    10.70363, 10.86506, 11.02656, 11.18813, 11.34976, 11.51145, 11.6732, 
    11.83501, 11.99688, 12.15881, 12.32079, 12.48282, 12.64491, 12.80704, 
    12.96922, 13.13146, 13.29373, 13.45606, 13.61842, 13.78083, 13.94327, 
    14.10576, 14.26828, 14.43083, 14.59342, 14.75604, 14.9187, 15.08138, 
    15.24409, 15.40682, 15.56958, 15.73237, 15.89517, 16.058, 16.22084, 
    16.3837, 16.54658, 16.70946, 16.87237, 17.03528, 17.1982, 17.36113, 
    17.52406, 17.687, 17.84994, 18.01289, 18.17583, 18.33877, 18.50171, 
    18.66465, 18.82757, 18.99049, 19.1534, 19.3163, 19.47919, 19.64206, 
    19.80492, 19.96776, 20.13058, 20.29338, 20.45616, 20.61892, 20.78165, 
    20.94436, 21.10703, 21.26968, 21.4323, 21.59488, 21.75743, 21.91995, 
    22.08243, 22.24487, 22.40727, 22.56962, 22.73194, 22.89421, 23.05643, 
    23.21861, 23.38074, 23.54281, 23.70484, 23.86681, 24.02873, 24.19059, 
    24.35239, 24.51413, 24.67582, 24.83743, 24.99899, 25.16048, 25.32191, 
    25.48326, 25.64455, 25.80576, 25.96691, 26.12797, 26.28897, 26.44988, 
    26.61072, 26.77148, 26.93216, 27.09276, 27.25327, 27.4137, 27.57404, 
    27.73429, 27.89446, 28.05453, 28.21451, 28.3744, 28.53419, 28.69389, 
    28.85349, 29.01299, 29.1724, 29.3317, 29.4909, 29.64999, 29.80898, 
    29.96787, 30.12664, 30.28531, 30.44387, 30.60232, 30.76065, 30.91887, 
    31.07697, 31.23496, 31.39283, 31.55058, 31.70822, 31.86573, 32.02312, 
    32.18038, 32.33752, 32.49454, 32.65142, 32.80818, 32.96481, 33.12131, 
    33.27768, 33.43392, 33.59002, 33.74599, 33.90182, 34.05751, 34.21307, 
    34.36848, 34.52376, 34.6789, 34.83389, 34.98874, 35.14344, 35.298, 
    35.45242, 35.60669, 35.7608, 35.91477, 36.06859, 36.22226, 36.37577, 
    36.52913, 36.68234, 36.83539, 36.98829, 37.14103, 37.29361, 37.44603, 
    37.59829, 37.75039, 37.90233, 38.05411, 38.20573, 38.35718, 38.50847, 
    38.65959, 38.81054, 38.96133, 39.11195, 39.2624, 39.41268, 39.56279, 
    39.71273, 39.8625, 40.0121, 40.16152, 40.31077, 40.45984, 40.60874, 
    40.75746, 40.906, 41.05437, 41.20256, 41.35057, 41.4984, 41.64605, 
    41.79351, 41.9408, 42.08791, 42.23483, 42.38157, 42.52813, 42.6745, 
    42.82068, 42.96668, 43.1125, 43.25812, 43.40356, 43.54881, 43.69387, 
    43.83875, 43.98343, 44.12793, 44.27223, 44.41634, 44.56027, 44.704,
  -21.24389, -21.11884, -20.99357, -20.86811, -20.74244, -20.61656, 
    -20.49048, -20.36419, -20.2377, -20.111, -19.9841, -19.85699, -19.72968, 
    -19.60216, -19.47443, -19.3465, -19.21836, -19.09001, -18.96146, 
    -18.8327, -18.70374, -18.57457, -18.44519, -18.31561, -18.18582, 
    -18.05582, -17.92561, -17.7952, -17.66458, -17.53376, -17.40273, 
    -17.27149, -17.14004, -17.00839, -16.87653, -16.74446, -16.61219, 
    -16.47971, -16.34702, -16.21413, -16.08103, -15.94772, -15.81421, 
    -15.68049, -15.54656, -15.41243, -15.27809, -15.14355, -15.0088, 
    -14.87384, -14.73868, -14.60331, -14.46774, -14.33196, -14.19597, 
    -14.05978, -13.92339, -13.78679, -13.64999, -13.51298, -13.37577, 
    -13.23835, -13.10073, -12.96291, -12.82488, -12.68665, -12.54821, 
    -12.40958, -12.27074, -12.1317, -11.99245, -11.85301, -11.71336, 
    -11.57351, -11.43347, -11.29322, -11.15277, -11.01212, -10.87127, 
    -10.73022, -10.58897, -10.44753, -10.30588, -10.16404, -10.022, 
    -9.879765, -9.73733, -9.594701, -9.451875, -9.308853, -9.165636, 
    -9.022224, -8.878618, -8.734818, -8.590825, -8.446639, -8.30226, 
    -8.15769, -8.012928, -7.867975, -7.722831, -7.577498, -7.431975, 
    -7.286263, -7.140362, -6.994274, -6.847998, -6.701536, -6.554887, 
    -6.408053, -6.261034, -6.113831, -5.966443, -5.818872, -5.67112, 
    -5.523185, -5.375068, -5.226771, -5.078295, -4.929638, -4.780804, 
    -4.631791, -4.482601, -4.333235, -4.183692, -4.033975, -3.884083, 
    -3.734018, -3.58378, -3.43337, -3.282788, -3.132036, -2.981114, 
    -2.830023, -2.678764, -2.527337, -2.375744, -2.223986, -2.072062, 
    -1.919975, -1.767724, -1.615311, -1.462736, -1.310001, -1.157107, 
    -1.004053, -0.8508421, -0.697474, -0.5439499, -0.3902707, -0.2364375, 
    -0.08245112, 0.07168744, 0.2259772, 0.3804172, 0.5350064, 0.6897439, 
    0.8446286, 0.9996595, 1.154836, 1.310156, 1.465619, 1.621225, 1.776971, 
    1.932858, 2.088883, 2.245046, 2.401346, 2.557781, 2.714351, 2.871054, 
    3.02789, 3.184856, 3.341953, 3.499178, 3.656531, 3.814011, 3.971616, 
    4.129345, 4.287197, 4.445171, 4.603265, 4.761479, 4.919811, 5.07826, 
    5.236825, 5.395503, 5.554296, 5.7132, 5.872214, 6.031339, 6.190571, 
    6.34991, 6.509355, 6.668904, 6.828556, 6.988309, 7.148164, 7.308116, 
    7.468167, 7.628314, 7.788557, 7.948892, 8.109321, 8.269839, 8.430448, 
    8.591145, 8.751928, 8.912797, 9.07375, 9.234786, 9.395903, 9.557099, 
    9.718374, 9.879726, 10.04115, 10.20266, 10.36423, 10.52588, 10.68759, 
    10.84938, 11.01123, 11.17314, 11.33512, 11.49717, 11.65927, 11.82144, 
    11.98366, 12.14594, 12.30827, 12.47066, 12.6331, 12.79559, 12.95813, 
    13.12072, 13.28335, 13.44603, 13.60875, 13.77151, 13.93431, 14.09715, 
    14.26003, 14.42295, 14.58589, 14.74887, 14.91189, 15.07493, 15.238, 
    15.40109, 15.56421, 15.72735, 15.89052, 16.0537, 16.2169, 16.38012, 
    16.54336, 16.70661, 16.86987, 17.03314, 17.19642, 17.35971, 17.52301, 
    17.68631, 17.84961, 18.01292, 18.17622, 18.33952, 18.50282, 18.66612, 
    18.8294, 18.99269, 19.15596, 19.31922, 19.48246, 19.6457, 19.80891, 
    19.97211, 20.1353, 20.29846, 20.4616, 20.62471, 20.7878, 20.95087, 
    21.1139, 21.27691, 21.43988, 21.60283, 21.76574, 21.92861, 22.09144, 
    22.25424, 22.417, 22.57971, 22.74238, 22.90501, 23.06759, 23.23012, 
    23.3926, 23.55503, 23.71741, 23.87974, 24.04201, 24.20422, 24.36637, 
    24.52847, 24.6905, 24.85247, 25.01438, 25.17622, 25.33799, 25.4997, 
    25.66133, 25.8229, 25.98439, 26.1458, 26.30714, 26.4684, 26.62959, 
    26.79069, 26.95172, 27.11266, 27.27351, 27.43428, 27.59496, 27.75556, 
    27.91606, 28.07648, 28.2368, 28.39702, 28.55716, 28.71719, 28.87713, 
    29.03697, 29.1967, 29.35634, 29.51587, 29.6753, 29.83462, 29.99384, 
    30.15295, 30.31194, 30.47083, 30.6296, 30.78827, 30.94681, 31.10524, 
    31.26356, 31.42175, 31.57983, 31.73778, 31.89561, 32.05332, 32.21091, 
    32.36837, 32.5257, 32.68291, 32.83998, 32.99693, 33.15374, 33.31042, 
    33.46697, 33.62339, 33.77967, 33.93581, 34.09181, 34.24767, 34.4034, 
    34.55898, 34.71442, 34.86972, 35.02487, 35.17988, 35.33474, 35.48946, 
    35.64402, 35.79844, 35.95271, 36.10682, 36.26078, 36.41459, 36.56824, 
    36.72174, 36.87509, 37.02827, 37.1813, 37.33417, 37.48688, 37.63943, 
    37.79182, 37.94404, 38.0961, 38.248, 38.39973, 38.5513, 38.7027, 
    38.85394, 39.005, 39.1559, 39.30662, 39.45717, 39.60756, 39.75777, 
    39.90781, 40.05767, 40.20736, 40.35687, 40.50621, 40.65537, 40.80436, 
    40.95317, 41.10179, 41.25024, 41.39851, 41.5466, 41.6945, 41.84223, 
    41.98977, 42.13713, 42.2843, 42.43129, 42.5781, 42.72472, 42.87115, 
    43.0174, 43.16345, 43.30933, 43.45501, 43.6005, 43.7458, 43.89092, 
    44.03584, 44.18057, 44.32511, 44.46946, 44.61362, 44.75758,
  -21.31444, -21.18925, -21.06385, -20.93825, -20.81244, -20.68643, 
    -20.56021, -20.43379, -20.30716, -20.18032, -20.05327, -19.92602, 
    -19.79856, -19.6709, -19.54303, -19.41495, -19.28666, -19.15817, 
    -19.02947, -18.90056, -18.77144, -18.64212, -18.51259, -18.38285, 
    -18.2529, -18.12275, -17.99239, -17.86182, -17.73104, -17.60005, 
    -17.46886, -17.33746, -17.20585, -17.07403, -16.94201, -16.80977, 
    -16.67733, -16.54468, -16.41183, -16.27876, -16.14549, -16.01201, 
    -15.87832, -15.74443, -15.61032, -15.47601, -15.3415, -15.20677, 
    -15.07184, -14.9367, -14.80136, -14.6658, -14.53004, -14.39408, 
    -14.25791, -14.12153, -13.98494, -13.84815, -13.71116, -13.57396, 
    -13.43655, -13.29894, -13.16112, -13.0231, -12.88487, -12.74644, 
    -12.60781, -12.46897, -12.32993, -12.19068, -12.05123, -11.91158, 
    -11.77173, -11.63167, -11.49141, -11.35095, -11.21029, -11.06943, 
    -10.92836, -10.7871, -10.64563, -10.50397, -10.36211, -10.22004, 
    -10.07778, -9.935322, -9.792664, -9.649809, -9.506756, -9.363507, 
    -9.220061, -9.07642, -8.932584, -8.788551, -8.644325, -8.499905, 
    -8.35529, -8.210484, -8.065484, -7.920291, -7.774908, -7.629333, 
    -7.483567, -7.337612, -7.191467, -7.045133, -6.89861, -6.751899, 
    -6.605001, -6.457917, -6.310646, -6.163189, -6.015548, -5.867723, 
    -5.719713, -5.571521, -5.423146, -5.27459, -5.125852, -4.976934, 
    -4.827837, -4.678559, -4.529104, -4.379471, -4.229661, -4.079676, 
    -3.929514, -3.779178, -3.628668, -3.477984, -3.327129, -3.176101, 
    -3.024903, -2.873534, -2.721997, -2.570291, -2.418417, -2.266376, 
    -2.11417, -1.961798, -1.809262, -1.656563, -1.503702, -1.350678, 
    -1.197494, -1.04415, -0.8906479, -0.7369873, -0.5831696, -0.429196, 
    -0.2750672, -0.1207842, 0.03365204, 0.1882405, 0.3429801, 0.49787, 
    0.6529092, 0.8080965, 0.9634311, 1.118912, 1.274538, 1.430308, 1.586221, 
    1.742276, 1.898472, 2.054807, 2.211282, 2.367894, 2.524642, 2.681526, 
    2.838545, 2.995696, 3.15298, 3.310394, 3.467938, 3.625611, 3.783411, 
    3.941337, 4.099389, 4.257564, 4.415862, 4.574281, 4.73282, 4.891479, 
    5.050254, 5.209147, 5.368155, 5.527277, 5.686512, 5.845858, 6.005313, 
    6.164879, 6.324552, 6.484331, 6.644215, 6.804203, 6.964293, 7.124484, 
    7.284775, 7.445164, 7.60565, 7.766232, 7.926908, 8.087678, 8.248539, 
    8.40949, 8.57053, 8.731657, 8.892871, 9.054169, 9.21555, 9.377013, 
    9.538557, 9.70018, 9.861879, 10.02366, 10.18551, 10.34743, 10.50943, 
    10.67149, 10.83363, 10.99583, 11.1581, 11.32043, 11.48283, 11.64529, 
    11.80781, 11.97038, 12.13301, 12.2957, 12.45845, 12.62124, 12.78409, 
    12.94698, 13.10993, 13.27292, 13.43595, 13.59903, 13.76215, 13.92532, 
    14.08852, 14.25175, 14.41503, 14.57833, 14.74167, 14.90505, 15.06845, 
    15.23188, 15.39533, 15.55881, 15.72231, 15.88584, 16.04939, 16.21295, 
    16.37653, 16.54013, 16.70374, 16.86736, 17.031, 17.19464, 17.35829, 
    17.52195, 17.68561, 17.84928, 18.01295, 18.17661, 18.34028, 18.50394, 
    18.66759, 18.83125, 18.99489, 19.15852, 19.32214, 19.48575, 19.64935, 
    19.81292, 19.97649, 20.14003, 20.30355, 20.46705, 20.63053, 20.79398, 
    20.9574, 21.1208, 21.28417, 21.4475, 21.6108, 21.77407, 21.9373, 22.1005, 
    22.26365, 22.42677, 22.58984, 22.75287, 22.91585, 23.07879, 23.24167, 
    23.40451, 23.5673, 23.73004, 23.89272, 24.05534, 24.21791, 24.38041, 
    24.54286, 24.70525, 24.86757, 25.02983, 25.19202, 25.35415, 25.5162, 
    25.67819, 25.8401, 26.00194, 26.1637, 26.32539, 26.487, 26.64853, 
    26.80998, 26.97135, 27.13264, 27.29384, 27.45495, 27.61598, 27.77691, 
    27.93776, 28.09851, 28.25918, 28.41974, 28.58021, 28.74059, 28.90086, 
    29.06104, 29.22111, 29.38108, 29.54095, 29.70071, 29.86037, 30.01992, 
    30.17936, 30.33868, 30.4979, 30.65701, 30.81599, 30.97487, 31.13363, 
    31.29227, 31.45079, 31.60919, 31.76747, 31.92562, 32.08365, 32.24156, 
    32.39934, 32.55699, 32.71452, 32.87191, 33.02917, 33.1863, 33.3433, 
    33.50016, 33.65689, 33.81348, 33.96993, 34.12624, 34.28242, 34.43845, 
    34.59434, 34.75009, 34.90569, 35.06115, 35.21646, 35.37162, 35.52664, 
    35.68151, 35.83622, 35.99079, 36.1452, 36.29946, 36.45356, 36.60751, 
    36.7613, 36.91494, 37.06842, 37.22174, 37.37489, 37.52789, 37.68073, 
    37.8334, 37.98591, 38.13826, 38.29044, 38.44245, 38.5943, 38.74598, 
    38.89749, 39.04883, 39.2, 39.351, 39.50183, 39.65249, 39.80297, 39.95328, 
    40.10341, 40.25337, 40.40315, 40.55276, 40.70218, 40.85143, 41.0005, 
    41.14939, 41.2981, 41.44663, 41.59497, 41.74314, 41.89112, 42.03891, 
    42.18653, 42.33395, 42.4812, 42.62825, 42.77512, 42.9218, 43.06829, 
    43.2146, 43.36071, 43.50664, 43.65237, 43.79792, 43.94327, 44.08843, 
    44.2334, 44.37818, 44.52276, 44.66715, 44.81135,
  -21.38518, -21.25986, -21.13433, -21.00859, -20.88265, -20.7565, -20.63014, 
    -20.50358, -20.37681, -20.24983, -20.12265, -19.99525, -19.86765, 
    -19.73984, -19.61182, -19.4836, -19.35517, -19.22652, -19.09767, 
    -18.96861, -18.83935, -18.70987, -18.58019, -18.45029, -18.32019, 
    -18.18988, -18.05936, -17.92863, -17.7977, -17.66655, -17.53519, 
    -17.40363, -17.27186, -17.13987, -17.00768, -16.87528, -16.74267, 
    -16.60986, -16.47683, -16.34359, -16.21015, -16.07649, -15.94263, 
    -15.80856, -15.67428, -15.53979, -15.4051, -15.27019, -15.13508, 
    -14.99976, -14.86423, -14.7285, -14.59255, -14.4564, -14.32004, 
    -14.18347, -14.0467, -13.90972, -13.77253, -13.63513, -13.49753, 
    -13.35973, -13.22171, -13.08349, -12.94507, -12.80644, -12.6676, 
    -12.52856, -12.38931, -12.24986, -12.11021, -11.97035, -11.83029, 
    -11.69002, -11.54955, -11.40888, -11.26801, -11.12693, -10.98565, 
    -10.84417, -10.70249, -10.56061, -10.41852, -10.27624, -10.13375, 
    -9.991072, -9.848189, -9.705109, -9.56183, -9.418353, -9.274678, 
    -9.130807, -8.986739, -8.842475, -8.698014, -8.553359, -8.408509, 
    -8.263465, -8.118227, -7.972795, -7.827171, -7.681354, -7.535346, 
    -7.389146, -7.242755, -7.096175, -6.949405, -6.802445, -6.655297, 
    -6.507962, -6.360439, -6.212729, -6.064833, -5.916752, -5.768486, 
    -5.620036, -5.471402, -5.322585, -5.173586, -5.024405, -4.875044, 
    -4.725502, -4.575781, -4.425881, -4.275803, -4.125548, -3.975116, 
    -3.824508, -3.673725, -3.522768, -3.371637, -3.220334, -3.068858, 
    -2.917211, -2.765394, -2.613408, -2.461252, -2.308929, -2.156439, 
    -2.003783, -1.850961, -1.697975, -1.544825, -1.391512, -1.238038, 
    -1.084403, -0.9306082, -0.7766541, -0.6225421, -0.4682729, -0.3138476, 
    -0.159267, -0.004532254, 0.1503558, 0.3053961, 0.4605876, 0.6159294, 
    0.7714204, 0.9270597, 1.082846, 1.238779, 1.394856, 1.551078, 1.707442, 
    1.863949, 2.020596, 2.177383, 2.334308, 2.491371, 2.648571, 2.805905, 
    2.963374, 3.120975, 3.278709, 3.436573, 3.594566, 3.752688, 3.910937, 
    4.069311, 4.22781, 4.386434, 4.545178, 4.704045, 4.86303, 5.022135, 
    5.181357, 5.340695, 5.500148, 5.659714, 5.819393, 5.979182, 6.139081, 
    6.299089, 6.459203, 6.619424, 6.779748, 6.940176, 7.100706, 7.261336, 
    7.422066, 7.582892, 7.743816, 7.904834, 8.065946, 8.22715, 8.388445, 
    8.549829, 8.711303, 8.872862, 9.034507, 9.196235, 9.358046, 9.519938, 
    9.681909, 9.843958, 10.00608, 10.16829, 10.33056, 10.49291, 10.65533, 
    10.81781, 10.98037, 11.14299, 11.30568, 11.46843, 11.63124, 11.79412, 
    11.95705, 12.12004, 12.28308, 12.44618, 12.60933, 12.77254, 12.93579, 
    13.0991, 13.26245, 13.42584, 13.58928, 13.75276, 13.91628, 14.07984, 
    14.24344, 14.40707, 14.57074, 14.73444, 14.89818, 15.06194, 15.22573, 
    15.38955, 15.55339, 15.71726, 15.88114, 16.04505, 16.20898, 16.37292, 
    16.53688, 16.70086, 16.86485, 17.02884, 17.19285, 17.35687, 17.52089, 
    17.68491, 17.84894, 18.01297, 18.177, 18.34103, 18.50506, 18.66908, 
    18.83309, 18.9971, 19.16109, 19.32508, 19.48905, 19.65301, 19.81695, 
    19.98088, 20.14478, 20.30867, 20.47253, 20.63637, 20.80018, 20.96397, 
    21.12773, 21.29145, 21.45515, 21.61881, 21.78244, 21.94603, 22.10959, 
    22.2731, 22.43658, 22.60001, 22.7634, 22.92674, 23.09003, 23.25328, 
    23.41648, 23.57962, 23.74271, 23.90575, 24.06873, 24.23165, 24.39452, 
    24.55732, 24.72006, 24.88274, 25.04535, 25.20789, 25.37037, 25.53278, 
    25.69511, 25.85738, 26.01957, 26.18168, 26.34372, 26.50568, 26.66755, 
    26.82935, 26.99107, 27.1527, 27.31425, 27.4757, 27.63708, 27.79836, 
    27.95955, 28.12064, 28.28165, 28.44255, 28.60336, 28.76408, 28.92469, 
    29.08521, 29.24562, 29.40593, 29.56613, 29.72623, 29.88622, 30.0461, 
    30.20587, 30.36553, 30.52508, 30.68452, 30.84384, 31.00304, 31.16213, 
    31.32109, 31.47994, 31.63867, 31.79727, 31.95575, 32.11411, 32.27233, 
    32.43044, 32.58841, 32.74625, 32.90396, 33.06154, 33.21899, 33.3763, 
    33.53348, 33.69053, 33.84743, 34.00419, 34.16082, 34.3173, 34.47364, 
    34.62984, 34.7859, 34.94181, 35.09757, 35.25319, 35.40865, 35.56397, 
    35.71914, 35.87416, 36.02902, 36.18373, 36.33829, 36.49269, 36.64693, 
    36.80102, 36.95495, 37.10872, 37.26233, 37.41578, 37.56906, 37.72219, 
    37.87514, 38.02794, 38.18057, 38.33303, 38.48533, 38.63746, 38.78942, 
    38.94121, 39.09283, 39.24428, 39.39555, 39.54666, 39.69759, 39.84834, 
    39.99892, 40.14933, 40.29956, 40.4496, 40.59948, 40.74917, 40.89868, 
    41.04802, 41.19717, 41.34614, 41.49493, 41.64353, 41.79195, 41.94019, 
    42.08824, 42.23611, 42.38379, 42.53128, 42.67859, 42.8257, 42.97263, 
    43.11937, 43.26593, 43.41228, 43.55846, 43.70443, 43.85022, 43.99581, 
    44.14121, 44.28642, 44.43143, 44.57626, 44.72088, 44.86531,
  -21.45613, -21.33067, -21.20501, -21.07914, -20.95306, -20.82677, 
    -20.70028, -20.57358, -20.44667, -20.31955, -20.19222, -20.06469, 
    -19.93694, -19.80899, -19.68082, -19.55245, -19.42387, -19.29508, 
    -19.16608, -19.03687, -18.90746, -18.77783, -18.64799, -18.51794, 
    -18.38769, -18.25722, -18.12654, -17.99565, -17.86456, -17.73325, 
    -17.60173, -17.47001, -17.33807, -17.20592, -17.07356, -16.941, 
    -16.80822, -16.67523, -16.54204, -16.40863, -16.27501, -16.14118, 
    -16.00715, -15.8729, -15.73845, -15.60378, -15.4689, -15.33382, 
    -15.19853, -15.06302, -14.92731, -14.79139, -14.65526, -14.51892, 
    -14.38237, -14.24562, -14.10865, -13.97148, -13.8341, -13.69651, 
    -13.55872, -13.42071, -13.2825, -13.14409, -13.00546, -12.86663, 
    -12.72759, -12.58835, -12.4489, -12.30924, -12.16938, -12.02932, 
    -11.88905, -11.74857, -11.60789, -11.46701, -11.32592, -11.18463, 
    -11.04313, -10.90144, -10.75954, -10.61744, -10.47513, -10.33263, 
    -10.18992, -10.04702, -9.90391, -9.760603, -9.617097, -9.473392, 
    -9.329488, -9.185386, -9.041086, -8.896588, -8.751895, -8.607004, 
    -8.461918, -8.316636, -8.171159, -8.025487, -7.879622, -7.733563, 
    -7.587311, -7.440866, -7.29423, -7.147403, -7.000384, -6.853176, 
    -6.705777, -6.55819, -6.410414, -6.262451, -6.1143, -5.965962, -5.817439, 
    -5.66873, -5.519836, -5.370758, -5.221497, -5.072053, -4.922428, 
    -4.77262, -4.622633, -4.472465, -4.322118, -4.171593, -4.020889, 
    -3.870009, -3.718953, -3.567721, -3.416315, -3.264734, -3.112981, 
    -2.961055, -2.808958, -2.65669, -2.504252, -2.351645, -2.198871, 
    -2.045928, -1.89282, -1.739546, -1.586107, -1.432505, -1.278739, 
    -1.124812, -0.970724, -0.8164757, -0.6620683, -0.5075027, -0.3527799, 
    -0.1979009, -0.04286657, 0.112322, 0.2676639, 0.4231581, 0.5788035, 
    0.7345992, 0.8905441, 1.046637, 1.202877, 1.359264, 1.515795, 1.67247, 
    1.829288, 1.986248, 2.143348, 2.300588, 2.457967, 2.615482, 2.773134, 
    2.930921, 3.088842, 3.246895, 3.40508, 3.563395, 3.72184, 3.880412, 
    4.039112, 4.197936, 4.356885, 4.515958, 4.675152, 4.834467, 4.993901, 
    5.153453, 5.313123, 5.472908, 5.632807, 5.792819, 5.952943, 6.113177, 
    6.273521, 6.433972, 6.594531, 6.755194, 6.915961, 7.07683, 7.237801, 
    7.398871, 7.56004, 7.721306, 7.882668, 8.044124, 8.205672, 8.367313, 
    8.529043, 8.690863, 8.852769, 9.014762, 9.176838, 9.338998, 9.50124, 
    9.663561, 9.825961, 9.988439, 10.15099, 10.31362, 10.47632, 10.63909, 
    10.80193, 10.96484, 11.12782, 11.29086, 11.45397, 11.61714, 11.78037, 
    11.94366, 12.10701, 12.27041, 12.43387, 12.59738, 12.76094, 12.92456, 
    13.08822, 13.25193, 13.41568, 13.57948, 13.74332, 13.90721, 14.07113, 
    14.23509, 14.39909, 14.56312, 14.72718, 14.89128, 15.0554, 15.21956, 
    15.38374, 15.54795, 15.71218, 15.87643, 16.0407, 16.20499, 16.3693, 
    16.53363, 16.69797, 16.86232, 17.02668, 17.19106, 17.35543, 17.51982, 
    17.68421, 17.84861, 18.013, 18.1774, 18.34179, 18.50618, 18.67057, 
    18.83495, 18.99932, 19.16368, 19.32803, 19.49237, 19.65669, 19.821, 
    19.98528, 20.14956, 20.3138, 20.47803, 20.64223, 20.80641, 20.97056, 
    21.13468, 21.29877, 21.46283, 21.62686, 21.79085, 21.9548, 22.11872, 
    22.2826, 22.44643, 22.61022, 22.77397, 22.93767, 23.10133, 23.26493, 
    23.42849, 23.59199, 23.75544, 23.91884, 24.08218, 24.24545, 24.40868, 
    24.57183, 24.73493, 24.89796, 25.06093, 25.22383, 25.38666, 25.54942, 
    25.71211, 25.87473, 26.03727, 26.19973, 26.36212, 26.52443, 26.68666, 
    26.8488, 27.01087, 27.17285, 27.33474, 27.49655, 27.65826, 27.81989, 
    27.98142, 28.14286, 28.30421, 28.46546, 28.62661, 28.78767, 28.94862, 
    29.10948, 29.27023, 29.43087, 29.59142, 29.75185, 29.91218, 30.07239, 
    30.2325, 30.39249, 30.55238, 30.71214, 30.87179, 31.03133, 31.19074, 
    31.35004, 31.50921, 31.66827, 31.8272, 31.986, 32.14468, 32.30323, 
    32.46165, 32.61995, 32.77811, 32.93615, 33.09405, 33.25181, 33.40944, 
    33.56694, 33.72429, 33.88151, 34.03859, 34.19553, 34.35232, 34.50898, 
    34.66549, 34.82185, 34.97807, 35.13413, 35.29005, 35.44583, 35.60145, 
    35.75692, 35.91224, 36.0674, 36.22241, 36.37727, 36.53196, 36.6865, 
    36.84089, 36.99511, 37.14917, 37.30307, 37.45681, 37.61039, 37.7638, 
    37.91705, 38.07013, 38.22305, 38.3758, 38.52838, 38.68079, 38.83303, 
    38.9851, 39.137, 39.28872, 39.44028, 39.59166, 39.74286, 39.89389, 
    40.04474, 40.19542, 40.34591, 40.49623, 40.64637, 40.79633, 40.94611, 
    41.09571, 41.24512, 41.39435, 41.5434, 41.69226, 41.84095, 41.98944, 
    42.13775, 42.28587, 42.4338, 42.58155, 42.72911, 42.87647, 43.02365, 
    43.17064, 43.31744, 43.46404, 43.61046, 43.75668, 43.90271, 44.04854, 
    44.19418, 44.33963, 44.48488, 44.62994, 44.7748, 44.91946,
  -21.52727, -21.40168, -21.27589, -21.14988, -21.02367, -20.89725, 
    -20.77061, -20.64378, -20.51673, -20.38947, -20.262, -20.13432, 
    -20.00643, -19.87834, -19.75003, -19.62151, -19.49278, -19.36385, 
    -19.2347, -19.10534, -18.97577, -18.84599, -18.716, -18.58579, -18.45538, 
    -18.32476, -18.19392, -18.06288, -17.93162, -17.80015, -17.66848, 
    -17.53659, -17.40449, -17.27217, -17.13965, -17.00692, -16.87397, 
    -16.74081, -16.60745, -16.47387, -16.34008, -16.20608, -16.07187, 
    -15.93745, -15.80281, -15.66797, -15.53292, -15.39765, -15.26218, 
    -15.12649, -14.99059, -14.85449, -14.71817, -14.58165, -14.44491, 
    -14.30797, -14.17081, -14.03345, -13.89588, -13.75809, -13.6201, 
    -13.4819, -13.3435, -13.20488, -13.06606, -12.92702, -12.78779, 
    -12.64834, -12.50869, -12.36883, -12.22876, -12.08848, -11.94801, 
    -11.80732, -11.66643, -11.52533, -11.38403, -11.24253, -11.10082, 
    -10.9589, -10.81679, -10.67447, -10.53194, -10.38921, -10.24629, 
    -10.10316, -9.959825, -9.816292, -9.672558, -9.528625, -9.384491, 
    -9.240158, -9.095626, -8.950895, -8.805966, -8.66084, -8.515517, 
    -8.369997, -8.22428, -8.078369, -7.932262, -7.78596, -7.639464, 
    -7.492774, -7.345892, -7.198817, -7.05155, -6.904091, -6.756442, 
    -6.608603, -6.460573, -6.312355, -6.163949, -6.015354, -5.866572, 
    -5.717604, -5.56845, -5.419111, -5.269587, -5.11988, -4.969989, 
    -4.819915, -4.66966, -4.519224, -4.368608, -4.217811, -4.066836, 
    -3.915683, -3.764352, -3.612845, -3.461162, -3.309304, -3.157272, 
    -3.005067, -2.852688, -2.700138, -2.547417, -2.394526, -2.241466, 
    -2.088238, -1.934841, -1.781278, -1.62755, -1.473657, -1.319599, 
    -1.165379, -1.010997, -0.8564532, -0.7017495, -0.5468866, -0.3918654, 
    -0.2366869, -0.08135205, 0.0741381, 0.2297826, 0.3855804, 0.5415304, 
    0.6976318, 0.8538834, 1.010284, 1.166833, 1.323529, 1.480371, 1.637358, 
    1.794488, 1.951762, 2.109177, 2.266732, 2.424427, 2.582261, 2.740231, 
    2.898337, 3.056578, 3.214953, 3.37346, 3.532098, 3.690866, 3.849764, 
    4.008789, 4.16794, 4.327217, 4.486618, 4.646141, 4.805786, 4.965551, 
    5.125435, 5.285437, 5.445555, 5.605788, 5.766136, 5.926596, 6.087167, 
    6.247848, 6.408637, 6.569534, 6.730537, 6.891644, 7.052855, 7.214168, 
    7.37558, 7.537093, 7.698702, 7.860409, 8.02221, 8.184105, 8.346092, 
    8.50817, 8.670337, 8.832592, 8.994934, 9.15736, 9.319871, 9.482463, 
    9.645137, 9.807889, 9.970719, 10.13363, 10.29661, 10.45966, 10.62279, 
    10.78599, 10.94925, 11.11259, 11.27598, 11.43945, 11.60298, 11.76656, 
    11.93021, 12.09392, 12.25768, 12.4215, 12.58537, 12.7493, 12.91327, 
    13.07729, 13.24136, 13.40548, 13.56964, 13.73385, 13.89809, 14.06238, 
    14.2267, 14.39106, 14.55546, 14.71989, 14.88435, 15.04884, 15.21336, 
    15.37791, 15.54248, 15.70707, 15.87169, 16.03633, 16.20099, 16.36567, 
    16.53036, 16.69506, 16.85978, 17.02451, 17.18925, 17.354, 17.51875, 
    17.68351, 17.84827, 18.01303, 18.17779, 18.34255, 18.50731, 18.67206, 
    18.83681, 19.00155, 19.16628, 19.33099, 19.4957, 19.66039, 19.82506, 
    19.98971, 20.15435, 20.31896, 20.48356, 20.64812, 20.81267, 20.97718, 
    21.14167, 21.30612, 21.47055, 21.63494, 21.79929, 21.96361, 22.12789, 
    22.29213, 22.45633, 22.62048, 22.78459, 22.94866, 23.11267, 23.27664, 
    23.44056, 23.60442, 23.76823, 23.93198, 24.09568, 24.25932, 24.4229, 
    24.58641, 24.74987, 24.91326, 25.07658, 25.23983, 25.40302, 25.56614, 
    25.72918, 25.89215, 26.05504, 26.21786, 26.3806, 26.54326, 26.70584, 
    26.86834, 27.03075, 27.19308, 27.35532, 27.51748, 27.67954, 27.84151, 
    28.00339, 28.16518, 28.32687, 28.48846, 28.64996, 28.81136, 28.97265, 
    29.13385, 29.29494, 29.45592, 29.6168, 29.77758, 29.93824, 30.09879, 
    30.25924, 30.41957, 30.57978, 30.73988, 30.89986, 31.05973, 31.21947, 
    31.3791, 31.5386, 31.69799, 31.85724, 32.01638, 32.17538, 32.33426, 
    32.493, 32.65162, 32.81011, 32.96846, 33.12668, 33.28477, 33.44271, 
    33.60052, 33.7582, 33.91573, 34.07312, 34.23038, 34.38749, 34.54445, 
    34.70127, 34.85794, 35.01447, 35.17084, 35.32707, 35.48315, 35.63908, 
    35.79485, 35.95047, 36.10593, 36.26125, 36.4164, 36.5714, 36.72623, 
    36.88091, 37.03543, 37.18979, 37.34398, 37.49801, 37.65188, 37.80558, 
    37.95912, 38.11249, 38.26569, 38.41872, 38.57159, 38.72428, 38.8768, 
    39.02916, 39.18133, 39.33334, 39.48517, 39.63682, 39.7883, 39.93961, 
    40.09073, 40.24168, 40.39244, 40.54303, 40.69344, 40.84367, 40.99371, 
    41.14357, 41.29325, 41.44275, 41.59206, 41.74118, 41.89012, 42.03887, 
    42.18744, 42.33581, 42.484, 42.632, 42.77981, 42.92743, 43.07486, 
    43.2221, 43.36914, 43.51599, 43.66265, 43.80912, 43.95539, 44.10146, 
    44.24734, 44.39303, 44.53852, 44.68381, 44.82891, 44.9738,
  -21.59862, -21.4729, -21.34697, -21.22083, -21.09448, -20.96792, -20.84116, 
    -20.71418, -20.58699, -20.45959, -20.33198, -20.20416, -20.07613, 
    -19.94789, -19.81944, -19.69077, -19.5619, -19.43281, -19.30351, 
    -19.17401, -19.04428, -18.91435, -18.78421, -18.65385, -18.52328, 
    -18.3925, -18.26151, -18.13031, -17.99889, -17.86726, -17.73542, 
    -17.60337, -17.47111, -17.33863, -17.20594, -17.07304, -16.93993, 
    -16.8066, -16.67306, -16.53931, -16.40535, -16.27118, -16.13679, 
    -16.0022, -15.86739, -15.73236, -15.59713, -15.46169, -15.32603, 
    -15.19016, -15.05408, -14.91779, -14.78129, -14.64458, -14.50765, 
    -14.37052, -14.23318, -14.09562, -13.95785, -13.81988, -13.68169, 
    -13.5433, -13.40469, -13.26588, -13.12686, -12.98762, -12.84818, 
    -12.70853, -12.56868, -12.42861, -12.28833, -12.14785, -12.00717, 
    -11.86627, -11.72517, -11.58386, -11.44234, -11.30062, -11.1587, 
    -11.01657, -10.87423, -10.73169, -10.58895, -10.446, -10.30285, 
    -10.15949, -10.01594, -9.872176, -9.728215, -9.584052, -9.439689, 
    -9.295124, -9.15036, -9.005396, -8.860232, -8.714869, -8.569309, 
    -8.423551, -8.277595, -8.131441, -7.985092, -7.838547, -7.691807, 
    -7.544872, -7.397742, -7.250419, -7.102903, -6.955194, -6.807293, 
    -6.659201, -6.510918, -6.362444, -6.213781, -6.064929, -5.915889, 
    -5.766661, -5.617246, -5.467645, -5.317857, -5.167885, -5.017729, 
    -4.867388, -4.716865, -4.56616, -4.415273, -4.264205, -4.112957, 
    -3.96153, -3.809925, -3.658142, -3.506181, -3.354045, -3.201734, 
    -3.049247, -2.896587, -2.743754, -2.590749, -2.437573, -2.284227, 
    -2.130711, -1.977026, -1.823174, -1.669154, -1.514969, -1.360619, 
    -1.206105, -1.051427, -0.8965877, -0.7415868, -0.5864256, -0.431105, 
    -0.2756261, -0.1199898, 0.03580284, 0.1917509, 0.3478533, 0.504109, 
    0.660517, 0.8170763, 0.9737858, 1.130644, 1.287651, 1.444805, 1.602104, 
    1.759549, 1.917137, 2.074868, 2.23274, 2.390753, 2.548904, 2.707194, 
    2.865621, 3.024183, 3.18288, 3.341711, 3.500673, 3.659767, 3.81899, 
    3.978342, 4.137821, 4.297426, 4.457157, 4.617011, 4.776987, 4.937084, 
    5.097301, 5.257637, 5.418089, 5.578659, 5.739342, 5.900139, 6.061048, 
    6.222067, 6.383197, 6.544434, 6.705778, 6.867227, 7.02878, 7.190435, 
    7.352192, 7.514049, 7.676004, 7.838057, 8.000205, 8.162447, 8.324782, 
    8.487208, 8.649725, 8.81233, 8.975022, 9.1378, 9.300663, 9.463608, 
    9.626634, 9.78974, 9.952925, 10.11619, 10.27952, 10.44293, 10.60642, 
    10.76997, 10.93359, 11.09729, 11.26104, 11.42487, 11.58875, 11.7527, 
    11.91671, 12.08077, 12.2449, 12.40908, 12.57331, 12.7376, 12.90194, 
    13.06632, 13.23076, 13.39524, 13.55976, 13.72433, 13.88894, 14.05359, 
    14.21828, 14.38301, 14.54777, 14.71256, 14.87739, 15.04225, 15.20713, 
    15.37205, 15.53699, 15.70195, 15.86694, 16.03194, 16.19697, 16.36201, 
    16.52707, 16.69214, 16.85723, 17.02233, 17.18744, 17.35255, 17.51767, 
    17.6828, 17.84793, 18.01306, 18.17819, 18.34332, 18.50845, 18.67357, 
    18.83868, 19.00379, 19.16888, 19.33397, 19.49904, 19.6641, 19.82914, 
    19.99416, 20.15916, 20.32415, 20.48911, 20.65404, 20.81895, 20.98383, 
    21.14868, 21.31351, 21.47829, 21.64305, 21.80777, 21.97245, 22.1371, 
    22.3017, 22.46626, 22.63078, 22.79526, 22.95968, 23.12406, 23.28839, 
    23.45267, 23.6169, 23.78107, 23.94518, 24.10924, 24.27324, 24.43718, 
    24.60105, 24.76487, 24.92861, 25.09229, 25.25591, 25.41945, 25.58292, 
    25.74632, 25.90965, 26.07289, 26.23607, 26.39916, 26.56217, 26.72511, 
    26.88795, 27.05072, 27.2134, 27.37599, 27.53849, 27.7009, 27.86322, 
    28.02545, 28.18758, 28.34962, 28.51156, 28.6734, 28.83514, 28.99678, 
    29.15832, 29.31975, 29.48108, 29.6423, 29.80341, 29.96441, 30.1253, 
    30.28608, 30.44675, 30.6073, 30.76773, 30.92805, 31.08825, 31.24833, 
    31.40828, 31.56812, 31.72783, 31.88741, 32.04688, 32.2062, 32.36541, 
    32.52448, 32.68342, 32.84223, 33.00091, 33.15945, 33.31786, 33.47612, 
    33.63425, 33.79224, 33.95009, 34.1078, 34.26537, 34.42279, 34.58006, 
    34.73719, 34.89418, 35.05101, 35.2077, 35.36423, 35.52062, 35.67685, 
    35.83293, 35.98885, 36.14462, 36.30023, 36.45568, 36.61098, 36.76612, 
    36.92109, 37.0759, 37.23056, 37.38504, 37.53937, 37.69353, 37.84752, 
    38.00135, 38.15501, 38.30849, 38.46181, 38.61496, 38.76794, 38.92075, 
    39.07338, 39.22584, 39.37812, 39.53023, 39.68216, 39.83392, 39.9855, 
    40.13689, 40.28811, 40.43915, 40.59001, 40.74069, 40.89118, 41.04149, 
    41.19162, 41.34156, 41.49132, 41.64089, 41.79028, 41.93948, 42.08849, 
    42.23731, 42.38594, 42.53439, 42.68264, 42.8307, 42.97857, 43.12625, 
    43.27374, 43.42103, 43.56813, 43.71503, 43.86174, 44.00826, 44.15458, 
    44.3007, 44.44662, 44.59235, 44.73788, 44.88321, 45.02834,
  -21.67017, -21.54432, -21.41825, -21.29198, -21.1655, -21.03881, -20.9119, 
    -20.78478, -20.65746, -20.52992, -20.40217, -20.27421, -20.14603, 
    -20.01765, -19.88905, -19.76024, -19.63122, -19.50199, -19.37254, 
    -19.24288, -19.11301, -18.98292, -18.85263, -18.72212, -18.59139, 
    -18.46046, -18.32931, -18.19795, -18.06637, -17.93458, -17.80258, 
    -17.67036, -17.53794, -17.40529, -17.27244, -17.13937, -17.00609, 
    -16.8726, -16.73889, -16.60497, -16.47083, -16.33648, -16.20193, 
    -16.06715, -15.93217, -15.79697, -15.66155, -15.52593, -15.39009, 
    -15.25404, -15.11778, -14.9813, -14.84461, -14.70772, -14.5706, 
    -14.43328, -14.29574, -14.158, -14.02004, -13.88187, -13.74349, -13.6049, 
    -13.46609, -13.32708, -13.18786, -13.04843, -12.90878, -12.76893, 
    -12.62887, -12.4886, -12.34811, -12.20743, -12.06653, -11.92542, 
    -11.78411, -11.64259, -11.50086, -11.35892, -11.21678, -11.07443, 
    -10.93188, -10.78912, -10.64615, -10.50298, -10.35961, -10.21603, 
    -10.07225, -9.928259, -9.78407, -9.639677, -9.495083, -9.350286, 
    -9.205289, -9.060091, -8.914692, -8.769093, -8.623295, -8.477297, 
    -8.3311, -8.184707, -8.038115, -7.891326, -7.74434, -7.597159, -7.449782, 
    -7.302211, -7.154445, -7.006485, -6.858332, -6.709986, -6.561448, 
    -6.412719, -6.263799, -6.114689, -5.96539, -5.815901, -5.666224, 
    -5.51636, -5.366309, -5.216072, -5.065649, -4.915041, -4.764249, 
    -4.613274, -4.462116, -4.310776, -4.159255, -4.007553, -3.855672, 
    -3.703612, -3.551373, -3.398958, -3.246366, -3.093598, -2.940656, 
    -2.787539, -2.634249, -2.480787, -2.327153, -2.173349, -2.019375, 
    -1.865232, -1.710921, -1.556444, -1.4018, -1.246991, -1.092017, 
    -0.9368805, -0.7815814, -0.6261209, -0.4705001, -0.3147198, -0.1587811, 
    -0.002684894, 0.1535677, 0.3099757, 0.4665381, 0.6232538, 0.7801218, 
    0.9371411, 1.094311, 1.251629, 1.409096, 1.566709, 1.724468, 1.882372, 
    2.04042, 2.19861, 2.356941, 2.515412, 2.674023, 2.832771, 2.991656, 
    3.150677, 3.309832, 3.46912, 3.628539, 3.78809, 3.94777, 4.107578, 
    4.267513, 4.427575, 4.58776, 4.748069, 4.908499, 5.069051, 5.229722, 
    5.39051, 5.551416, 5.712437, 5.873572, 6.034821, 6.19618, 6.35765, 
    6.519228, 6.680914, 6.842707, 7.004604, 7.166604, 7.328706, 7.490909, 
    7.653211, 7.815611, 7.978107, 8.140697, 8.303383, 8.466159, 8.629026, 
    8.791983, 8.955028, 9.118157, 9.281373, 9.444673, 9.608053, 9.771514, 
    9.935054, 10.09867, 10.26237, 10.42613, 10.58997, 10.75389, 10.91787, 
    11.08192, 11.24604, 11.41022, 11.57447, 11.73878, 11.90315, 12.06757, 
    12.23206, 12.3966, 12.5612, 12.72585, 12.89055, 13.0553, 13.2201, 
    13.38495, 13.54984, 13.71478, 13.87975, 14.04477, 14.20983, 14.37492, 
    14.54005, 14.70521, 14.8704, 15.03563, 15.20088, 15.36617, 15.53147, 
    15.6968, 15.86216, 16.02753, 16.19293, 16.35834, 16.52377, 16.68921, 
    16.85467, 17.02014, 17.18562, 17.3511, 17.51659, 17.68209, 17.84759, 
    18.01309, 18.17859, 18.34409, 18.50959, 18.67508, 18.84056, 19.00604, 
    19.1715, 19.33696, 19.5024, 19.66782, 19.83323, 19.99863, 20.164, 
    20.32935, 20.49468, 20.65998, 20.82526, 20.99051, 21.15573, 21.32092, 
    21.48608, 21.6512, 21.81629, 21.98134, 22.14635, 22.31132, 22.47624, 
    22.64113, 22.80597, 22.97076, 23.1355, 23.3002, 23.46484, 23.62943, 
    23.79396, 23.95844, 24.12286, 24.28722, 24.45152, 24.61576, 24.77993, 
    24.94403, 25.10807, 25.27205, 25.43595, 25.59978, 25.76353, 25.92722, 
    26.09082, 26.25435, 26.4178, 26.58117, 26.74445, 26.90765, 27.07077, 
    27.2338, 27.39674, 27.5596, 27.72236, 27.88503, 28.0476, 28.21008, 
    28.37247, 28.53476, 28.69694, 28.85903, 29.02101, 29.18289, 29.34467, 
    29.50634, 29.6679, 29.82935, 29.99069, 30.15192, 30.31304, 30.47404, 
    30.63493, 30.7957, 30.95635, 31.11689, 31.2773, 31.43759, 31.59775, 
    31.75779, 31.91771, 32.0775, 32.23716, 32.39669, 32.55609, 32.71535, 
    32.87449, 33.03349, 33.19235, 33.35107, 33.50967, 33.66811, 33.82642, 
    33.98459, 34.14262, 34.3005, 34.45823, 34.61582, 34.77327, 34.93056, 
    35.08771, 35.2447, 35.40155, 35.55824, 35.71478, 35.87116, 36.02739, 
    36.18346, 36.33937, 36.49513, 36.65072, 36.80616, 36.96143, 37.11654, 
    37.27149, 37.42627, 37.58089, 37.73534, 37.88963, 38.04374, 38.19769, 
    38.35147, 38.50507, 38.65851, 38.81177, 38.96486, 39.11777, 39.27052, 
    39.42308, 39.57547, 39.72768, 39.87971, 40.03156, 40.18324, 40.33473, 
    40.48604, 40.63717, 40.78811, 40.93888, 41.08945, 41.23985, 41.39006, 
    41.54008, 41.68991, 41.83956, 41.98902, 42.13829, 42.28737, 42.43626, 
    42.58496, 42.73346, 42.88178, 43.0299, 43.17783, 43.32557, 43.47311, 
    43.62045, 43.7676, 43.91456, 44.06132, 44.20788, 44.35424, 44.5004, 
    44.64637, 44.79214, 44.93771, 45.08307,
  -21.74192, -21.61594, -21.48974, -21.36334, -21.23672, -21.10989, 
    -20.98285, -20.8556, -20.72813, -20.60045, -20.47256, -20.34446, 
    -20.21614, -20.08761, -19.95887, -19.82992, -19.70075, -19.57137, 
    -19.44177, -19.31196, -19.18194, -19.0517, -18.92125, -18.79059, 
    -18.65971, -18.52862, -18.39731, -18.26579, -18.13406, -18.00211, 
    -17.86994, -17.73757, -17.60497, -17.47217, -17.33915, -17.20591, 
    -17.07246, -16.9388, -16.80492, -16.67083, -16.53652, -16.402, -16.26727, 
    -16.13232, -15.99715, -15.86178, -15.72618, -15.59038, -15.45436, 
    -15.31813, -15.18168, -15.04502, -14.90815, -14.77106, -14.63376, 
    -14.49625, -14.35852, -14.22058, -14.08243, -13.94407, -13.80549, 
    -13.6667, -13.5277, -13.38849, -13.24907, -13.10943, -12.96959, 
    -12.82953, -12.68926, -12.54879, -12.4081, -12.2672, -12.12609, 
    -11.98478, -11.84325, -11.70152, -11.55958, -11.41743, -11.27507, 
    -11.1325, -10.98973, -10.84675, -10.70356, -10.56017, -10.41657, 
    -10.27276, -10.12875, -9.984541, -9.840122, -9.6955, -9.550675, 
    -9.405647, -9.260416, -9.114983, -8.969348, -8.823512, -8.677475, 
    -8.531239, -8.384801, -8.238165, -8.091331, -7.944297, -7.797066, 
    -7.649638, -7.502014, -7.354193, -7.206176, -7.057965, -6.909559, 
    -6.76096, -6.612166, -6.463181, -6.314004, -6.164635, -6.015076, 
    -5.865326, -5.715387, -5.565259, -5.414943, -5.26444, -5.11375, 
    -4.962874, -4.811812, -4.660567, -4.509137, -4.357524, -4.205729, 
    -4.053752, -3.901594, -3.749257, -3.59674, -3.444044, -3.291171, 
    -3.138121, -2.984895, -2.831494, -2.677918, -2.524169, -2.370248, 
    -2.216154, -2.06189, -1.907456, -1.752853, -1.598081, -1.443143, 
    -1.288038, -1.132767, -0.9773327, -0.8217345, -0.6659738, -0.5100517, 
    -0.3539691, -0.1977269, -0.04132627, 0.1152319, 0.2719465, 0.4288166, 
    0.585841, 0.7430188, 0.9003488, 1.05783, 1.215461, 1.373242, 1.53117, 
    1.689245, 1.847466, 2.005831, 2.16434, 2.322992, 2.481784, 2.640716, 
    2.799787, 2.958996, 3.118341, 3.277822, 3.437436, 3.597184, 3.757063, 
    3.917072, 4.07721, 4.237477, 4.39787, 4.558388, 4.719031, 4.879796, 
    5.040683, 5.20169, 5.362816, 5.52406, 5.68542, 5.846895, 6.008483, 
    6.170184, 6.331996, 6.493917, 6.655947, 6.818084, 6.980326, 7.142672, 
    7.305121, 7.467671, 7.630321, 7.79307, 7.955915, 8.118856, 8.281892, 
    8.445021, 8.60824, 8.771549, 8.934947, 9.098432, 9.262002, 9.425656, 
    9.589393, 9.75321, 9.917108, 10.08108, 10.24513, 10.40926, 10.57346, 
    10.73773, 10.90208, 11.06649, 11.23097, 11.39551, 11.56012, 11.72479, 
    11.88953, 12.05432, 12.21917, 12.38408, 12.54904, 12.71405, 12.87912, 
    13.04424, 13.2094, 13.37462, 13.53988, 13.70518, 13.87052, 14.03591, 
    14.20133, 14.36679, 14.53229, 14.69782, 14.86339, 15.02898, 15.1946, 
    15.36026, 15.52593, 15.69164, 15.85736, 16.02311, 16.18887, 16.35466, 
    16.52046, 16.68627, 16.8521, 17.01794, 17.18379, 17.34964, 17.51551, 
    17.68138, 17.84725, 18.01312, 18.17899, 18.34486, 18.51073, 18.67659, 
    18.84245, 19.0083, 19.17413, 19.33996, 19.50577, 19.67157, 19.83735, 
    20.00311, 20.16886, 20.33458, 20.50027, 20.66595, 20.8316, 20.99722, 
    21.16281, 21.32837, 21.49389, 21.65938, 21.82484, 21.99026, 22.15564, 
    22.32097, 22.48627, 22.65152, 22.81672, 22.98188, 23.14699, 23.31205, 
    23.47706, 23.64201, 23.80691, 23.97175, 24.13654, 24.30126, 24.46592, 
    24.63052, 24.79506, 24.95952, 25.12392, 25.28826, 25.45252, 25.6167, 
    25.78082, 25.94486, 26.10882, 26.27271, 26.43651, 26.60024, 26.76388, 
    26.92743, 27.09091, 27.25429, 27.41759, 27.58079, 27.7439, 27.90693, 
    28.06985, 28.23268, 28.39541, 28.55805, 28.72058, 28.88301, 29.04535, 
    29.20757, 29.36969, 29.5317, 29.69361, 29.8554, 30.01708, 30.17866, 
    30.34011, 30.50145, 30.66268, 30.82379, 30.98478, 31.14564, 31.30639, 
    31.46701, 31.62751, 31.78788, 31.94813, 32.10825, 32.26824, 32.42809, 
    32.58782, 32.74741, 32.90687, 33.0662, 33.22538, 33.38443, 33.54334, 
    33.70211, 33.86074, 34.01923, 34.17757, 34.33577, 34.49382, 34.65173, 
    34.80948, 34.96709, 35.12455, 35.28185, 35.43901, 35.59601, 35.75285, 
    35.90954, 36.06608, 36.22245, 36.37867, 36.53473, 36.69062, 36.84636, 
    37.00193, 37.15734, 37.31258, 37.46766, 37.62257, 37.77732, 37.9319, 
    38.0863, 38.24054, 38.39461, 38.5485, 38.70222, 38.85577, 39.00914, 
    39.16234, 39.31536, 39.46821, 39.62088, 39.77337, 39.92567, 40.0778, 
    40.22975, 40.38152, 40.5331, 40.68451, 40.83572, 40.98675, 41.1376, 
    41.28826, 41.43873, 41.58902, 41.73912, 41.88903, 42.03875, 42.18827, 
    42.33761, 42.48676, 42.63572, 42.78448, 42.93305, 43.08142, 43.2296, 
    43.37759, 43.52538, 43.67297, 43.82037, 43.96757, 44.11457, 44.26138, 
    44.40798, 44.55438, 44.70059, 44.8466, 44.9924, 45.138,
  -21.81388, -21.68777, -21.56144, -21.4349, -21.30815, -21.18118, -21.05401, 
    -20.92662, -20.79901, -20.67119, -20.54316, -20.41492, -20.28646, 
    -20.15779, -20.0289, -19.8998, -19.77048, -19.64095, -19.51121, 
    -19.38125, -19.25108, -19.12069, -18.99009, -18.85927, -18.72824, 
    -18.59699, -18.46552, -18.33385, -18.20195, -18.06984, -17.93752, 
    -17.80498, -17.67222, -17.53925, -17.40606, -17.27266, -17.13904, 
    -17.00521, -16.87116, -16.7369, -16.60242, -16.46773, -16.33282, 
    -16.19769, -16.06235, -15.92679, -15.79102, -15.65504, -15.51884, 
    -15.38242, -15.24579, -15.10894, -14.97189, -14.83461, -14.69712, 
    -14.55942, -14.4215, -14.28337, -14.14503, -14.00647, -13.8677, 
    -13.72871, -13.58952, -13.45011, -13.31048, -13.17065, -13.0306, 
    -12.89034, -12.74987, -12.60918, -12.46829, -12.32718, -12.18587, 
    -12.04434, -11.9026, -11.76065, -11.6185, -11.47613, -11.33356, 
    -11.19077, -11.04778, -10.90458, -10.76117, -10.61755, -10.47373, 
    -10.3297, -10.18546, -10.04102, -9.896376, -9.751523, -9.606466, 
    -9.461205, -9.315741, -9.170073, -9.024201, -8.878128, -8.731853, 
    -8.585376, -8.438698, -8.291819, -8.14474, -7.997463, -7.849986, 
    -7.70231, -7.554437, -7.406367, -7.258099, -7.109636, -6.960977, 
    -6.812123, -6.663074, -6.513832, -6.364396, -6.214768, -6.064948, 
    -5.914937, -5.764735, -5.614343, -5.463761, -5.312992, -5.162034, 
    -5.010889, -4.859558, -4.70804, -4.556338, -4.404451, -4.252381, 
    -4.100128, -3.947694, -3.795077, -3.642281, -3.489305, -3.33615, 
    -3.182817, -3.029306, -2.87562, -2.721758, -2.567721, -2.413511, 
    -2.259127, -2.104572, -1.949846, -1.794949, -1.639883, -1.484649, 
    -1.329247, -1.173679, -1.017946, -0.8620473, -0.7059855, -0.5497611, 
    -0.3933752, -0.2368286, -0.08012246, 0.07674225, 0.2337645, 0.3909433, 
    0.5482774, 0.705766, 0.8634079, 1.021202, 1.179147, 1.337243, 1.495487, 
    1.653879, 1.812418, 1.971102, 2.129931, 2.288903, 2.448018, 2.607273, 
    2.766668, 2.926202, 3.085873, 3.24568, 3.405622, 3.565699, 3.725907, 
    3.886247, 4.046717, 4.207316, 4.368042, 4.528894, 4.689872, 4.850973, 
    5.012197, 5.173542, 5.335006, 5.496589, 5.658289, 5.820106, 5.982036, 
    6.144079, 6.306235, 6.4685, 6.630875, 6.793357, 6.955946, 7.118639, 
    7.281436, 7.444335, 7.607335, 7.770433, 7.93363, 8.096923, 8.26031, 
    8.423792, 8.587365, 8.751028, 8.914782, 9.078622, 9.242548, 9.406559, 
    9.570653, 9.734829, 9.899084, 10.06342, 10.22783, 10.39232, 10.55688, 
    10.72151, 10.88622, 11.05099, 11.21583, 11.38074, 11.54571, 11.71075, 
    11.87585, 12.04101, 12.20622, 12.3715, 12.53682, 12.70221, 12.86764, 
    13.03312, 13.19866, 13.36424, 13.52987, 13.69554, 13.86125, 14.02701, 
    14.1928, 14.35863, 14.5245, 14.6904, 14.85634, 15.0223, 15.1883, 
    15.35432, 15.52037, 15.68645, 15.85254, 16.01866, 16.1848, 16.35096, 
    16.51713, 16.68332, 16.84952, 17.01573, 17.18195, 17.34818, 17.51442, 
    17.68066, 17.8469, 18.01315, 18.17939, 18.34564, 18.51188, 18.67811, 
    18.84434, 19.01056, 19.17677, 19.34297, 19.50916, 19.67533, 19.84148, 
    20.00762, 20.17373, 20.33983, 20.5059, 20.67194, 20.83796, 21.00395, 
    21.16991, 21.33584, 21.50174, 21.6676, 21.83343, 21.99922, 22.16496, 
    22.33067, 22.49634, 22.66195, 22.82753, 22.99306, 23.15853, 23.32396, 
    23.48933, 23.65465, 23.81992, 23.98512, 24.15027, 24.31536, 24.48039, 
    24.64535, 24.81025, 24.97508, 25.13984, 25.30453, 25.46916, 25.63371, 
    25.79818, 25.96258, 26.1269, 26.29115, 26.45531, 26.61939, 26.78339, 
    26.9473, 27.11113, 27.27487, 27.43852, 27.60207, 27.76554, 27.92891, 
    28.09219, 28.25537, 28.41846, 28.58144, 28.74432, 28.9071, 29.06978, 
    29.23235, 29.39482, 29.55717, 29.71942, 29.88156, 30.04359, 30.2055, 
    30.3673, 30.52898, 30.69054, 30.85199, 31.01331, 31.17452, 31.3356, 
    31.49656, 31.65739, 31.8181, 31.97868, 32.13913, 32.29944, 32.45963, 
    32.61969, 32.77961, 32.93939, 33.09904, 33.25856, 33.41793, 33.57716, 
    33.73625, 33.8952, 34.05401, 34.21267, 34.37119, 34.52956, 34.68777, 
    34.84585, 35.00377, 35.16154, 35.31916, 35.47662, 35.63393, 35.79108, 
    35.94808, 36.10492, 36.2616, 36.41813, 36.57449, 36.73068, 36.88672, 
    37.04259, 37.1983, 37.35384, 37.50922, 37.66442, 37.81946, 37.97433, 
    38.12903, 38.28356, 38.43792, 38.5921, 38.74611, 38.89994, 39.0536, 
    39.20708, 39.36039, 39.51352, 39.66646, 39.81923, 39.97182, 40.12423, 
    40.27645, 40.42849, 40.58035, 40.73202, 40.88351, 41.03481, 41.18592, 
    41.33685, 41.48759, 41.63815, 41.78851, 41.93868, 42.08866, 42.23845, 
    42.38805, 42.53745, 42.68666, 42.83568, 42.9845, 43.13313, 43.28157, 
    43.4298, 43.57784, 43.72569, 43.87333, 44.02077, 44.16802, 44.31507, 
    44.46191, 44.60856, 44.755, 44.90125, 45.04729, 45.19313,
  -21.88605, -21.75981, -21.63335, -21.50667, -21.37979, -21.25269, 
    -21.12537, -20.99784, -20.8701, -20.74215, -20.61397, -20.48559, 
    -20.35699, -20.22817, -20.09914, -19.96989, -19.84043, -19.71075, 
    -19.58086, -19.45075, -19.32043, -19.18989, -19.05913, -18.92816, 
    -18.79697, -18.66557, -18.53395, -18.40211, -18.27006, -18.13779, 
    -18.0053, -17.8726, -17.73968, -17.60654, -17.47319, -17.33962, 
    -17.20584, -17.07183, -16.93762, -16.80318, -16.66853, -16.53366, 
    -16.39858, -16.26328, -16.12776, -15.99202, -15.85607, -15.71991, 
    -15.58352, -15.44693, -15.31011, -15.17308, -15.03584, -14.89837, 
    -14.7607, -14.6228, -14.4847, -14.34637, -14.20784, -14.06908, -13.93012, 
    -13.79094, -13.65154, -13.51193, -13.37211, -13.23207, -13.09182, 
    -12.95135, -12.81068, -12.66979, -12.52869, -12.38737, -12.24584, 
    -12.10411, -11.96216, -11.81999, -11.67762, -11.53504, -11.39225, 
    -11.24924, -11.10603, -10.96261, -10.81898, -10.67514, -10.53109, 
    -10.38684, -10.24238, -10.09771, -9.952829, -9.807747, -9.662458, 
    -9.516964, -9.371265, -9.225362, -9.079253, -8.932942, -8.786427, 
    -8.63971, -8.49279, -8.345669, -8.198346, -8.050823, -7.9031, -7.755177, 
    -7.607055, -7.458734, -7.310215, -7.161499, -7.012586, -6.863477, 
    -6.714172, -6.564672, -6.414978, -6.26509, -6.115008, -5.964735, 
    -5.814269, -5.663612, -5.512765, -5.361728, -5.210502, -5.059087, 
    -4.907485, -4.755696, -4.60372, -4.451559, -4.299213, -4.146684, 
    -3.993971, -3.841076, -3.687999, -3.534741, -3.381303, -3.227686, 
    -3.073891, -2.919919, -2.765769, -2.611444, -2.456944, -2.30227, 
    -2.147422, -1.992403, -1.837212, -1.681851, -1.52632, -1.370621, 
    -1.214754, -1.05872, -0.902521, -0.7461571, -0.5896295, -0.4329393, 
    -0.2760873, -0.1190747, 0.03809764, 0.1954286, 0.352917, 0.510562, 
    0.6683624, 0.8263173, 0.9844254, 1.142686, 1.301097, 1.459658, 1.618369, 
    1.777227, 1.936231, 2.095381, 2.254676, 2.414113, 2.573693, 2.733413, 
    2.893272, 3.053271, 3.213406, 3.373677, 3.534083, 3.694622, 3.855294, 
    4.016097, 4.177029, 4.33809, 4.499278, 4.660592, 4.82203, 4.983592, 
    5.145276, 5.30708, 5.469004, 5.631045, 5.793203, 5.955477, 6.117865, 
    6.280365, 6.442976, 6.605697, 6.768526, 6.931463, 7.094505, 7.257651, 
    7.4209, 7.58425, 7.747701, 7.91125, 8.074896, 8.238637, 8.402472, 
    8.566401, 8.73042, 8.894529, 9.058726, 9.22301, 9.38738, 9.551833, 
    9.716368, 9.880983, 10.04568, 10.21045, 10.3753, 10.54022, 10.70522, 
    10.87029, 11.03543, 11.20063, 11.36591, 11.53124, 11.69665, 11.86211, 
    12.02763, 12.19322, 12.35886, 12.52456, 12.69031, 12.85611, 13.02196, 
    13.18787, 13.35382, 13.51982, 13.68586, 13.85194, 14.01807, 14.18423, 
    14.35044, 14.51668, 14.68295, 14.84926, 15.0156, 15.18196, 15.34836, 
    15.51478, 15.68123, 15.8477, 16.0142, 16.18071, 16.34724, 16.51379, 
    16.68035, 16.84692, 17.01351, 17.18011, 17.34671, 17.51332, 17.67994, 
    17.84656, 18.01318, 18.1798, 18.34642, 18.51303, 18.67964, 18.84625, 
    19.01284, 19.17943, 19.346, 19.51256, 19.6791, 19.84563, 20.01214, 
    20.17863, 20.3451, 20.51154, 20.67796, 20.84435, 21.01072, 21.17705, 
    21.34335, 21.50962, 21.67586, 21.84205, 22.00821, 22.17433, 22.34041, 
    22.50644, 22.67244, 22.83838, 23.00428, 23.17012, 23.33592, 23.50166, 
    23.66735, 23.83298, 23.99855, 24.16407, 24.32952, 24.49492, 24.66024, 
    24.8255, 24.9907, 25.15583, 25.32088, 25.48587, 25.65078, 25.81562, 
    25.98038, 26.14506, 26.30966, 26.47419, 26.63863, 26.80298, 26.96725, 
    27.13144, 27.29553, 27.45954, 27.62345, 27.78727, 27.951, 28.11463, 
    28.27816, 28.4416, 28.60493, 28.76816, 28.93129, 29.09432, 29.25724, 
    29.42005, 29.58275, 29.74535, 29.90783, 30.0702, 30.23245, 30.39459, 
    30.55662, 30.71852, 30.88031, 31.04197, 31.20352, 31.36493, 31.52623, 
    31.6874, 31.84844, 32.00935, 32.17013, 32.33078, 32.4913, 32.65168, 
    32.81194, 32.97205, 33.13202, 33.29186, 33.45156, 33.61112, 33.77053, 
    33.9298, 34.08893, 34.24791, 34.40675, 34.56543, 34.72397, 34.88236, 
    35.0406, 35.19868, 35.35661, 35.51439, 35.672, 35.82947, 35.98677, 
    36.14392, 36.30091, 36.45774, 36.6144, 36.7709, 36.92724, 37.08341, 
    37.23942, 37.39526, 37.55093, 37.70644, 37.86177, 38.01694, 38.17193, 
    38.32675, 38.4814, 38.63587, 38.79016, 38.94429, 39.09823, 39.252, 
    39.40559, 39.55899, 39.71223, 39.86527, 40.01814, 40.17082, 40.32333, 
    40.47564, 40.62777, 40.77972, 40.93148, 41.08305, 41.23444, 41.38563, 
    41.53664, 41.68746, 41.83808, 41.98852, 42.13876, 42.28881, 42.43867, 
    42.58833, 42.7378, 42.88708, 43.03616, 43.18504, 43.33372, 43.48221, 
    43.6305, 43.77859, 43.92648, 44.07417, 44.22166, 44.36895, 44.51604, 
    44.66293, 44.80962, 44.9561, 45.10238, 45.24846,
  -21.95843, -21.83205, -21.70546, -21.57866, -21.45163, -21.3244, -21.19695, 
    -21.06928, -20.9414, -20.8133, -20.68499, -20.55647, -20.42772, 
    -20.29876, -20.16959, -20.0402, -19.91059, -19.78077, -19.65072, 
    -19.52047, -19.38999, -19.2593, -19.12839, -18.99726, -18.86592, 
    -18.73436, -18.60258, -18.47059, -18.33838, -18.20595, -18.0733, 
    -17.94043, -17.80735, -17.67405, -17.54053, -17.4068, -17.27284, 
    -17.13867, -17.00428, -16.86967, -16.73485, -16.59981, -16.46455, 
    -16.32907, -16.19338, -16.05746, -15.92134, -15.78499, -15.64843, 
    -15.51164, -15.37465, -15.23743, -15.1, -14.96235, -14.82448, -14.6864, 
    -14.5481, -14.40959, -14.27086, -14.13191, -13.99275, -13.85337, 
    -13.71377, -13.57397, -13.43394, -13.2937, -13.15325, -13.01258, 
    -12.8717, -12.7306, -12.58929, -12.44777, -12.30603, -12.16408, 
    -12.02192, -11.87954, -11.73696, -11.59416, -11.45115, -11.30793, 
    -11.16449, -11.02085, -10.877, -10.73293, -10.58866, -10.44418, 
    -10.29949, -10.15459, -10.00949, -9.864173, -9.718652, -9.572925, 
    -9.426991, -9.28085, -9.134506, -8.987956, -8.841202, -8.694243, 
    -8.547082, -8.399717, -8.25215, -8.104381, -7.95641, -7.808239, 
    -7.659867, -7.511296, -7.362525, -7.213556, -7.064388, -6.915023, 
    -6.765461, -6.615704, -6.46575, -6.315601, -6.165258, -6.014721, 
    -5.863992, -5.713069, -5.561955, -5.41065, -5.259155, -5.10747, 
    -4.955596, -4.803535, -4.651285, -4.498849, -4.346227, -4.193419, 
    -4.040428, -3.887253, -3.733895, -3.580354, -3.426633, -3.272732, 
    -3.118651, -2.964391, -2.809953, -2.655339, -2.500548, -2.345582, 
    -2.190442, -2.035129, -1.879643, -1.723985, -1.568157, -1.412159, 
    -1.255992, -1.099658, -0.9431568, -0.7864898, -0.6296581, -0.4726625, 
    -0.3155042, -0.158184, -0.000703152, 0.1569374, 0.3147367, 0.4726935, 
    0.6308068, 0.7890756, 0.9474987, 1.106075, 1.264804, 1.423683, 1.582713, 
    1.741891, 1.901217, 2.060689, 2.220307, 2.380068, 2.539973, 2.70002, 
    2.860207, 3.020533, 3.180997, 3.341599, 3.502336, 3.663207, 3.824212, 
    3.985348, 4.146616, 4.308012, 4.469537, 4.631188, 4.792965, 4.954866, 
    5.11689, 5.279036, 5.441301, 5.603686, 5.766188, 5.928806, 6.091538, 
    6.254385, 6.417343, 6.580411, 6.743589, 6.906875, 7.070267, 7.233765, 
    7.397365, 7.561068, 7.724871, 7.888773, 8.052773, 8.21687, 8.381062, 
    8.545346, 8.709723, 8.87419, 9.038746, 9.203389, 9.368118, 9.532931, 
    9.697827, 9.862805, 10.02786, 10.193, 10.35821, 10.5235, 10.68886, 
    10.85429, 11.01979, 11.18537, 11.35101, 11.51671, 11.68248, 11.84831, 
    12.0142, 12.18016, 12.34617, 12.51223, 12.67835, 12.84453, 13.01075, 
    13.17703, 13.34335, 13.50972, 13.67613, 13.84259, 14.00909, 14.17563, 
    14.3422, 14.50882, 14.67547, 14.84215, 15.00886, 15.1756, 15.34238, 
    15.50917, 15.676, 15.84284, 16.00971, 16.1766, 16.34351, 16.51043, 
    16.67737, 16.84432, 17.01128, 17.17825, 17.34523, 17.51222, 17.67921, 
    17.84621, 18.01321, 18.18021, 18.3472, 18.51419, 18.68118, 18.84816, 
    19.01513, 19.18209, 19.34904, 19.51598, 19.6829, 19.8498, 20.01669, 
    20.18355, 20.35039, 20.51721, 20.68401, 20.85077, 21.01751, 21.18422, 
    21.3509, 21.51754, 21.68415, 21.85072, 22.01725, 22.18374, 22.35019, 
    22.5166, 22.68296, 22.84928, 23.01554, 23.18176, 23.34793, 23.51404, 
    23.6801, 23.8461, 24.01204, 24.17792, 24.34375, 24.5095, 24.6752, 
    24.84083, 25.00639, 25.17188, 25.33731, 25.50265, 25.66793, 25.83313, 
    25.99825, 26.1633, 26.32826, 26.49314, 26.65795, 26.82266, 26.98729, 
    27.15183, 27.31628, 27.48065, 27.64492, 27.80909, 27.97318, 28.13716, 
    28.30105, 28.46483, 28.62852, 28.7921, 28.95559, 29.11896, 29.28223, 
    29.44539, 29.60844, 29.77138, 29.93421, 30.09693, 30.25953, 30.42201, 
    30.58437, 30.74662, 30.90875, 31.07075, 31.23263, 31.39439, 31.55602, 
    31.71753, 31.8789, 32.04015, 32.20126, 32.36225, 32.5231, 32.68382, 
    32.84439, 33.00484, 33.16514, 33.32531, 33.48533, 33.64521, 33.80495, 
    33.96455, 34.124, 34.2833, 34.44245, 34.60146, 34.76031, 34.91902, 
    35.07757, 35.23597, 35.39421, 35.5523, 35.71024, 35.86801, 36.02562, 
    36.18308, 36.34037, 36.49751, 36.65448, 36.81128, 36.96792, 37.1244, 
    37.28071, 37.43685, 37.59282, 37.74862, 37.90425, 38.05971, 38.21499, 
    38.37011, 38.52504, 38.67981, 38.8344, 38.9888, 39.14304, 39.29709, 
    39.45096, 39.60465, 39.75817, 39.9115, 40.06464, 40.2176, 40.37038, 
    40.52298, 40.67538, 40.8276, 40.97963, 41.13148, 41.28313, 41.4346, 
    41.58587, 41.73695, 41.88785, 42.03855, 42.18905, 42.33937, 42.48948, 
    42.6394, 42.78913, 42.93866, 43.088, 43.23713, 43.38607, 43.53481, 
    43.68335, 43.83169, 43.97983, 44.12777, 44.27551, 44.42304, 44.57037, 
    44.7175, 44.86443, 45.01115, 45.15767, 45.30398,
  -22.03102, -21.90451, -21.77778, -21.65084, -21.52369, -21.39632, 
    -21.26873, -21.14093, -21.01291, -20.88468, -20.75623, -20.62756, 
    -20.49867, -20.36957, -20.24025, -20.11071, -19.98096, -19.85099, 
    -19.7208, -19.59039, -19.45976, -19.32892, -19.19786, -19.06658, 
    -18.93508, -18.80337, -18.67143, -18.53928, -18.40691, -18.27432, 
    -18.14151, -18.00848, -17.87523, -17.74177, -17.60809, -17.47418, 
    -17.34006, -17.20572, -17.07116, -16.93638, -16.80139, -16.66617, 
    -16.53074, -16.39508, -16.25921, -16.12312, -15.98681, -15.85028, 
    -15.71354, -15.57657, -15.43939, -15.30199, -15.16437, -15.02654, 
    -14.88848, -14.75021, -14.61172, -14.47301, -14.33409, -14.19495, 
    -14.05559, -13.91601, -13.77622, -13.63621, -13.49599, -13.35554, 
    -13.21489, -13.07401, -12.93293, -12.79162, -12.65011, -12.50837, 
    -12.36643, -12.22426, -12.08189, -11.9393, -11.7965, -11.65348, 
    -11.51025, -11.36681, -11.22316, -11.0793, -10.93522, -10.79093, 
    -10.64644, -10.50173, -10.35681, -10.21168, -10.06635, -9.920802, 
    -9.775049, -9.629087, -9.482919, -9.336542, -9.18996, -9.043171, 
    -8.896176, -8.748977, -8.601573, -8.453964, -8.306152, -8.158136, 
    -8.009918, -7.861498, -7.712876, -7.564054, -7.41503, -7.265807, 
    -7.116385, -6.966763, -6.816945, -6.666928, -6.516714, -6.366304, 
    -6.215699, -6.064898, -5.913903, -5.762715, -5.611334, -5.45976, 
    -5.307995, -5.156039, -5.003893, -4.851558, -4.699033, -4.546321, 
    -4.393422, -4.240337, -4.087066, -3.93361, -3.77997, -3.626147, 
    -3.472141, -3.317954, -3.163586, -3.009038, -2.854312, -2.699407, 
    -2.544325, -2.389067, -2.233633, -2.078024, -1.922242, -1.766287, 
    -1.610161, -1.453864, -1.297396, -1.14076, -0.983956, -0.826985, 
    -0.6698481, -0.5125462, -0.3550805, -0.1974518, -0.03966132, 0.11829, 
    0.276401, 0.4346707, 0.593098, 0.7516818, 0.9104211, 1.069315, 1.228361, 
    1.38756, 1.54691, 1.70641, 1.866058, 2.025854, 2.185796, 2.345883, 
    2.506114, 2.666488, 2.827003, 2.987659, 3.148454, 3.309387, 3.470456, 
    3.631661, 3.793, 3.954472, 4.116075, 4.277809, 4.439671, 4.601662, 
    4.763778, 4.92602, 5.088386, 5.250873, 5.413482, 5.57621, 5.739058, 
    5.902021, 6.065101, 6.228294, 6.391601, 6.555019, 6.718546, 6.882183, 
    7.045927, 7.209776, 7.373729, 7.537786, 7.701943, 7.866201, 8.030558, 
    8.19501, 8.359559, 8.524202, 8.688937, 8.853764, 9.01868, 9.183683, 
    9.348773, 9.513948, 9.679207, 9.844547, 10.00997, 10.17547, 10.34105, 
    10.5067, 10.67242, 10.83822, 11.00409, 11.17003, 11.33604, 11.50212, 
    11.66825, 11.83445, 12.00072, 12.16704, 12.33342, 12.49986, 12.66635, 
    12.8329, 12.99949, 13.16614, 13.33284, 13.49958, 13.66637, 13.8332, 
    14.00007, 14.16698, 14.33394, 14.50093, 14.66795, 14.83501, 15.0021, 
    15.16922, 15.33636, 15.50354, 15.67074, 15.83796, 16.00521, 16.17247, 
    16.33976, 16.50706, 16.67437, 16.8417, 17.00904, 17.17639, 17.34375, 
    17.51112, 17.67849, 17.84586, 18.01324, 18.18061, 18.34799, 18.51536, 
    18.68272, 18.85008, 19.01743, 19.18477, 19.35209, 19.51941, 19.68671, 
    19.85399, 20.02125, 20.18849, 20.35571, 20.52291, 20.69008, 20.85722, 
    21.02434, 21.19142, 21.35847, 21.52549, 21.69247, 21.85942, 22.02633, 
    22.19319, 22.36002, 22.5268, 22.69353, 22.86022, 23.02686, 23.19345, 
    23.35999, 23.52647, 23.6929, 23.85927, 24.02559, 24.19184, 24.35803, 
    24.52416, 24.69022, 24.85622, 25.02215, 25.18801, 25.3538, 25.51951, 
    25.68515, 25.85072, 26.0162, 26.18161, 26.34694, 26.51219, 26.67735, 
    26.84242, 27.00741, 27.17232, 27.33713, 27.50185, 27.66648, 27.83101, 
    27.99545, 28.15979, 28.32403, 28.48817, 28.65221, 28.81615, 28.97998, 
    29.14371, 29.30733, 29.47084, 29.63424, 29.79753, 29.9607, 30.12376, 
    30.28671, 30.44954, 30.61225, 30.77484, 30.93731, 31.09965, 31.26188, 
    31.42397, 31.58594, 31.74778, 31.9095, 32.07108, 32.23253, 32.39385, 
    32.55503, 32.71608, 32.87699, 33.03776, 33.1984, 33.35889, 33.51924, 
    33.67945, 33.83952, 33.99943, 34.15921, 34.31883, 34.47831, 34.63763, 
    34.79681, 34.95583, 35.1147, 35.27341, 35.43197, 35.59037, 35.74862, 
    35.90671, 36.06463, 36.2224, 36.38, 36.53744, 36.69472, 36.85183, 
    37.00877, 37.16555, 37.32216, 37.4786, 37.63487, 37.79097, 37.9469, 
    38.10265, 38.25823, 38.41364, 38.56887, 38.72392, 38.8788, 39.0335, 
    39.18801, 39.34236, 39.49651, 39.65049, 39.80429, 39.9579, 40.11132, 
    40.26456, 40.41762, 40.57049, 40.72317, 40.87567, 41.02797, 41.18009, 
    41.33202, 41.48375, 41.63529, 41.78664, 41.9378, 42.08876, 42.23954, 
    42.39011, 42.54049, 42.69067, 42.84066, 42.99044, 43.14003, 43.28942, 
    43.43862, 43.58761, 43.7364, 43.88499, 44.03338, 44.18156, 44.32955, 
    44.47733, 44.6249, 44.77227, 44.91944, 45.06641, 45.21316, 45.35971,
  -22.10381, -21.97717, -21.85032, -21.72325, -21.59596, -21.46845, 
    -21.34073, -21.21279, -21.08463, -20.95626, -20.82767, -20.69886, 
    -20.56983, -20.44059, -20.31112, -20.18144, -20.05154, -19.92142, 
    -19.79109, -19.66053, -19.52975, -19.39876, -19.26755, -19.13611, 
    -19.00446, -18.87259, -18.7405, -18.60818, -18.47565, -18.3429, 
    -18.20993, -18.07674, -17.94333, -17.8097, -17.67585, -17.54178, 
    -17.40749, -17.27299, -17.13826, -17.00331, -16.86814, -16.73275, 
    -16.59714, -16.46131, -16.32526, -16.18899, -16.0525, -15.91579, 
    -15.77887, -15.64172, -15.50435, -15.36677, -15.22896, -15.09094, 
    -14.95269, -14.81423, -14.67555, -14.53665, -14.39753, -14.25819, 
    -14.11864, -13.97887, -13.83888, -13.69867, -13.55824, -13.4176, 
    -13.27674, -13.13566, -12.99437, -12.85286, -12.71113, -12.56919, 
    -12.42703, -12.28466, -12.14207, -11.99927, -11.85625, -11.71302, 
    -11.56957, -11.42591, -11.28204, -11.13795, -10.99365, -10.84914, 
    -10.70442, -10.55948, -10.41434, -10.26898, -10.12341, -9.977637, 
    -9.831651, -9.685454, -9.53905, -9.392437, -9.245617, -9.098589, 
    -8.951354, -8.803912, -8.656264, -8.508411, -8.360354, -8.212091, 
    -8.063625, -7.914956, -7.766084, -7.617009, -7.467733, -7.318255, 
    -7.168577, -7.018699, -6.868622, -6.718346, -6.567872, -6.4172, 
    -6.266331, -6.115266, -5.964006, -5.812551, -5.660902, -5.509059, 
    -5.357023, -5.204795, -5.052376, -4.899767, -4.746967, -4.593978, 
    -4.440802, -4.287437, -4.133885, -3.980148, -3.826225, -3.672118, 
    -3.517828, -3.363354, -3.208699, -3.053863, -2.898846, -2.74365, 
    -2.588276, -2.432724, -2.276995, -2.121091, -1.965012, -1.808759, 
    -1.652333, -1.495736, -1.338967, -1.182028, -1.02492, -0.8676438, 
    -0.7102007, -0.5525916, -0.3948174, -0.2368792, -0.07877808, 0.07948495, 
    0.2379088, 0.3964925, 0.5552348, 0.7141348, 0.8731912, 1.032403, 
    1.191769, 1.351288, 1.51096, 1.670782, 1.830753, 1.990874, 2.151141, 
    2.311555, 2.472114, 2.632817, 2.793662, 2.954648, 3.115775, 3.27704, 
    3.438443, 3.599982, 3.761657, 3.923465, 4.085406, 4.247478, 4.409679, 
    4.57201, 4.734468, 4.897051, 5.05976, 5.222591, 5.385545, 5.548619, 
    5.711812, 5.875123, 6.03855, 6.202093, 6.365749, 6.529517, 6.693397, 
    6.857385, 7.021482, 7.185684, 7.349992, 7.514404, 7.678917, 7.843532, 
    8.008245, 8.173057, 8.337964, 8.502966, 8.668061, 8.833248, 8.998526, 
    9.163892, 9.329345, 9.494884, 9.660506, 9.826211, 9.991997, 10.15786, 
    10.32381, 10.48983, 10.65592, 10.82209, 10.98833, 11.15463, 11.32101, 
    11.48746, 11.65396, 11.82054, 11.98717, 12.15387, 12.32062, 12.48743, 
    12.65429, 12.82121, 12.98818, 13.15521, 13.32228, 13.4894, 13.65656, 
    13.82376, 13.99101, 14.1583, 14.32563, 14.493, 14.6604, 14.82783, 
    14.9953, 15.1628, 15.33032, 15.49788, 15.66546, 15.83306, 16.00068, 
    16.16833, 16.33599, 16.50367, 16.67136, 16.83907, 17.00679, 17.17452, 
    17.34226, 17.51001, 17.67776, 17.84551, 18.01327, 18.18102, 18.34878, 
    18.51653, 18.68427, 18.85201, 19.01974, 19.18746, 19.35516, 19.52286, 
    19.69053, 19.85819, 20.02584, 20.19345, 20.36105, 20.52863, 20.69618, 
    20.8637, 21.03119, 21.19865, 21.36608, 21.53348, 21.70084, 21.86816, 
    22.03544, 22.20269, 22.36989, 22.53704, 22.70415, 22.87122, 23.03823, 
    23.20519, 23.3721, 23.53896, 23.70576, 23.87251, 24.03919, 24.20582, 
    24.37238, 24.53888, 24.70531, 24.87168, 25.03798, 25.2042, 25.37036, 
    25.53644, 25.70245, 25.86838, 26.03423, 26.20001, 26.3657, 26.53131, 
    26.69683, 26.86227, 27.02762, 27.19289, 27.35806, 27.52314, 27.68813, 
    27.85302, 28.01782, 28.18251, 28.34711, 28.51161, 28.67601, 28.8403, 
    29.00448, 29.16856, 29.33253, 29.4964, 29.66015, 29.82378, 29.98731, 
    30.15072, 30.31401, 30.47718, 30.64024, 30.80317, 30.96599, 31.12868, 
    31.29124, 31.45368, 31.61599, 31.77817, 31.94022, 32.10214, 32.26393, 
    32.42558, 32.5871, 32.74848, 32.90972, 33.07083, 33.23179, 33.39261, 
    33.5533, 33.71383, 33.87422, 34.03447, 34.19456, 34.35451, 34.51431, 
    34.67395, 34.83345, 34.99279, 35.15198, 35.31101, 35.46989, 35.6286, 
    35.78716, 35.94556, 36.1038, 36.26188, 36.41978, 36.57753, 36.73512, 
    36.89253, 37.04978, 37.20686, 37.36378, 37.52052, 37.67709, 37.83349, 
    37.98971, 38.14576, 38.30164, 38.45734, 38.61287, 38.76821, 38.92338, 
    39.07837, 39.23317, 39.3878, 39.54225, 39.69651, 39.85059, 40.00448, 
    40.15819, 40.31171, 40.46505, 40.61819, 40.77115, 40.92392, 41.0765, 
    41.22889, 41.38108, 41.53309, 41.6849, 41.83652, 41.98795, 42.13918, 
    42.29021, 42.44105, 42.59169, 42.74213, 42.89238, 43.04242, 43.19227, 
    43.34192, 43.49136, 43.6406, 43.78965, 43.93849, 44.08712, 44.23556, 
    44.38379, 44.53181, 44.67963, 44.82725, 44.97466, 45.12186, 45.26886, 
    45.41564,
  -22.17682, -22.05005, -21.92307, -21.79586, -21.66844, -21.5408, -21.41294, 
    -21.28487, -21.15657, -21.02806, -20.89933, -20.77038, -20.64121, 
    -20.51182, -20.38221, -20.25239, -20.12234, -19.99207, -19.86159, 
    -19.73088, -19.59996, -19.46881, -19.33744, -19.20586, -19.07405, 
    -18.94202, -18.80977, -18.67731, -18.54462, -18.41171, -18.27857, 
    -18.14522, -18.01165, -17.87785, -17.74384, -17.6096, -17.47514, 
    -17.34047, -17.20557, -17.07044, -16.9351, -16.79954, -16.66376, 
    -16.52775, -16.39152, -16.25508, -16.11841, -15.98152, -15.84441, 
    -15.70708, -15.56953, -15.43176, -15.29377, -15.15555, -15.01712, 
    -14.87847, -14.7396, -14.6005, -14.46119, -14.32166, -14.18191, 
    -14.04194, -13.90175, -13.76134, -13.62071, -13.47987, -13.3388, 
    -13.19752, -13.05602, -12.91431, -12.77237, -12.63022, -12.48785, 
    -12.34526, -12.20246, -12.05944, -11.91621, -11.77276, -11.6291, 
    -11.48522, -11.34112, -11.19681, -11.05229, -10.90756, -10.76261, 
    -10.61745, -10.47207, -10.32649, -10.18069, -10.03468, -9.888458, 
    -9.742028, -9.595387, -9.448537, -9.301478, -9.15421, -9.006734, 
    -8.859051, -8.71116, -8.563062, -8.414758, -8.266248, -8.117534, 
    -7.968614, -7.81949, -7.670163, -7.520633, -7.370901, -7.220967, 
    -7.070831, -6.920495, -6.769959, -6.619224, -6.468289, -6.317157, 
    -6.165827, -6.014301, -5.862578, -5.71066, -5.558547, -5.40624, -5.25374, 
    -5.101048, -4.948163, -4.795087, -4.641821, -4.488366, -4.334722, 
    -4.180889, -4.026869, -3.872663, -3.718271, -3.563694, -3.408934, 
    -3.25399, -3.098864, -2.943557, -2.788069, -2.632402, -2.476556, 
    -2.320532, -2.16433, -2.007954, -1.851402, -1.694676, -1.537776, 
    -1.380705, -1.223462, -1.066049, -0.9084675, -0.7507172, -0.5927998, 
    -0.4347162, -0.2764675, -0.1180547, 0.04052117, 0.199259, 0.3581576, 
    0.517216, 0.6764332, 0.8358079, 0.9953392, 1.155026, 1.314866, 1.47486, 
    1.635006, 1.795302, 1.955748, 2.116343, 2.277085, 2.437972, 2.599005, 
    2.76018, 2.921499, 3.082958, 3.244557, 3.406295, 3.56817, 3.730181, 
    3.892327, 4.054607, 4.217018, 4.37956, 4.542233, 4.705033, 4.867959, 
    5.031012, 5.194189, 5.357488, 5.520909, 5.68445, 5.84811, 6.011887, 
    6.175779, 6.339786, 6.503906, 6.668138, 6.83248, 6.996931, 7.161489, 
    7.326153, 7.490921, 7.655792, 7.820764, 7.985837, 8.151008, 8.316275, 
    8.481638, 8.647095, 8.812644, 8.978285, 9.144014, 9.309832, 9.475735, 
    9.641723, 9.807795, 9.973948, 10.14018, 10.30649, 10.47288, 10.63934, 
    10.80588, 10.97249, 11.13917, 11.30592, 11.47273, 11.63961, 11.80656, 
    11.97357, 12.14063, 12.30776, 12.47495, 12.64219, 12.80948, 12.97683, 
    13.14422, 13.31167, 13.47917, 13.64671, 13.81429, 13.98192, 14.14958, 
    14.31729, 14.48503, 14.65281, 14.82063, 14.98848, 15.15635, 15.32426, 
    15.49219, 15.66015, 15.82813, 15.99614, 16.16416, 16.33221, 16.50027, 
    16.66834, 16.83643, 17.00454, 17.17265, 17.34077, 17.50889, 17.67703, 
    17.84516, 18.0133, 18.18143, 18.34957, 18.5177, 18.68583, 18.85395, 
    19.02206, 19.19016, 19.35824, 19.52632, 19.69438, 19.86242, 20.03044, 
    20.19844, 20.36642, 20.53437, 20.7023, 20.8702, 21.03808, 21.20592, 
    21.37373, 21.5415, 21.70924, 21.87694, 22.0446, 22.21222, 22.3798, 
    22.54733, 22.71482, 22.88226, 23.04965, 23.21699, 23.38427, 23.5515, 
    23.71868, 23.8858, 24.05286, 24.21985, 24.38679, 24.55366, 24.72046, 
    24.8872, 25.05387, 25.22047, 25.38699, 25.55345, 25.71982, 25.88612, 
    26.05234, 26.21848, 26.38454, 26.55051, 26.7164, 26.88221, 27.04792, 
    27.21355, 27.37908, 27.54453, 27.70988, 27.87513, 28.04028, 28.20534, 
    28.37029, 28.53515, 28.6999, 28.86455, 29.02909, 29.19352, 29.35785, 
    29.52206, 29.68616, 29.85015, 30.01403, 30.17779, 30.34143, 30.50495, 
    30.66835, 30.83163, 30.99479, 31.15782, 31.32073, 31.48351, 31.64616, 
    31.80868, 31.97107, 32.13333, 32.29546, 32.45744, 32.6193, 32.78101, 
    32.94259, 33.10403, 33.26532, 33.42648, 33.58749, 33.74835, 33.90907, 
    34.06964, 34.23006, 34.39034, 34.55046, 34.71043, 34.87024, 35.02991, 
    35.18941, 35.34876, 35.50795, 35.66699, 35.82586, 35.98457, 36.14312, 
    36.30151, 36.45973, 36.61779, 36.77568, 36.93341, 37.09096, 37.24835, 
    37.40556, 37.56261, 37.71948, 37.87618, 38.0327, 38.18905, 38.34522, 
    38.50122, 38.65704, 38.81268, 38.96814, 39.12341, 39.27851, 39.43343, 
    39.58816, 39.74271, 39.89707, 40.05125, 40.20523, 40.35904, 40.51265, 
    40.66608, 40.81931, 40.97236, 41.12521, 41.27788, 41.43035, 41.58262, 
    41.7347, 41.88659, 42.03828, 42.18978, 42.34108, 42.49218, 42.64308, 
    42.79379, 42.94429, 43.09459, 43.2447, 43.3946, 43.5443, 43.6938, 
    43.84309, 43.99218, 44.14107, 44.28975, 44.43823, 44.5865, 44.73457, 
    44.88243, 45.03008, 45.17752, 45.32475, 45.47178,
  -22.25005, -22.12315, -21.99603, -21.86869, -21.74113, -21.61336, 
    -21.48537, -21.35715, -21.22872, -21.10007, -20.9712, -20.84211, 
    -20.7128, -20.58327, -20.45352, -20.32355, -20.19336, -20.06294, 
    -19.93231, -19.80145, -19.67038, -19.53908, -19.40756, -19.27582, 
    -19.14386, -19.01168, -18.87927, -18.74664, -18.6138, -18.48072, 
    -18.34743, -18.21392, -18.08018, -17.94622, -17.81204, -17.67764, 
    -17.54301, -17.40816, -17.27309, -17.1378, -17.00229, -16.86655, 
    -16.73059, -16.59441, -16.45801, -16.32138, -16.18453, -16.04746, 
    -15.91017, -15.77266, -15.63492, -15.49697, -15.35879, -15.22039, 
    -15.08177, -14.94292, -14.80386, -14.66457, -14.52507, -14.38534, 
    -14.24539, -14.10523, -13.96484, -13.82423, -13.6834, -13.54235, 
    -13.40108, -13.2596, -13.11789, -12.97597, -12.83382, -12.69146, 
    -12.54888, -12.40608, -12.26307, -12.11983, -11.97639, -11.83272, 
    -11.68884, -11.54473, -11.40042, -11.25589, -11.11114, -10.96618, 
    -10.82101, -10.67562, -10.53001, -10.3842, -10.23817, -10.09193, 
    -9.945474, -9.798808, -9.651931, -9.504843, -9.357545, -9.210037, 
    -9.06232, -8.914392, -8.766258, -8.617915, -8.469364, -8.320607, 
    -8.171643, -8.022473, -7.873098, -7.723518, -7.573734, -7.423746, 
    -7.273555, -7.123161, -6.972566, -6.821769, -6.670772, -6.519575, 
    -6.368178, -6.216583, -6.064789, -5.912798, -5.760611, -5.608228, 
    -5.455649, -5.302876, -5.149909, -4.996748, -4.843396, -4.689852, 
    -4.536117, -4.382192, -4.228077, -4.073774, -3.919284, -3.764606, 
    -3.609743, -3.454695, -3.299462, -3.144045, -2.988446, -2.832666, 
    -2.676704, -2.520563, -2.364242, -2.207744, -2.051068, -1.894216, 
    -1.737189, -1.579987, -1.422612, -1.265065, -1.107346, -0.9494573, 
    -0.7913989, -0.6331722, -0.4747781, -0.3162178, -0.1574923, 0.001397389, 
    0.1604501, 0.3196649, 0.4790405, 0.6385759, 0.79827, 0.9581217, 1.11813, 
    1.278293, 1.438611, 1.599081, 1.759704, 1.920477, 2.081399, 2.24247, 
    2.403687, 2.565051, 2.726559, 2.88821, 3.050004, 3.211938, 3.374012, 
    3.536224, 3.698573, 3.861058, 4.023677, 4.18643, 4.349314, 4.512329, 
    4.675472, 4.838744, 5.002142, 5.165665, 5.329312, 5.493081, 5.656971, 
    5.82098, 5.985108, 6.149352, 6.313712, 6.478185, 6.642771, 6.807468, 
    6.972274, 7.137189, 7.30221, 7.467336, 7.632566, 7.797898, 7.96333, 
    8.128862, 8.294492, 8.460217, 8.626038, 8.79195, 8.957955, 9.12405, 
    9.290233, 9.456503, 9.622858, 9.789297, 9.955818, 10.12242, 10.2891, 
    10.45586, 10.62269, 10.7896, 10.95658, 11.12363, 11.29075, 11.45794, 
    11.6252, 11.79252, 11.9599, 12.12734, 12.29484, 12.46241, 12.63002, 
    12.79769, 12.96542, 13.13319, 13.30102, 13.46889, 13.63681, 13.80477, 
    13.97278, 14.14083, 14.30891, 14.47704, 14.6452, 14.81339, 14.98162, 
    15.14988, 15.31817, 15.48648, 15.65482, 15.82319, 15.99157, 16.15998, 
    16.32841, 16.49685, 16.66531, 16.83378, 17.00227, 17.17076, 17.33926, 
    17.50777, 17.67629, 17.84481, 18.01333, 18.18185, 18.35037, 18.51888, 
    18.68739, 18.85589, 19.02439, 19.19287, 19.36134, 19.5298, 19.69824, 
    19.86666, 20.03506, 20.20345, 20.37181, 20.54015, 20.70846, 20.87674, 
    21.04499, 21.21321, 21.3814, 21.54956, 21.71768, 21.88576, 22.0538, 
    22.2218, 22.38976, 22.55767, 22.72553, 22.89335, 23.06112, 23.22883, 
    23.3965, 23.5641, 23.73166, 23.89915, 24.06658, 24.23396, 24.40126, 
    24.56851, 24.73569, 24.9028, 25.06984, 25.23681, 25.4037, 25.57052, 
    25.73727, 25.90394, 26.07053, 26.23704, 26.40346, 26.5698, 26.73606, 
    26.90223, 27.06831, 27.2343, 27.4002, 27.566, 27.73171, 27.89733, 
    28.06285, 28.22826, 28.39358, 28.55879, 28.7239, 28.8889, 29.0538, 
    29.21859, 29.38327, 29.54784, 29.7123, 29.87664, 30.04086, 30.20497, 
    30.36896, 30.53283, 30.69658, 30.86021, 31.02371, 31.18709, 31.35034, 
    31.51347, 31.67646, 31.83932, 32.00206, 32.16465, 32.32712, 32.48944, 
    32.65163, 32.81369, 32.9756, 33.13737, 33.299, 33.46048, 33.62183, 
    33.78302, 33.94407, 34.10497, 34.26571, 34.42631, 34.58676, 34.74705, 
    34.90719, 35.06717, 35.227, 35.38667, 35.54618, 35.70553, 35.86472, 
    36.02375, 36.18261, 36.34131, 36.49984, 36.65821, 36.81641, 36.97445, 
    37.13231, 37.29, 37.44752, 37.60487, 37.76204, 37.91904, 38.07586, 
    38.23251, 38.38898, 38.54527, 38.70139, 38.85732, 39.01307, 39.16864, 
    39.32403, 39.47923, 39.63425, 39.78909, 39.94373, 40.09819, 40.25247, 
    40.40655, 40.56045, 40.71415, 40.86767, 41.02099, 41.17412, 41.32705, 
    41.4798, 41.63235, 41.7847, 41.93686, 42.08881, 42.24058, 42.39214, 
    42.54351, 42.69467, 42.84563, 42.9964, 43.14697, 43.29733, 43.44749, 
    43.59744, 43.74719, 43.89674, 44.04608, 44.19522, 44.34415, 44.49288, 
    44.6414, 44.7897, 44.93781, 45.0857, 45.23338, 45.38086, 45.52813,
  -22.32348, -22.19645, -22.0692, -21.94173, -21.81404, -21.68614, -21.55801, 
    -21.42966, -21.30109, -21.1723, -21.04329, -20.91406, -20.78461, 
    -20.65494, -20.52504, -20.39492, -20.26459, -20.13403, -20.00324, 
    -19.87224, -19.74101, -19.60957, -19.4779, -19.346, -19.21389, -19.08155, 
    -18.94899, -18.8162, -18.68319, -18.54996, -18.41651, -18.28283, 
    -18.14893, -18.01481, -17.88046, -17.74589, -17.6111, -17.47608, 
    -17.34084, -17.20538, -17.06969, -16.93378, -16.79765, -16.66129, 
    -16.52471, -16.3879, -16.25088, -16.11363, -15.97615, -15.83846, 
    -15.70054, -15.56239, -15.42403, -15.28544, -15.14663, -15.0076, 
    -14.86834, -14.72886, -14.58916, -14.44924, -14.3091, -14.16873, 
    -14.02814, -13.88733, -13.7463, -13.60505, -13.46358, -13.32189, 
    -13.17998, -13.03784, -12.89549, -12.75292, -12.61013, -12.46712, 
    -12.32389, -12.18044, -12.03677, -11.89289, -11.74879, -11.60447, 
    -11.45993, -11.31518, -11.17021, -11.02502, -10.87962, -10.734, 
    -10.58817, -10.44212, -10.29586, -10.14939, -10.0027, -9.855797, 
    -9.708683, -9.561357, -9.413819, -9.26607, -9.118111, -8.969941, 
    -8.821562, -8.672973, -8.524176, -8.37517, -8.225956, -8.076535, 
    -7.926908, -7.777074, -7.627035, -7.476791, -7.326343, -7.175691, 
    -7.024836, -6.873778, -6.722518, -6.571057, -6.419395, -6.267534, 
    -6.115473, -5.963213, -5.810756, -5.658101, -5.50525, -5.352202, 
    -5.19896, -5.045524, -4.891893, -4.73807, -4.584055, -4.429849, 
    -4.275452, -4.120865, -3.966089, -3.811126, -3.655975, -3.500638, 
    -3.345114, -3.189407, -3.033515, -2.877441, -2.721185, -2.564747, 
    -2.408129, -2.251332, -2.094357, -1.937204, -1.779874, -1.62237, 
    -1.46469, -1.306837, -1.148812, -0.9906146, -0.832247, -0.6737099, 
    -0.5150044, -0.3561315, -0.1970922, -0.03788763, 0.1214811, 0.281013, 
    0.4407069, 0.6005618, 0.7605764, 0.9207497, 1.08108, 1.241568, 1.40221, 
    1.563007, 1.723956, 1.885057, 2.046308, 2.207709, 2.369258, 2.530954, 
    2.692795, 2.854781, 3.01691, 3.17918, 3.341591, 3.504142, 3.66683, 
    3.829655, 3.992616, 4.155711, 4.318938, 4.482297, 4.645786, 4.809403, 
    4.973148, 5.137019, 5.301014, 5.465133, 5.629373, 5.793734, 5.958214, 
    6.122811, 6.287525, 6.452353, 6.617294, 6.782348, 6.947511, 7.112783, 
    7.278163, 7.443649, 7.609239, 7.774932, 7.940726, 8.106621, 8.272614, 
    8.438703, 8.604887, 8.771166, 8.937536, 9.103998, 9.270549, 9.437186, 
    9.60391, 9.770719, 9.93761, 10.10458, 10.27163, 10.43876, 10.60597, 
    10.77325, 10.9406, 11.10803, 11.27553, 11.44309, 11.61072, 11.77841, 
    11.94617, 12.11399, 12.28187, 12.44981, 12.61781, 12.78586, 12.95396, 
    13.12211, 13.29032, 13.45857, 13.62687, 13.79521, 13.9636, 14.13203, 
    14.3005, 14.469, 14.63755, 14.80612, 14.97473, 15.14338, 15.31205, 
    15.48074, 15.64947, 15.81822, 15.98699, 16.15578, 16.32459, 16.49342, 
    16.66226, 16.83112, 16.99999, 17.16887, 17.33776, 17.50665, 17.67555, 
    17.84445, 18.01336, 18.18226, 18.35117, 18.52007, 18.68896, 18.85785, 
    19.02673, 19.19559, 19.36445, 19.53329, 19.70211, 19.87092, 20.03971, 
    20.20848, 20.37722, 20.54594, 20.71464, 20.8833, 21.05194, 21.22054, 
    21.38912, 21.55765, 21.72615, 21.89462, 22.06304, 22.23142, 22.39976, 
    22.56805, 22.73629, 22.90449, 23.07264, 23.24073, 23.40877, 23.57676, 
    23.74469, 23.91256, 24.08037, 24.24812, 24.4158, 24.58342, 24.75097, 
    24.91846, 25.08587, 25.25322, 25.42048, 25.58768, 25.7548, 25.92184, 
    26.08879, 26.25567, 26.42247, 26.58918, 26.7558, 26.92234, 27.08879, 
    27.25514, 27.42141, 27.58758, 27.75365, 27.91963, 28.08551, 28.25129, 
    28.41696, 28.58253, 28.748, 28.91337, 29.07862, 29.24377, 29.4088, 
    29.57373, 29.73854, 29.90323, 30.06781, 30.23227, 30.39661, 30.56084, 
    30.72494, 30.88891, 31.05276, 31.21649, 31.38008, 31.54355, 31.70689, 
    31.8701, 32.03317, 32.19611, 32.35891, 32.52158, 32.68411, 32.8465, 
    33.00875, 33.17085, 33.33282, 33.49463, 33.65631, 33.81783, 33.97921, 
    34.14044, 34.30151, 34.46244, 34.62321, 34.78383, 34.94429, 35.1046, 
    35.26475, 35.42474, 35.58456, 35.74423, 35.90374, 36.06308, 36.22226, 
    36.38128, 36.54012, 36.6988, 36.85731, 37.01565, 37.17382, 37.33182, 
    37.48964, 37.6473, 37.80477, 37.96207, 38.1192, 38.27615, 38.43291, 
    38.5895, 38.74591, 38.90214, 39.05819, 39.21405, 39.36973, 39.52522, 
    39.68053, 39.83565, 39.99059, 40.14533, 40.29989, 40.45425, 40.60843, 
    40.76242, 40.91621, 41.06981, 41.22321, 41.37643, 41.52944, 41.68226, 
    41.83488, 41.98731, 42.13954, 42.29157, 42.4434, 42.59503, 42.74646, 
    42.89769, 43.04871, 43.19954, 43.35015, 43.50057, 43.65078, 43.80079, 
    43.95059, 44.10019, 44.24957, 44.39875, 44.54773, 44.69649, 44.84505, 
    44.99339, 45.14153, 45.28946, 45.43717, 45.58467,
  -22.39713, -22.26997, -22.14259, -22.01499, -21.88717, -21.75913, 
    -21.63087, -21.50238, -21.37368, -21.24475, -21.1156, -20.98623, 
    -20.85663, -20.72682, -20.59678, -20.46652, -20.33604, -20.20533, 
    -20.0744, -19.94325, -19.81187, -19.68027, -19.54845, -19.4164, 
    -19.28413, -19.15164, -19.01892, -18.88598, -18.75281, -18.61942, 
    -18.48581, -18.35197, -18.2179, -18.08362, -17.9491, -17.81437, 
    -17.67941, -17.54422, -17.40881, -17.27317, -17.13731, -17.00123, 
    -16.86492, -16.72839, -16.59163, -16.45465, -16.31744, -16.18001, 
    -16.04235, -15.90447, -15.76637, -15.62804, -15.48949, -15.35071, 
    -15.21171, -15.07249, -14.93304, -14.79337, -14.65347, -14.51336, 
    -14.37302, -14.23245, -14.09167, -13.95066, -13.80943, -13.66797, 
    -13.5263, -13.3844, -13.24228, -13.09994, -12.95738, -12.8146, -12.67159, 
    -12.52837, -12.38492, -12.24126, -12.09738, -11.95327, -11.80895, 
    -11.66441, -11.51965, -11.37468, -11.22948, -11.08407, -10.93844, 
    -10.7926, -10.64653, -10.50026, -10.35376, -10.20706, -10.06013, 
    -9.912995, -9.765644, -9.61808, -9.470303, -9.322312, -9.17411, 
    -9.025697, -8.877072, -8.728237, -8.579192, -8.429937, -8.280474, 
    -8.130801, -7.980921, -7.830834, -7.680539, -7.530039, -7.379333, 
    -7.228421, -7.077305, -6.925986, -6.774463, -6.622737, -6.47081, 
    -6.318682, -6.166353, -6.013824, -5.861095, -5.708169, -5.555044, 
    -5.401722, -5.248204, -5.09449, -4.940582, -4.786479, -4.632183, 
    -4.477694, -4.323014, -4.168142, -4.013081, -3.85783, -3.702391, 
    -3.546764, -3.39095, -3.23495, -3.078765, -2.922396, -2.765844, -2.60911, 
    -2.452193, -2.295097, -2.137821, -1.980366, -1.822734, -1.664925, 
    -1.50694, -1.34878, -1.190447, -1.031941, -0.8732628, -0.7144144, 
    -0.5553964, -0.3962098, -0.2368557, -0.07733514, 0.08235074, 0.2422009, 
    0.4022142, 0.5623895, 0.7227257, 0.8832217, 1.043876, 1.204688, 1.365657, 
    1.52678, 1.688058, 1.849488, 2.01107, 2.172802, 2.334684, 2.496713, 
    2.658889, 2.82121, 2.983675, 3.146283, 3.309033, 3.471923, 3.634952, 
    3.798119, 3.961422, 4.12486, 4.288432, 4.452136, 4.615972, 4.779936, 
    4.944029, 5.108249, 5.272595, 5.437064, 5.601656, 5.76637, 5.931203, 
    6.096155, 6.261224, 6.426408, 6.591707, 6.757118, 6.92264, 7.088272, 
    7.254012, 7.419858, 7.58581, 7.751866, 7.918024, 8.084282, 8.250639, 
    8.417094, 8.583645, 8.75029, 8.917028, 9.083858, 9.250777, 9.417785, 
    9.584879, 9.752058, 9.91932, 10.08666, 10.25409, 10.42159, 10.58917, 
    10.75683, 10.92456, 11.09236, 11.26023, 11.42817, 11.59618, 11.76425, 
    11.93238, 12.10058, 12.26884, 12.43716, 12.60553, 12.77396, 12.94245, 
    13.11098, 13.27957, 13.4482, 13.61689, 13.78561, 13.95438, 14.12319, 
    14.29204, 14.46093, 14.62986, 14.79882, 14.96782, 15.13684, 15.3059, 
    15.47498, 15.64409, 15.81322, 15.98238, 16.15156, 16.32076, 16.48997, 
    16.6592, 16.82844, 16.9977, 17.16697, 17.33624, 17.50552, 17.67481, 
    17.8441, 18.01339, 18.18268, 18.35197, 18.52126, 18.69054, 18.85981, 
    19.02908, 19.19833, 19.36757, 19.5368, 19.70601, 19.8752, 20.04438, 
    20.21353, 20.38266, 20.55177, 20.72085, 20.8899, 21.05892, 21.22791, 
    21.39686, 21.56578, 21.73467, 21.90351, 22.07232, 22.24108, 22.4098, 
    22.57847, 22.7471, 22.91568, 23.08421, 23.25268, 23.4211, 23.58947, 
    23.75778, 23.92603, 24.09422, 24.26234, 24.4304, 24.5984, 24.76633, 
    24.93419, 25.10198, 25.2697, 25.43734, 25.60491, 25.7724, 25.93981, 
    26.10714, 26.27439, 26.44156, 26.60864, 26.77563, 26.94254, 27.10935, 
    27.27608, 27.44271, 27.60924, 27.77568, 27.94202, 28.10827, 28.27441, 
    28.44045, 28.60638, 28.77221, 28.93793, 29.10355, 29.26905, 29.43445, 
    29.59973, 29.76489, 29.92994, 30.09488, 30.25969, 30.42439, 30.58896, 
    30.75341, 30.91774, 31.08194, 31.24601, 31.40995, 31.57377, 31.73745, 
    31.901, 32.06442, 32.2277, 32.39085, 32.55385, 32.71672, 32.87945, 
    33.04203, 33.20448, 33.36678, 33.52893, 33.69093, 33.85279, 34.0145, 
    34.17606, 34.33746, 34.49872, 34.65982, 34.82076, 34.98155, 35.14218, 
    35.30265, 35.46296, 35.62311, 35.7831, 35.94292, 36.10258, 36.26207, 
    36.4214, 36.58056, 36.73955, 36.89837, 37.05703, 37.2155, 37.37381, 
    37.53194, 37.6899, 37.84768, 38.00528, 38.16271, 38.31996, 38.47703, 
    38.63391, 38.79062, 38.94714, 39.10349, 39.25964, 39.41561, 39.57139, 
    39.72699, 39.8824, 40.03762, 40.19265, 40.3475, 40.50214, 40.6566, 
    40.81087, 40.96494, 41.11882, 41.2725, 41.42599, 41.57928, 41.73237, 
    41.88527, 42.03796, 42.19046, 42.34276, 42.49486, 42.64675, 42.79845, 
    42.94994, 43.10122, 43.25231, 43.40319, 43.55386, 43.70433, 43.85459, 
    44.00464, 44.15449, 44.30413, 44.45356, 44.60278, 44.75179, 44.9006, 
    45.04919, 45.19757, 45.34574, 45.49369, 45.64144,
  -22.471, -22.34371, -22.2162, -22.08847, -21.96052, -21.83234, -21.70394, 
    -21.57532, -21.44648, -21.31741, -21.18813, -21.05861, -20.92888, 
    -20.79892, -20.66874, -20.53834, -20.40771, -20.27685, -20.14578, 
    -20.01447, -19.88295, -19.7512, -19.61922, -19.48702, -19.3546, 
    -19.22195, -19.08908, -18.95598, -18.82265, -18.6891, -18.55532, 
    -18.42132, -18.2871, -18.15265, -18.01797, -17.88306, -17.74793, 
    -17.61258, -17.477, -17.34119, -17.20516, -17.0689, -16.93242, -16.79571, 
    -16.65877, -16.52161, -16.38422, -16.24661, -16.10877, -15.97071, 
    -15.83242, -15.69391, -15.55517, -15.4162, -15.27701, -15.1376, 
    -14.99796, -14.8581, -14.71801, -14.57769, -14.43716, -14.2964, 
    -14.15541, -14.0142, -13.87277, -13.73111, -13.58923, -13.44713, 
    -13.3048, -13.16225, -13.01948, -12.87649, -12.73327, -12.58984, 
    -12.44618, -12.3023, -12.1582, -12.01388, -11.86934, -11.72457, 
    -11.57959, -11.43439, -11.28897, -11.14334, -10.99748, -10.85141, 
    -10.70511, -10.55861, -10.41188, -10.26494, -10.11778, -9.970406, 
    -9.822817, -9.675014, -9.526996, -9.378764, -9.230319, -9.081662, 
    -8.932792, -8.78371, -8.634417, -8.484912, -8.335197, -8.185273, 
    -8.03514, -7.884798, -7.734248, -7.583489, -7.432525, -7.281354, 
    -7.129977, -6.978395, -6.826608, -6.674618, -6.522424, -6.370028, 
    -6.21743, -6.064631, -5.911631, -5.758432, -5.605033, -5.451436, 
    -5.297641, -5.14365, -4.989462, -4.835079, -4.680501, -4.52573, 
    -4.370765, -4.215608, -4.06026, -3.904721, -3.748992, -3.593075, 
    -3.43697, -3.280677, -3.124198, -2.967533, -2.810684, -2.653652, 
    -2.496437, -2.33904, -2.181462, -2.023704, -1.865768, -1.707653, 
    -1.549362, -1.390895, -1.232253, -1.073437, -0.9144477, -0.7552869, 
    -0.5959553, -0.436454, -0.276784, -0.1169464, 0.04305766, 0.2032271, 
    0.3635609, 0.5240578, 0.6847168, 0.8455366, 1.006516, 1.167654, 1.32895, 
    1.490402, 1.652009, 1.813769, 1.975683, 2.137748, 2.299963, 2.462327, 
    2.624838, 2.787496, 2.950299, 3.113246, 3.276336, 3.439567, 3.602938, 
    3.766448, 3.930094, 4.093877, 4.257795, 4.421846, 4.586029, 4.750342, 
    4.914785, 5.079356, 5.244052, 5.408875, 5.57382, 5.738887, 5.904076, 
    6.069384, 6.234809, 6.400351, 6.566008, 6.731778, 6.89766, 7.063653, 
    7.229754, 7.395964, 7.562279, 7.728698, 7.895221, 8.061845, 8.228568, 
    8.39539, 8.562308, 8.729322, 8.89643, 9.063629, 9.230919, 9.398297, 
    9.565763, 9.733315, 9.90095, 10.06867, 10.23647, 10.40434, 10.5723, 
    10.74033, 10.90844, 11.07661, 11.24486, 11.41318, 11.58157, 11.75002, 
    11.91854, 12.08711, 12.25575, 12.42445, 12.59321, 12.76202, 12.93089, 
    13.0998, 13.26877, 13.43779, 13.60686, 13.77597, 13.94512, 14.11432, 
    14.28355, 14.45283, 14.62214, 14.79149, 14.96087, 15.13028, 15.29972, 
    15.46919, 15.63869, 15.80821, 15.97775, 16.14732, 16.3169, 16.48651, 
    16.65612, 16.82576, 16.9954, 17.16505, 17.33472, 17.50439, 17.67406, 
    17.84374, 18.01342, 18.1831, 18.35278, 18.52245, 18.69212, 18.86178, 
    19.03144, 19.20108, 19.37071, 19.54032, 19.70992, 19.8795, 20.04907, 
    20.21861, 20.38812, 20.55762, 20.72708, 20.89652, 21.06593, 21.2353, 
    21.40464, 21.57395, 21.74322, 21.91245, 22.08164, 22.25079, 22.41989, 
    22.58895, 22.75796, 22.92692, 23.09583, 23.26469, 23.43349, 23.60224, 
    23.77093, 23.93956, 24.10813, 24.27663, 24.44507, 24.61345, 24.78176, 
    24.94999, 25.11816, 25.28625, 25.45427, 25.62222, 25.79008, 25.95787, 
    26.12557, 26.2932, 26.46073, 26.62819, 26.79555, 26.96283, 27.13001, 
    27.2971, 27.4641, 27.631, 27.79781, 27.96452, 28.13113, 28.29763, 
    28.46404, 28.63033, 28.79653, 28.96261, 29.12859, 29.29445, 29.46021, 
    29.62584, 29.79137, 29.95677, 30.12206, 30.28723, 30.45228, 30.61721, 
    30.78201, 30.94669, 31.11124, 31.27566, 31.43995, 31.60411, 31.76814, 
    31.93204, 32.0958, 32.25943, 32.42291, 32.58626, 32.74947, 32.91254, 
    33.07546, 33.23824, 33.40088, 33.56337, 33.72571, 33.8879, 34.04994, 
    34.21183, 34.37357, 34.53515, 34.69658, 34.85785, 35.01896, 35.17991, 
    35.34071, 35.50134, 35.66181, 35.82212, 35.98226, 36.14224, 36.30205, 
    36.4617, 36.62117, 36.78048, 36.93961, 37.09857, 37.25736, 37.41597, 
    37.57441, 37.73268, 37.89076, 38.04867, 38.2064, 38.36395, 38.52132, 
    38.6785, 38.83551, 38.99233, 39.14896, 39.30541, 39.46167, 39.61775, 
    39.77364, 39.92934, 40.08485, 40.24017, 40.39529, 40.55022, 40.70497, 
    40.85951, 41.01387, 41.16802, 41.32198, 41.47575, 41.62931, 41.78268, 
    41.93585, 42.08881, 42.24158, 42.39415, 42.54651, 42.69867, 42.85063, 
    43.00239, 43.15393, 43.30528, 43.45642, 43.60735, 43.75808, 43.90859, 
    44.0589, 44.209, 44.35889, 44.50858, 44.65805, 44.8073, 44.95636, 
    45.10519, 45.25381, 45.40223, 45.55042, 45.69841,
  -22.54509, -22.41767, -22.29003, -22.16217, -22.03408, -21.90577, 
    -21.77724, -21.64848, -21.5195, -21.3903, -21.26087, -21.13122, 
    -21.00135, -20.87125, -20.74092, -20.61037, -20.4796, -20.3486, 
    -20.21737, -20.08592, -19.95425, -19.82235, -19.69022, -19.55787, 
    -19.42529, -19.29249, -19.15945, -19.0262, -18.89271, -18.759, -18.62507, 
    -18.4909, -18.35651, -18.2219, -18.08705, -17.95198, -17.81668, 
    -17.68116, -17.54541, -17.40943, -17.27323, -17.1368, -17.00014, 
    -16.86325, -16.72614, -16.5888, -16.45123, -16.31344, -16.17542, 
    -16.03717, -15.8987, -15.76, -15.62107, -15.48192, -15.34254, -15.20294, 
    -15.0631, -14.92305, -14.78276, -14.64225, -14.50152, -14.36056, 
    -14.21937, -14.07796, -13.93633, -13.79447, -13.65238, -13.51008, 
    -13.36754, -13.22479, -13.08181, -12.9386, -12.79517, -12.65152, 
    -12.50765, -12.36355, -12.21924, -12.0747, -11.92994, -11.78495, 
    -11.63975, -11.49433, -11.34868, -11.20282, -11.05673, -10.91043, 
    -10.76391, -10.61717, -10.47021, -10.32303, -10.17564, -10.02803, 
    -9.880202, -9.73216, -9.5839, -9.435428, -9.286739, -9.137836, -8.988721, 
    -8.839392, -8.689849, -8.540095, -8.390129, -8.239953, -8.089565, 
    -7.938968, -7.788161, -7.637146, -7.485922, -7.33449, -7.182851, 
    -7.031006, -6.878956, -6.7267, -6.574239, -6.421575, -6.268707, 
    -6.115637, -5.962365, -5.808892, -5.655219, -5.501346, -5.347274, 
    -5.193004, -5.038536, -4.883872, -4.729012, -4.573956, -4.418707, 
    -4.263264, -4.107628, -3.9518, -3.795781, -3.639573, -3.483175, 
    -3.326588, -3.169814, -3.012853, -2.855706, -2.698375, -2.54086, 
    -2.383162, -2.225281, -2.06722, -1.908978, -1.750558, -1.591959, 
    -1.433183, -1.274231, -1.115104, -0.9558028, -0.7963286, -0.6366824, 
    -0.4768653, -0.3168784, -0.1567227, 0.003600628, 0.1640905, 0.3247459, 
    0.4855655, 0.6465483, 0.8076932, 0.9689989, 1.130464, 1.292088, 1.45387, 
    1.615807, 1.777899, 1.940145, 2.102544, 2.265094, 2.427794, 2.590642, 
    2.753639, 2.916781, 3.080068, 3.243499, 3.407072, 3.570786, 3.73464, 
    3.898632, 4.062761, 4.227026, 4.391425, 4.555957, 4.72062, 4.885414, 
    5.050336, 5.215386, 5.380562, 5.545862, 5.711285, 5.87683, 6.042495, 
    6.208279, 6.374179, 6.540196, 6.706327, 6.872571, 7.038926, 7.205391, 
    7.371964, 7.538644, 7.705429, 7.872317, 8.039309, 8.2064, 8.37359, 
    8.540878, 8.708261, 8.87574, 9.04331, 9.210972, 9.378723, 9.546563, 
    9.714488, 9.882499, 10.05059, 10.21877, 10.38702, 10.55535, 10.72376, 
    10.89225, 11.0608, 11.22943, 11.39813, 11.56689, 11.73573, 11.90462, 
    12.07358, 12.24261, 12.41169, 12.58083, 12.75002, 12.91927, 13.08857, 
    13.25793, 13.42733, 13.59678, 13.76628, 13.93582, 14.1054, 14.27502, 
    14.44469, 14.61439, 14.78412, 14.95389, 15.12369, 15.29352, 15.46338, 
    15.63326, 15.80317, 15.97311, 16.14306, 16.31304, 16.48303, 16.65303, 
    16.82306, 16.99309, 17.16313, 17.33319, 17.50325, 17.67331, 17.84338, 
    18.01345, 18.18352, 18.35359, 18.52365, 18.69371, 18.86377, 19.03381, 
    19.20384, 19.37386, 19.54386, 19.71385, 19.88382, 20.05377, 20.2237, 
    20.39361, 20.56349, 20.73335, 20.90317, 21.07297, 21.24273, 21.41246, 
    21.58215, 21.75181, 21.92143, 22.091, 22.26054, 22.43003, 22.59947, 
    22.76887, 22.93821, 23.10751, 23.27675, 23.44593, 23.61506, 23.78414, 
    23.95315, 24.1221, 24.29099, 24.45981, 24.62856, 24.79725, 24.96587, 
    25.13441, 25.30288, 25.47128, 25.6396, 25.80784, 25.976, 26.14408, 
    26.31208, 26.47999, 26.64782, 26.81556, 26.9832, 27.15076, 27.31822, 
    27.48559, 27.65286, 27.82004, 27.98711, 28.15409, 28.32096, 28.48773, 
    28.65439, 28.82095, 28.9874, 29.15373, 29.31996, 29.48607, 29.65207, 
    29.81795, 29.98372, 30.14936, 30.31489, 30.4803, 30.64557, 30.81073, 
    30.97576, 31.14066, 31.30544, 31.47008, 31.63459, 31.79897, 31.96321, 
    32.12732, 32.29129, 32.45512, 32.61881, 32.78236, 32.94577, 33.10904, 
    33.27216, 33.43513, 33.59795, 33.76063, 33.92316, 34.08553, 34.24775, 
    34.40982, 34.57173, 34.73349, 34.89509, 35.05653, 35.21781, 35.37893, 
    35.53988, 35.70068, 35.86131, 36.02177, 36.18207, 36.3422, 36.50216, 
    36.66195, 36.82157, 36.98101, 37.14029, 37.29939, 37.45831, 37.61706, 
    37.77563, 37.93402, 38.09224, 38.25027, 38.40812, 38.56579, 38.72327, 
    38.88058, 39.03769, 39.19463, 39.35137, 39.50793, 39.6643, 39.82047, 
    39.97646, 40.13226, 40.28786, 40.44328, 40.5985, 40.75352, 40.90835, 
    41.06298, 41.21742, 41.37166, 41.5257, 41.67954, 41.83318, 41.98663, 
    42.13986, 42.2929, 42.44574, 42.59837, 42.7508, 42.90302, 43.05504, 
    43.20685, 43.35846, 43.50986, 43.66105, 43.81203, 43.9628, 44.11337, 
    44.26372, 44.41386, 44.5638, 44.71352, 44.86303, 45.01232, 45.1614, 
    45.31027, 45.45893, 45.60737, 45.75559,
  -22.6194, -22.49185, -22.36408, -22.23608, -22.10786, -21.97942, -21.85075, 
    -21.72186, -21.59275, -21.46341, -21.33384, -21.20405, -21.07403, 
    -20.94379, -20.81332, -20.68263, -20.55171, -20.42057, -20.2892, 
    -20.1576, -20.02577, -19.89372, -19.76144, -19.62894, -19.4962, 
    -19.36325, -19.23006, -19.09664, -18.963, -18.82913, -18.69503, 
    -18.56071, -18.42616, -18.29137, -18.15636, -18.02113, -17.88566, 
    -17.74997, -17.61405, -17.4779, -17.34152, -17.20492, -17.06808, 
    -16.93102, -16.79373, -16.65621, -16.51847, -16.38049, -16.24229, 
    -16.10386, -15.9652, -15.82631, -15.6872, -15.54786, -15.40829, 
    -15.26849, -15.12847, -14.98822, -14.84774, -14.70704, -14.56611, 
    -14.42495, -14.28356, -14.14195, -14.00011, -13.85805, -13.71576, 
    -13.57325, -13.43051, -13.28754, -13.14435, -13.00093, -12.8573, 
    -12.71343, -12.56934, -12.42503, -12.2805, -12.13574, -11.99076, 
    -11.84555, -11.70013, -11.55448, -11.40861, -11.26252, -11.1162, 
    -10.96967, -10.82292, -10.67595, -10.52876, -10.38134, -10.23372, 
    -10.08587, -9.937801, -9.789518, -9.641019, -9.492303, -9.343371, 
    -9.194223, -9.044861, -8.895284, -8.745493, -8.595489, -8.445271, 
    -8.294841, -8.144198, -7.993346, -7.842282, -7.691008, -7.539525, 
    -7.387832, -7.235931, -7.083822, -6.931507, -6.778984, -6.626256, 
    -6.473323, -6.320185, -6.166843, -6.013299, -5.859551, -5.705603, 
    -5.551453, -5.397103, -5.242554, -5.087805, -4.932859, -4.777716, 
    -4.622376, -4.46684, -4.31111, -4.155186, -3.999069, -3.842759, 
    -3.686258, -3.529566, -3.372685, -3.215615, -3.058357, -2.900912, 
    -2.743281, -2.585464, -2.427464, -2.26928, -2.110914, -1.952366, 
    -1.793639, -1.634732, -1.475646, -1.316383, -1.156944, -0.9973296, 
    -0.8375409, -0.6775791, -0.5174451, -0.3571402, -0.1966653, -0.03602163, 
    0.1247898, 0.2857678, 0.4469113, 0.6082191, 0.7696902, 0.9313231, 
    1.093117, 1.25507, 1.417182, 1.579452, 1.741877, 1.904457, 2.06719, 
    2.230077, 2.393113, 2.5563, 2.719636, 2.883118, 3.046747, 3.21052, 
    3.374437, 3.538496, 3.702695, 3.867033, 4.03151, 4.196123, 4.360872, 
    4.525754, 4.690769, 4.855915, 5.021191, 5.186595, 5.352126, 5.517782, 
    5.683562, 5.849464, 6.015488, 6.181632, 6.347893, 6.514271, 6.680764, 
    6.847371, 7.01409, 7.18092, 7.347858, 7.514904, 7.682056, 7.849313, 
    8.016672, 8.184133, 8.351693, 8.519352, 8.687107, 8.854958, 9.022902, 
    9.190937, 9.359062, 9.527277, 9.695578, 9.863964, 10.03243, 10.20099, 
    10.36962, 10.53833, 10.70712, 10.87598, 11.04492, 11.21393, 11.38301, 
    11.55215, 11.72137, 11.89065, 12.05999, 12.2294, 12.39886, 12.56839, 
    12.73797, 12.90761, 13.07729, 13.24703, 13.41682, 13.58666, 13.75655, 
    13.92647, 14.09645, 14.26646, 14.43651, 14.6066, 14.77672, 14.94688, 
    15.11707, 15.28729, 15.45754, 15.62781, 15.79811, 15.96844, 16.13878, 
    16.30915, 16.47953, 16.64993, 16.82034, 16.99077, 17.16121, 17.33165, 
    17.5021, 17.67256, 17.84302, 18.01348, 18.18394, 18.3544, 18.52486, 
    18.69531, 18.86576, 19.03619, 19.20661, 19.37702, 19.54742, 19.7178, 
    19.88816, 20.0585, 20.22882, 20.39912, 20.56939, 20.73964, 20.90985, 
    21.08004, 21.25019, 21.42031, 21.59039, 21.76044, 21.93044, 22.10041, 
    22.27033, 22.44021, 22.61004, 22.77982, 22.94955, 23.11923, 23.28886, 
    23.45843, 23.62795, 23.7974, 23.9668, 24.13613, 24.3054, 24.47461, 
    24.64374, 24.81281, 24.98181, 25.15074, 25.31959, 25.48836, 25.65706, 
    25.82568, 25.99422, 26.16268, 26.33105, 26.49934, 26.66754, 26.83565, 
    27.00367, 27.1716, 27.33944, 27.50718, 27.67482, 27.84236, 28.00981, 
    28.17715, 28.34439, 28.51153, 28.67856, 28.84548, 29.01229, 29.17899, 
    29.34558, 29.51205, 29.67842, 29.84466, 30.01078, 30.17679, 30.34267, 
    30.50843, 30.67407, 30.83958, 31.00496, 31.17022, 31.33534, 31.50034, 
    31.6652, 31.82993, 31.99452, 32.15897, 32.32329, 32.48746, 32.6515, 
    32.8154, 32.97915, 33.14275, 33.30621, 33.46952, 33.63269, 33.7957, 
    33.95856, 34.12127, 34.28382, 34.44623, 34.60847, 34.77056, 34.93249, 
    35.09425, 35.25586, 35.41731, 35.57859, 35.73971, 35.90066, 36.06144, 
    36.22206, 36.38251, 36.54279, 36.70289, 36.86283, 37.02259, 37.18217, 
    37.34159, 37.50082, 37.65988, 37.81876, 37.97746, 38.13598, 38.29432, 
    38.45247, 38.61044, 38.76823, 38.92583, 39.08324, 39.24047, 39.39751, 
    39.55436, 39.71103, 39.8675, 40.02378, 40.17986, 40.33576, 40.49146, 
    40.64696, 40.80227, 40.95738, 41.1123, 41.26701, 41.42153, 41.57585, 
    41.72997, 41.88388, 42.0376, 42.19111, 42.34442, 42.49753, 42.65043, 
    42.80312, 42.95562, 43.1079, 43.25997, 43.41184, 43.5635, 43.71495, 
    43.86619, 44.01722, 44.16804, 44.31865, 44.46905, 44.61923, 44.7692, 
    44.91896, 45.0685, 45.21783, 45.36694, 45.51584, 45.66452, 45.81299,
  -22.69393, -22.56625, -22.43835, -22.31022, -22.18187, -22.05329, 
    -21.92449, -21.79547, -21.66621, -21.53674, -21.40703, -21.2771, 
    -21.14695, -21.01656, -20.88595, -20.75512, -20.62405, -20.49276, 
    -20.36124, -20.22949, -20.09752, -19.96532, -19.83289, -19.70023, 
    -19.56734, -19.43423, -19.30088, -19.16731, -19.03351, -18.89948, 
    -18.76522, -18.63074, -18.49602, -18.36108, -18.2259, -18.0905, 
    -17.95486, -17.819, -17.68291, -17.54659, -17.41004, -17.27326, 
    -17.13625, -16.99901, -16.86155, -16.72385, -16.58592, -16.44777, 
    -16.30938, -16.17077, -16.03193, -15.89286, -15.75355, -15.61403, 
    -15.47427, -15.33428, -15.19406, -15.05362, -14.91295, -14.77205, 
    -14.63092, -14.48956, -14.34798, -14.20616, -14.06412, -13.92186, 
    -13.77936, -13.63664, -13.49369, -13.35052, -13.20712, -13.06349, 
    -12.91964, -12.77556, -12.63126, -12.48673, -12.34198, -12.197, -12.0518, 
    -11.90637, -11.76072, -11.61485, -11.46875, -11.32243, -11.17589, 
    -11.02913, -10.88215, -10.73494, -10.58752, -10.43987, -10.29201, 
    -10.14392, -9.995617, -9.847094, -9.698352, -9.549393, -9.400216, 
    -9.250823, -9.101213, -8.951388, -8.801348, -8.651093, -8.500623, 
    -8.349938, -8.199042, -8.047933, -7.896611, -7.745078, -7.593334, 
    -7.44138, -7.289217, -7.136844, -6.984262, -6.831473, -6.678476, 
    -6.525274, -6.371865, -6.218251, -6.064433, -5.910411, -5.756186, 
    -5.601759, -5.44713, -5.2923, -5.137271, -4.982042, -4.826614, -4.67099, 
    -4.515167, -4.359149, -4.202936, -4.046528, -3.889927, -3.733133, 
    -3.576147, -3.41897, -3.261603, -3.104046, -2.946302, -2.78837, 
    -2.630252, -2.471948, -2.31346, -2.154788, -1.995934, -1.836898, 
    -1.677681, -1.518285, -1.35871, -1.198958, -1.039029, -0.8789252, 
    -0.7186466, -0.5581948, -0.3975708, -0.2367756, -0.07581042, 0.08532366, 
    0.2466255, 0.408094, 0.569728, 0.7315262, 0.8934876, 1.055611, 1.217895, 
    1.380339, 1.542941, 1.705701, 1.868616, 2.031686, 2.194909, 2.358284, 
    2.521811, 2.685487, 2.849311, 3.013282, 3.177399, 3.341661, 3.506065, 
    3.670611, 3.835298, 4.000124, 4.165086, 4.330186, 4.49542, 4.660788, 
    4.826288, 4.991918, 5.157678, 5.323565, 5.489579, 5.655717, 5.821979, 
    5.988363, 6.154868, 6.321491, 6.488232, 6.655088, 6.82206, 6.989144, 
    7.15634, 7.323646, 7.491059, 7.65858, 7.826206, 7.993936, 8.161767, 
    8.3297, 8.49773, 8.665859, 8.834083, 9.002401, 9.170812, 9.339314, 
    9.507904, 9.676582, 9.845346, 10.0142, 10.18313, 10.35214, 10.52123, 
    10.6904, 10.85964, 11.02896, 11.19835, 11.36782, 11.53735, 11.70695, 
    11.87661, 12.04634, 12.21613, 12.38598, 12.55589, 12.72586, 12.89589, 
    13.06596, 13.23609, 13.40627, 13.5765, 13.74677, 13.91709, 14.08745, 
    14.25785, 14.42829, 14.59877, 14.76929, 14.93984, 15.11042, 15.28103, 
    15.45167, 15.62234, 15.79303, 15.96375, 16.13449, 16.30524, 16.47602, 
    16.64681, 16.81762, 16.98844, 17.15927, 17.33011, 17.50095, 17.6718, 
    17.84266, 18.01351, 18.18437, 18.35522, 18.52607, 18.69692, 18.86776, 
    19.03858, 19.2094, 19.38021, 19.55099, 19.72177, 19.89252, 20.06326, 
    20.23397, 20.40466, 20.57532, 20.74596, 20.91657, 21.08714, 21.25769, 
    21.4282, 21.59867, 21.76911, 21.9395, 22.10986, 22.28017, 22.45044, 
    22.62065, 22.79082, 22.96095, 23.13101, 23.30103, 23.47099, 23.64089, 
    23.81073, 23.98051, 24.15023, 24.31988, 24.48947, 24.65899, 24.82845, 
    24.99783, 25.16713, 25.33637, 25.50552, 25.6746, 25.8436, 26.01252, 
    26.18135, 26.35011, 26.51877, 26.68735, 26.85583, 27.02423, 27.19253, 
    27.36074, 27.52886, 27.69687, 27.86479, 28.0326, 28.20032, 28.36793, 
    28.53543, 28.70283, 28.87012, 29.03729, 29.20436, 29.37131, 29.53815, 
    29.70487, 29.87148, 30.03796, 30.20433, 30.37057, 30.53669, 30.70268, 
    30.86855, 31.03429, 31.1999, 31.36538, 31.53073, 31.69594, 31.86102, 
    32.02596, 32.19076, 32.35543, 32.51995, 32.68433, 32.84857, 33.01266, 
    33.17661, 33.34042, 33.50407, 33.66757, 33.83092, 33.99412, 34.15717, 
    34.32006, 34.48279, 34.64537, 34.80779, 34.97004, 35.13214, 35.29408, 
    35.45585, 35.61746, 35.7789, 35.94018, 36.10128, 36.26222, 36.42299, 
    36.58359, 36.74401, 36.90426, 37.06434, 37.22424, 37.38396, 37.54351, 
    37.70288, 37.86207, 38.02107, 38.1799, 38.33854, 38.497, 38.65528, 
    38.81337, 38.97127, 39.12898, 39.28651, 39.44384, 39.60099, 39.75795, 
    39.91471, 40.07128, 40.22766, 40.38384, 40.53983, 40.69562, 40.85122, 
    41.00661, 41.16181, 41.31681, 41.4716, 41.6262, 41.78059, 41.93479, 
    42.08878, 42.24257, 42.39614, 42.54952, 42.70269, 42.85566, 43.00841, 
    43.16096, 43.3133, 43.46543, 43.61735, 43.76906, 43.92056, 44.07185, 
    44.22293, 44.37379, 44.52444, 44.67487, 44.8251, 44.9751, 45.12489, 
    45.27447, 45.42383, 45.57297, 45.72189, 45.8706,
  -22.76868, -22.64087, -22.51284, -22.38458, -22.2561, -22.12739, -21.99846, 
    -21.86929, -21.7399, -21.61029, -21.48045, -21.35038, -21.22008, 
    -21.08956, -20.9588, -20.82782, -20.69661, -20.56518, -20.43351, 
    -20.30162, -20.16949, -20.03714, -19.90456, -19.77175, -19.63871, 
    -19.50544, -19.37194, -19.23821, -19.10425, -18.97006, -18.83564, 
    -18.70099, -18.56611, -18.43101, -18.29567, -18.1601, -18.02429, 
    -17.88826, -17.752, -17.61551, -17.47879, -17.34183, -17.20465, 
    -17.06724, -16.92959, -16.79172, -16.65361, -16.51527, -16.37671, 
    -16.23791, -16.09888, -15.95962, -15.82014, -15.68042, -15.54047, 
    -15.40029, -15.25988, -15.11924, -14.97838, -14.83728, -14.69595, 
    -14.5544, -14.41261, -14.2706, -14.12836, -13.98589, -13.84319, 
    -13.70026, -13.5571, -13.41372, -13.27011, -13.12627, -12.98221, 
    -12.83791, -12.69339, -12.54865, -12.40368, -12.25848, -12.11306, 
    -11.96741, -11.82154, -11.67544, -11.52912, -11.38257, -11.2358, 
    -11.08881, -10.9416, -10.79416, -10.6465, -10.49862, -10.35052, 
    -10.20219, -10.05365, -9.904884, -9.755901, -9.606699, -9.457277, 
    -9.307638, -9.157781, -9.007707, -8.857416, -8.706909, -8.556187, 
    -8.405249, -8.254096, -8.10273, -7.95115, -7.799358, -7.647353, 
    -7.495137, -7.34271, -7.190072, -7.037224, -6.884167, -6.730902, 
    -6.577429, -6.423749, -6.269862, -6.11577, -5.961472, -5.80697, 
    -5.652265, -5.497356, -5.342246, -5.186934, -5.031422, -4.87571, 
    -4.719799, -4.563689, -4.407382, -4.250879, -4.09418, -3.937286, 
    -3.780198, -3.622916, -3.465443, -3.307778, -3.149923, -2.991878, 
    -2.833645, -2.675224, -2.516616, -2.357822, -2.198844, -2.039681, 
    -1.880336, -1.720809, -1.561101, -1.401214, -1.241148, -1.080903, 
    -0.9204827, -0.7598864, -0.5991156, -0.4381714, -0.2770548, -0.115767, 
    0.0456908, 0.2073176, 0.3691122, 0.5310735, 0.6932002, 0.8554912, 
    1.017945, 1.180562, 1.343338, 1.506275, 1.669369, 1.832621, 1.996028, 
    2.15959, 2.323305, 2.487173, 2.651191, 2.815358, 2.979673, 3.144135, 
    3.308743, 3.473494, 3.638388, 3.803424, 3.9686, 4.133914, 4.299366, 
    4.464953, 4.630675, 4.79653, 4.962516, 5.128633, 5.294878, 5.461251, 
    5.627749, 5.794373, 5.961118, 6.127985, 6.294972, 6.462077, 6.629299, 
    6.796637, 6.964087, 7.131651, 7.299325, 7.467108, 7.634999, 7.802996, 
    7.971097, 8.139301, 8.307607, 8.476012, 8.644515, 8.813114, 8.981809, 
    9.150597, 9.319475, 9.488444, 9.657501, 9.826646, 9.995874, 10.16519, 
    10.33458, 10.50405, 10.6736, 10.84323, 11.01294, 11.18271, 11.35256, 
    11.52248, 11.69246, 11.86251, 12.03263, 12.20281, 12.37305, 12.54334, 
    12.7137, 12.88411, 13.05458, 13.2251, 13.39567, 13.56628, 13.73695, 
    13.90766, 14.07841, 14.2492, 14.42004, 14.59091, 14.76182, 14.93276, 
    15.10374, 15.27474, 15.44578, 15.61684, 15.78793, 15.95904, 16.13017, 
    16.30132, 16.47249, 16.64368, 16.81488, 16.9861, 17.15732, 17.32856, 
    17.4998, 17.67104, 17.84229, 18.01354, 18.1848, 18.35604, 18.52729, 
    18.69853, 18.86976, 19.04099, 19.2122, 19.3834, 19.55458, 19.72575, 
    19.8969, 20.06803, 20.23914, 20.41022, 20.58128, 20.75231, 20.92331, 
    21.09428, 21.26522, 21.43612, 21.60699, 21.77781, 21.9486, 22.11935, 
    22.29005, 22.46071, 22.63132, 22.80188, 22.97239, 23.14285, 23.31325, 
    23.4836, 23.65389, 23.82412, 23.99429, 24.16439, 24.33443, 24.50441, 
    24.67431, 24.84415, 25.01391, 25.18361, 25.35322, 25.52276, 25.69222, 
    25.8616, 26.0309, 26.20012, 26.36925, 26.53829, 26.70724, 26.87611, 
    27.04488, 27.21356, 27.38214, 27.55063, 27.71902, 27.88731, 28.0555, 
    28.22359, 28.39157, 28.55944, 28.72721, 28.89486, 29.06241, 29.22984, 
    29.39716, 29.56436, 29.73145, 29.89842, 30.06527, 30.23199, 30.3986, 
    30.56507, 30.73143, 30.89765, 31.06375, 31.22971, 31.39555, 31.56125, 
    31.72681, 31.89224, 32.05754, 32.22269, 32.3877, 32.55258, 32.7173, 
    32.88189, 33.04633, 33.21062, 33.37476, 33.53876, 33.7026, 33.86629, 
    34.02983, 34.19321, 34.35644, 34.51951, 34.68242, 34.84517, 35.00776, 
    35.17019, 35.33246, 35.49456, 35.65649, 35.81826, 35.97986, 36.14129, 
    36.30255, 36.46364, 36.62456, 36.7853, 36.94587, 37.10626, 37.26648, 
    37.42652, 37.58638, 37.74606, 37.90556, 38.06487, 38.224, 38.38295, 
    38.54172, 38.70029, 38.85869, 39.01689, 39.17491, 39.33273, 39.49036, 
    39.64781, 39.80506, 39.96212, 40.11898, 40.27565, 40.43212, 40.5884, 
    40.74447, 40.90035, 41.05603, 41.21152, 41.36679, 41.52187, 41.67675, 
    41.83142, 41.98589, 42.14016, 42.29422, 42.44807, 42.60172, 42.75516, 
    42.90839, 43.06142, 43.21423, 43.36684, 43.51923, 43.67141, 43.82338, 
    43.97514, 44.12669, 44.27802, 44.42914, 44.58004, 44.73073, 44.8812, 
    45.03146, 45.1815, 45.33132, 45.48093, 45.63031, 45.77948, 45.92843,
  -22.84365, -22.71572, -22.58755, -22.45917, -22.33055, -22.20171, 
    -22.07264, -21.94335, -21.81382, -21.68407, -21.55409, -21.42388, 
    -21.29344, -21.16278, -21.03188, -20.90076, -20.7694, -20.63782, 
    -20.50601, -20.37397, -20.24169, -20.10919, -19.97646, -19.84349, 
    -19.7103, -19.57688, -19.44322, -19.30934, -19.17522, -19.04087, 
    -18.90629, -18.77148, -18.63644, -18.50116, -18.36566, -18.22992, 
    -18.09395, -17.95775, -17.82132, -17.68466, -17.54776, -17.41063, 
    -17.27328, -17.13569, -16.99786, -16.85981, -16.72153, -16.58301, 
    -16.44426, -16.30528, -16.16607, -16.02662, -15.88694, -15.74704, 
    -15.6069, -15.46653, -15.32593, -15.1851, -15.04404, -14.90274, 
    -14.76122, -14.61946, -14.47748, -14.33526, -14.19282, -14.05014, 
    -13.90724, -13.76411, -13.62074, -13.47715, -13.33333, -13.18928, 
    -13.045, -12.90049, -12.75576, -12.6108, -12.46561, -12.32019, -12.17455, 
    -12.02868, -11.88258, -11.73626, -11.58971, -11.44293, -11.29594, 
    -11.14871, -11.00127, -10.8536, -10.7057, -10.55758, -10.40924, 
    -10.26068, -10.1119, -9.962894, -9.813668, -9.664222, -9.514555, 
    -9.364669, -9.214564, -9.06424, -8.913699, -8.76294, -8.611964, 
    -8.460772, -8.309363, -8.15774, -8.005901, -7.853849, -7.701582, 
    -7.549103, -7.396412, -7.243508, -7.090394, -6.937069, -6.783534, 
    -6.62979, -6.475838, -6.321678, -6.16731, -6.012736, -5.857957, 
    -5.702972, -5.547784, -5.392392, -5.236797, -5.081, -4.925003, -4.768805, 
    -4.612407, -4.455811, -4.299016, -4.142025, -3.984838, -3.827455, 
    -3.669878, -3.512107, -3.354143, -3.195988, -3.037642, -2.879106, 
    -2.720381, -2.561468, -2.402368, -2.243082, -2.083611, -1.923955, 
    -1.764117, -1.604097, -1.443895, -1.283514, -1.122953, -0.9622149, 
    -0.8012997, -0.6402088, -0.4789433, -0.3175043, -0.1558928, 0.005889919, 
    0.1678428, 0.3299647, 0.4922543, 0.6547107, 0.8173326, 0.9801187, 
    1.143068, 1.306179, 1.469451, 1.632882, 1.796471, 1.960217, 2.124119, 
    2.288175, 2.452384, 2.616745, 2.781257, 2.945918, 3.110726, 3.275681, 
    3.440781, 3.606025, 3.771411, 3.936939, 4.102605, 4.268411, 4.434353, 
    4.60043, 4.766642, 4.932986, 5.099461, 5.266066, 5.432799, 5.599658, 
    5.766644, 5.933752, 6.100983, 6.268335, 6.435806, 6.603395, 6.7711, 
    6.93892, 7.106852, 7.274896, 7.44305, 7.611313, 7.779682, 7.948157, 
    8.116735, 8.285416, 8.454196, 8.623075, 8.792052, 8.961124, 9.13029, 
    9.299548, 9.468897, 9.638335, 9.807859, 9.97747, 10.14716, 10.31694, 
    10.4868, 10.65673, 10.82675, 10.99684, 11.167, 11.33723, 11.50754, 
    11.67791, 11.84835, 12.01885, 12.18942, 12.36005, 12.53074, 12.70148, 
    12.87229, 13.04314, 13.21405, 13.38501, 13.55602, 13.72708, 13.89818, 
    14.06933, 14.24052, 14.41175, 14.58301, 14.75432, 14.92565, 15.09702, 
    15.26843, 15.43986, 15.61131, 15.7828, 15.95431, 16.12584, 16.29738, 
    16.46895, 16.64054, 16.81213, 16.98375, 17.15537, 17.327, 17.49864, 
    17.67028, 17.84193, 18.01358, 18.18522, 18.35687, 18.52851, 18.70015, 
    18.87178, 19.0434, 19.21501, 19.38661, 19.55819, 19.72975, 19.9013, 
    20.07283, 20.24433, 20.41581, 20.58726, 20.75869, 20.93009, 21.10145, 
    21.27278, 21.44408, 21.61534, 21.78656, 21.95774, 22.12889, 22.29998, 
    22.47103, 22.64203, 22.81298, 22.98389, 23.15474, 23.32553, 23.49627, 
    23.66695, 23.83757, 24.00812, 24.17862, 24.34905, 24.51941, 24.6897, 
    24.85992, 25.03008, 25.20015, 25.37015, 25.54008, 25.70992, 25.87968, 
    26.04937, 26.21896, 26.38847, 26.5579, 26.72723, 26.89647, 27.06563, 
    27.23468, 27.40364, 27.57251, 27.74127, 27.90994, 28.0785, 28.24696, 
    28.41531, 28.58356, 28.75169, 28.91972, 29.08764, 29.25544, 29.42312, 
    29.59069, 29.75814, 29.92548, 30.09269, 30.25978, 30.42674, 30.59358, 
    30.7603, 30.92688, 31.09334, 31.25966, 31.42585, 31.59191, 31.75783, 
    31.92361, 32.08926, 32.25476, 32.42012, 32.58535, 32.75042, 32.91536, 
    33.08014, 33.24478, 33.40926, 33.5736, 33.73779, 33.90182, 34.0657, 
    34.22942, 34.39298, 34.55639, 34.71964, 34.88272, 35.04564, 35.2084, 
    35.371, 35.53343, 35.69569, 35.85779, 36.01971, 36.18147, 36.34305, 
    36.50446, 36.6657, 36.82677, 36.98765, 37.14837, 37.3089, 37.46925, 
    37.62942, 37.78941, 37.94922, 38.10885, 38.26829, 38.42755, 38.58662, 
    38.7455, 38.9042, 39.0627, 39.22102, 39.37914, 39.53708, 39.69482, 
    39.85236, 40.00972, 40.16687, 40.32383, 40.48059, 40.63716, 40.79353, 
    40.94969, 41.10566, 41.26143, 41.41698, 41.57235, 41.7275, 41.88245, 
    42.0372, 42.19174, 42.34608, 42.50021, 42.65413, 42.80783, 42.96134, 
    43.11463, 43.26771, 43.42058, 43.57324, 43.72568, 43.87791, 44.02993, 
    44.18174, 44.33333, 44.4847, 44.63586, 44.7868, 44.93753, 45.08804, 
    45.23832, 45.38839, 45.53825, 45.68788, 45.83729, 45.98648,
  -22.91885, -22.79078, -22.66249, -22.53398, -22.40523, -22.27626, 
    -22.14705, -22.01762, -21.88796, -21.75808, -21.62796, -21.49761, 
    -21.36703, -21.23623, -21.10519, -20.97392, -20.84242, -20.71069, 
    -20.57874, -20.44654, -20.31412, -20.18147, -20.04859, -19.91547, 
    -19.78212, -19.64854, -19.51473, -19.38069, -19.24641, -19.11191, 
    -18.97717, -18.84219, -18.70699, -18.57155, -18.43588, -18.29998, 
    -18.16384, -18.02747, -17.89087, -17.75404, -17.61697, -17.47967, 
    -17.34213, -17.20437, -17.06637, -16.92813, -16.78967, -16.65097, 
    -16.51204, -16.37288, -16.23348, -16.09385, -15.95398, -15.81389, 
    -15.67356, -15.533, -15.39221, -15.25118, -15.10992, -14.96843, 
    -14.82671, -14.68476, -14.54257, -14.40016, -14.25751, -14.11463, 
    -13.97152, -13.82818, -13.68461, -13.54081, -13.39677, -13.25251, 
    -13.10802, -12.9633, -12.81835, -12.67317, -12.52776, -12.38212, 
    -12.23626, -12.09016, -11.94384, -11.7973, -11.65052, -11.50352, 
    -11.35629, -11.20884, -11.06116, -10.91325, -10.76513, -10.61677, 
    -10.46819, -10.31939, -10.17037, -10.02112, -9.871655, -9.721964, 
    -9.572051, -9.421918, -9.271564, -9.120992, -8.970199, -8.819187, 
    -8.667957, -8.51651, -8.364845, -8.212963, -8.060865, -7.908552, 
    -7.756024, -7.603281, -7.450325, -7.297155, -7.143774, -6.99018, 
    -6.836375, -6.682359, -6.528134, -6.373699, -6.219056, -6.064205, 
    -5.909148, -5.753883, -5.598414, -5.442739, -5.286861, -5.130779, 
    -4.974495, -4.818009, -4.661323, -4.504436, -4.34735, -4.190066, 
    -4.032584, -3.874906, -3.717031, -3.558962, -3.400699, -3.242243, 
    -3.083595, -2.924755, -2.765726, -2.606507, -2.447099, -2.287505, 
    -2.127723, -1.967757, -1.807606, -1.647272, -1.486756, -1.326058, 
    -1.16518, -1.004123, -0.8428879, -0.6814759, -0.519888, -0.3581254, 
    -0.1961891, -0.03408032, 0.1281998, 0.2906501, 0.4532694, 0.6160565, 
    0.7790104, 0.9421296, 1.105413, 1.26886, 1.432468, 1.596237, 1.760165, 
    1.924251, 2.088494, 2.252893, 2.417445, 2.582151, 2.747008, 2.912015, 
    3.077171, 3.242475, 3.407925, 3.57352, 3.739258, 3.905138, 4.071159, 
    4.237319, 4.403617, 4.570052, 4.736621, 4.903324, 5.070159, 5.237125, 
    5.40422, 5.571443, 5.738791, 5.906265, 6.073862, 6.24158, 6.409418, 
    6.577375, 6.745449, 6.913639, 7.081942, 7.250358, 7.418885, 7.587521, 
    7.756264, 7.925113, 8.094068, 8.263124, 8.432281, 8.601539, 8.770894, 
    8.940346, 9.109892, 9.279531, 9.449262, 9.619081, 9.788989, 9.958982, 
    10.12906, 10.29922, 10.46947, 10.63979, 10.81019, 10.98066, 11.15121, 
    11.32183, 11.49253, 11.66329, 11.83412, 12.00501, 12.17597, 12.34699, 
    12.51807, 12.68921, 12.86041, 13.03166, 13.20296, 13.37431, 13.54572, 
    13.71717, 13.88867, 14.06021, 14.23179, 14.40342, 14.57508, 14.74678, 
    14.91851, 15.09028, 15.26208, 15.43391, 15.60576, 15.77765, 15.94955, 
    16.12148, 16.29343, 16.46539, 16.63737, 16.80937, 16.98138, 17.1534, 
    17.32543, 17.49747, 17.66951, 17.84156, 18.01361, 18.18566, 18.3577, 
    18.52974, 18.70178, 18.87381, 19.04583, 19.21784, 19.38983, 19.56181, 
    19.73377, 19.90572, 20.07764, 20.24954, 20.42142, 20.59327, 20.7651, 
    20.93689, 21.10865, 21.28038, 21.45208, 21.62373, 21.79535, 21.96693, 
    22.13846, 22.30995, 22.4814, 22.65279, 22.82414, 22.99544, 23.16668, 
    23.33786, 23.509, 23.68007, 23.85108, 24.02202, 24.19291, 24.36373, 
    24.53448, 24.70516, 24.87577, 25.04631, 25.21677, 25.38716, 25.55747, 
    25.7277, 25.89785, 26.06791, 26.23789, 26.40779, 26.57759, 26.74731, 
    26.91693, 27.08647, 27.2559, 27.42524, 27.59448, 27.76362, 27.93266, 
    28.1016, 28.27044, 28.43916, 28.60778, 28.77629, 28.94469, 29.11297, 
    29.28115, 29.4492, 29.61714, 29.78496, 29.95266, 30.12024, 30.28769, 
    30.45502, 30.62222, 30.7893, 30.95624, 31.12305, 31.28974, 31.45628, 
    31.6227, 31.78897, 31.95511, 32.12111, 32.28697, 32.45268, 32.61826, 
    32.78368, 32.94896, 33.1141, 33.27908, 33.44391, 33.60859, 33.77312, 
    33.9375, 34.10172, 34.26578, 34.42968, 34.59342, 34.75701, 34.92043, 
    35.08368, 35.24678, 35.40971, 35.57246, 35.73506, 35.89748, 36.05973, 
    36.22182, 36.38372, 36.54546, 36.70702, 36.8684, 37.02961, 37.19064, 
    37.35149, 37.51216, 37.67265, 37.83295, 37.99307, 38.15301, 38.31276, 
    38.47233, 38.63171, 38.79089, 38.94989, 39.1087, 39.26732, 39.42575, 
    39.58398, 39.74202, 39.89986, 40.05751, 40.21496, 40.37221, 40.52927, 
    40.68612, 40.84278, 40.99923, 41.15548, 41.31153, 41.46738, 41.62302, 
    41.77846, 41.93369, 42.08871, 42.24353, 42.39814, 42.55254, 42.70674, 
    42.86072, 43.01449, 43.16805, 43.3214, 43.47453, 43.62746, 43.78017, 
    43.93266, 44.08494, 44.237, 44.38885, 44.54048, 44.69189, 44.84309, 
    44.99407, 45.14482, 45.29536, 45.44568, 45.59578, 45.74566, 45.89531, 
    46.04475,
  -22.99427, -22.86608, -22.73766, -22.60901, -22.48014, -22.35103, 
    -22.22169, -22.09213, -21.96233, -21.83231, -21.70205, -21.57157, 
    -21.44085, -21.3099, -21.17872, -21.04731, -20.91567, -20.7838, 
    -20.65169, -20.51935, -20.38678, -20.25398, -20.12094, -19.98768, 
    -19.85418, -19.72044, -19.58648, -19.45228, -19.31784, -19.18318, 
    -19.04827, -18.91314, -18.77777, -18.64217, -18.50634, -18.37027, 
    -18.23396, -18.09743, -17.96065, -17.82365, -17.68641, -17.54893, 
    -17.41122, -17.27328, -17.1351, -16.99669, -16.85805, -16.71917, 
    -16.58005, -16.4407, -16.30112, -16.16131, -16.02126, -15.88097, 
    -15.74045, -15.5997, -15.45872, -15.3175, -15.17604, -15.03436, 
    -14.89244, -14.75029, -14.6079, -14.46528, -14.32243, -14.17935, 
    -14.03603, -13.89248, -13.7487, -13.60469, -13.46045, -13.31597, 
    -13.17127, -13.02633, -12.88116, -12.73577, -12.59014, -12.44428, 
    -12.29819, -12.15188, -12.00533, -11.85856, -11.71156, -11.56433, 
    -11.41687, -11.26919, -11.12127, -10.97314, -10.82477, -10.67618, 
    -10.52737, -10.37833, -10.22906, -10.07957, -9.929861, -9.779925, 
    -9.629767, -9.479386, -9.328784, -9.17796, -9.026917, -8.875652, 
    -8.724168, -8.572464, -8.420542, -8.268402, -8.116044, -7.96347, 
    -7.810678, -7.657672, -7.50445, -7.351014, -7.197364, -7.0435, -6.889424, 
    -6.735137, -6.580638, -6.425928, -6.271009, -6.11588, -5.960544, 
    -5.804999, -5.649248, -5.49329, -5.337127, -5.18076, -5.024189, 
    -4.867414, -4.710438, -4.55326, -4.395881, -4.238303, -4.080526, 
    -3.922551, -3.764379, -3.606011, -3.447447, -3.288689, -3.129738, 
    -2.970594, -2.811259, -2.651733, -2.492017, -2.332113, -2.172021, 
    -2.011742, -1.851278, -1.690629, -1.529797, -1.368782, -1.207585, 
    -1.046209, -0.8846524, -0.7229182, -0.5610068, -0.3989194, -0.2366572, 
    -0.07422127, 0.08838721, 0.2511671, 0.4141172, 0.5772363, 0.7405233, 
    0.9039769, 1.067596, 1.231379, 1.395325, 1.559433, 1.723702, 1.888129, 
    2.052714, 2.217456, 2.382354, 2.547405, 2.712609, 2.877964, 3.043469, 
    3.209123, 3.374924, 3.540871, 3.706963, 3.873198, 4.039574, 4.20609, 
    4.372746, 4.539539, 4.706468, 4.873531, 5.040728, 5.208056, 5.375514, 
    5.543101, 5.710815, 5.878654, 6.046618, 6.214705, 6.382912, 6.551239, 
    6.719683, 6.888244, 7.05692, 7.225709, 7.39461, 7.563621, 7.732739, 
    7.901966, 8.071297, 8.240731, 8.410268, 8.579906, 8.74964, 8.919474, 
    9.089401, 9.259422, 9.429536, 9.59974, 9.770032, 9.940412, 10.11088, 
    10.28142, 10.45205, 10.62276, 10.79355, 10.96441, 11.13535, 11.30637, 
    11.47745, 11.6486, 11.81982, 11.99111, 12.16246, 12.33387, 12.50535, 
    12.67688, 12.84847, 13.02012, 13.19182, 13.36357, 13.53537, 13.70721, 
    13.87911, 14.05105, 14.22303, 14.39505, 14.56711, 14.73921, 14.91134, 
    15.08351, 15.2557, 15.42793, 15.60019, 15.77247, 15.94477, 16.1171, 
    16.28945, 16.46182, 16.6342, 16.8066, 16.97901, 17.15143, 17.32386, 
    17.4963, 17.66874, 17.84119, 18.01364, 18.18609, 18.35854, 18.53098, 
    18.70341, 18.87584, 19.04827, 19.22067, 19.39307, 19.56545, 19.73781, 
    19.91016, 20.08248, 20.25479, 20.42706, 20.59931, 20.77154, 20.94373, 
    21.11589, 21.28802, 21.46011, 21.63216, 21.80418, 21.97615, 22.14809, 
    22.31997, 22.49181, 22.66361, 22.83535, 23.00704, 23.17867, 23.35026, 
    23.52178, 23.69324, 23.86465, 24.03599, 24.20727, 24.37848, 24.54962, 
    24.72069, 24.89169, 25.06262, 25.23347, 25.40425, 25.57494, 25.74556, 
    25.91609, 26.08655, 26.25691, 26.42719, 26.59738, 26.76748, 26.93748, 
    27.1074, 27.27722, 27.44694, 27.61656, 27.78608, 27.9555, 28.12481, 
    28.29402, 28.46312, 28.63211, 28.801, 28.96977, 29.13843, 29.30697, 
    29.4754, 29.6437, 29.81189, 29.97996, 30.1479, 30.31572, 30.48342, 
    30.65098, 30.81842, 30.98573, 31.1529, 31.31995, 31.48685, 31.65363, 
    31.82026, 31.98675, 32.15311, 32.31932, 32.48539, 32.65131, 32.81709, 
    32.98272, 33.1482, 33.31353, 33.47871, 33.64374, 33.80861, 33.97333, 
    34.13789, 34.30229, 34.46654, 34.63062, 34.79454, 34.9583, 35.12189, 
    35.28532, 35.44858, 35.61167, 35.77459, 35.93735, 36.09993, 36.26234, 
    36.42457, 36.58663, 36.74851, 36.91022, 37.07175, 37.2331, 37.39426, 
    37.55525, 37.71605, 37.87667, 38.03711, 38.19736, 38.35742, 38.5173, 
    38.67698, 38.83648, 38.99578, 39.1549, 39.31382, 39.47254, 39.63108, 
    39.78941, 39.94755, 40.1055, 40.26324, 40.42079, 40.57814, 40.73528, 
    40.89223, 41.04897, 41.20551, 41.36184, 41.51797, 41.6739, 41.82962, 
    41.98513, 42.14043, 42.29553, 42.45042, 42.60509, 42.75956, 42.91381, 
    43.06785, 43.22168, 43.3753, 43.5287, 43.68189, 43.83486, 43.98762, 
    44.14016, 44.29248, 44.44459, 44.59648, 44.74815, 44.89959, 45.05082, 
    45.20183, 45.35262, 45.50319, 45.65353, 45.80366, 45.95356, 46.10324,
  -23.06992, -22.9416, -22.81306, -22.68428, -22.55527, -22.42603, -22.29656, 
    -22.16686, -22.03693, -21.90677, -21.77638, -21.64576, -21.5149, 
    -21.38381, -21.25249, -21.12094, -20.98915, -20.85713, -20.72488, 
    -20.59239, -20.45967, -20.32672, -20.19353, -20.06012, -19.92646, 
    -19.79257, -19.65845, -19.52409, -19.3895, -19.25468, -19.11962, 
    -18.98432, -18.84879, -18.71302, -18.57702, -18.44079, -18.30432, 
    -18.16761, -18.03067, -17.89349, -17.75608, -17.61843, -17.48055, 
    -17.34243, -17.20407, -17.06548, -16.92666, -16.7876, -16.6483, 
    -16.50877, -16.369, -16.229, -16.08876, -15.94829, -15.80758, -15.66663, 
    -15.52546, -15.38404, -15.2424, -15.10051, -14.9584, -14.81604, 
    -14.67346, -14.53064, -14.38758, -14.24429, -14.10077, -13.95702, 
    -13.81303, -13.66881, -13.52435, -13.37967, -13.23475, -13.08959, 
    -12.94421, -12.7986, -12.65275, -12.50667, -12.36036, -12.21382, 
    -12.06705, -11.92005, -11.77282, -11.62537, -11.47768, -11.32976, 
    -11.18162, -11.03325, -10.88465, -10.73582, -10.58676, -10.43748, 
    -10.28798, -10.13825, -9.988291, -9.83811, -9.687705, -9.537076, 
    -9.386225, -9.23515, -9.083854, -8.932336, -8.780596, -8.628636, 
    -8.476457, -8.324058, -8.171439, -8.018602, -7.865548, -7.712277, 
    -7.558789, -7.405086, -7.251167, -7.097033, -6.942686, -6.788125, 
    -6.633352, -6.478366, -6.32317, -6.167763, -6.012147, -5.856321, 
    -5.700287, -5.544046, -5.387598, -5.230944, -5.074084, -4.917021, 
    -4.759753, -4.602283, -4.444612, -4.286739, -4.128666, -3.970393, 
    -3.811923, -3.653254, -3.494389, -3.335329, -3.176073, -3.016624, 
    -2.856982, -2.697148, -2.537123, -2.376908, -2.216504, -2.055912, 
    -1.895134, -1.734169, -1.57302, -1.411686, -1.25017, -1.088473, 
    -0.9265946, -0.764537, -0.602301, -0.4398878, -0.2772985, -0.1145343, 
    0.04840375, 0.2115144, 0.3747965, 0.5382487, 0.7018701, 0.8656593, 
    1.029615, 1.193736, 1.358021, 1.52247, 1.687079, 1.851849, 2.016778, 
    2.181865, 2.347109, 2.512507, 2.678059, 2.843764, 3.009619, 3.175625, 
    3.341779, 3.508079, 3.674525, 3.841116, 4.007849, 4.174724, 4.341738, 
    4.508891, 4.67618, 4.843606, 5.011165, 5.178857, 5.34668, 5.514633, 
    5.682714, 5.850921, 6.019253, 6.187709, 6.356287, 6.524984, 6.693801, 
    6.862735, 7.031785, 7.200949, 7.370225, 7.539613, 7.709109, 7.878713, 
    8.048423, 8.218238, 8.388155, 8.558173, 8.728291, 8.898505, 9.068817, 
    9.239223, 9.40972, 9.58031, 9.750989, 9.921755, 10.09261, 10.26354, 
    10.43456, 10.60566, 10.77684, 10.94809, 11.11942, 11.29083, 11.4623, 
    11.63385, 11.80546, 11.97714, 12.14889, 12.3207, 12.49257, 12.66449, 
    12.83648, 13.00852, 13.18062, 13.35277, 13.52496, 13.69721, 13.8695, 
    14.04184, 14.21422, 14.38664, 14.5591, 14.7316, 14.90413, 15.0767, 
    15.2493, 15.42193, 15.59459, 15.76727, 15.93998, 16.11271, 16.28546, 
    16.45822, 16.63101, 16.80381, 16.97662, 17.14945, 17.32228, 17.49512, 
    17.66797, 17.84082, 18.01367, 18.18652, 18.35937, 18.53222, 18.70506, 
    18.87789, 19.05071, 19.22353, 19.39632, 19.56911, 19.74187, 19.91462, 
    20.08735, 20.26005, 20.43273, 20.60538, 20.778, 20.9506, 21.12316, 
    21.29569, 21.46818, 21.64063, 21.81305, 21.98542, 22.15775, 22.33004, 
    22.50228, 22.67447, 22.84661, 23.0187, 23.19073, 23.36271, 23.53462, 
    23.70648, 23.87828, 24.05002, 24.22169, 24.39329, 24.56483, 24.73629, 
    24.90768, 25.079, 25.25024, 25.42141, 25.5925, 25.7635, 25.93443, 
    26.10526, 26.27602, 26.44668, 26.61726, 26.78774, 26.95813, 27.12843, 
    27.29863, 27.46873, 27.63873, 27.80863, 27.97843, 28.14812, 28.31771, 
    28.48719, 28.65656, 28.82582, 28.99496, 29.164, 29.33291, 29.50171, 
    29.67039, 29.83895, 30.00738, 30.1757, 30.34388, 30.51194, 30.67988, 
    30.84768, 31.01535, 31.18289, 31.35029, 31.51756, 31.68469, 31.85168, 
    32.01854, 32.18525, 32.35181, 32.51824, 32.68451, 32.85064, 33.01662, 
    33.18246, 33.34814, 33.51367, 33.67904, 33.84426, 34.00932, 34.17422, 
    34.33897, 34.50356, 34.66798, 34.83224, 34.99633, 35.16026, 35.32402, 
    35.48762, 35.65104, 35.8143, 35.97738, 36.14029, 36.30303, 36.46559, 
    36.62798, 36.79018, 36.95221, 37.11406, 37.27573, 37.43722, 37.59852, 
    37.75964, 37.92058, 38.08133, 38.24189, 38.40226, 38.56245, 38.72244, 
    38.88225, 39.04186, 39.20128, 39.3605, 39.51953, 39.67837, 39.837, 
    39.99544, 40.15368, 40.31173, 40.46957, 40.6272, 40.78465, 40.94188, 
    41.09891, 41.25574, 41.41236, 41.56878, 41.72498, 41.88099, 42.03678, 
    42.19236, 42.34773, 42.5029, 42.65785, 42.81259, 42.96711, 43.12143, 
    43.27553, 43.42941, 43.58308, 43.73654, 43.88977, 44.04279, 44.19559, 
    44.34818, 44.50054, 44.65269, 44.80462, 44.95632, 45.1078, 45.25906, 
    45.4101, 45.56092, 45.71151, 45.86188, 46.01203, 46.16195,
  -23.1458, -23.01735, -22.88868, -22.75977, -22.63063, -22.50126, -22.37166, 
    -22.24183, -22.11176, -21.98147, -21.85094, -21.72017, -21.58918, 
    -21.45795, -21.32649, -21.19479, -21.06286, -20.9307, -20.7983, 
    -20.66566, -20.5328, -20.3997, -20.26636, -20.13279, -19.99898, 
    -19.86494, -19.73066, -19.59615, -19.4614, -19.32641, -19.19119, 
    -19.05573, -18.92004, -18.78411, -18.64795, -18.51154, -18.3749, 
    -18.23803, -18.10092, -17.96357, -17.82598, -17.68816, -17.5501, 
    -17.41181, -17.27328, -17.13451, -16.9955, -16.85626, -16.71678, 
    -16.57707, -16.43711, -16.29692, -16.1565, -16.01584, -15.87494, 
    -15.7338, -15.59243, -15.45082, -15.30898, -15.1669, -15.02459, 
    -14.88203, -14.73925, -14.59623, -14.45297, -14.30947, -14.16575, 
    -14.02178, -13.87759, -13.73316, -13.58849, -13.44359, -13.29846, 
    -13.15309, -13.00749, -12.86166, -12.71559, -12.56929, -12.42276, 
    -12.276, -12.129, -11.98178, -11.83432, -11.68663, -11.53871, -11.39056, 
    -11.24219, -11.09358, -10.94474, -10.79568, -10.64639, -10.49687, 
    -10.34712, -10.19715, -10.04694, -9.896518, -9.745866, -9.594989, 
    -9.443887, -9.292561, -9.141012, -8.98924, -8.837245, -8.685028, 
    -8.53259, -8.37993, -8.227052, -8.073953, -7.920635, -7.767098, 
    -7.613344, -7.459372, -7.305183, -7.150779, -6.99616, -6.841325, 
    -6.686277, -6.531015, -6.375542, -6.219855, -6.063958, -5.907851, 
    -5.751534, -5.595007, -5.438273, -5.281332, -5.124184, -4.96683, 
    -4.809271, -4.651509, -4.493543, -4.335374, -4.177004, -4.018434, 
    -3.859663, -3.700694, -3.541527, -3.382162, -3.222602, -3.062846, 
    -2.902897, -2.742754, -2.582418, -2.421892, -2.261175, -2.100269, 
    -1.939175, -1.777894, -1.616426, -1.454773, -1.292937, -1.130917, 
    -0.9687158, -0.8063338, -0.6437721, -0.4810319, -0.3181144, -0.1550207, 
    0.008248037, 0.1716906, 0.3353058, 0.4990925, 0.6630494, 0.8271754, 
    0.9914691, 1.155929, 1.320555, 1.485345, 1.650297, 1.815411, 1.980685, 
    2.146118, 2.311709, 2.477456, 2.643357, 2.809412, 2.97562, 3.141978, 
    3.308486, 3.475142, 3.641944, 3.808892, 3.975983, 4.143217, 4.310591, 
    4.478106, 4.645758, 4.813546, 4.98147, 5.149527, 5.317717, 5.486036, 
    5.654485, 5.823062, 5.991764, 6.160591, 6.329541, 6.498612, 6.667802, 
    6.837111, 7.006536, 7.176077, 7.34573, 7.515496, 7.685371, 7.855355, 
    8.025445, 8.195642, 8.36594, 8.536342, 8.706842, 8.877442, 9.048139, 
    9.21893, 9.389815, 9.560791, 9.731858, 9.903012, 10.07425, 10.24558, 
    10.41699, 10.58848, 10.76005, 10.9317, 11.10342, 11.27522, 11.44709, 
    11.61903, 11.79104, 11.96311, 12.13525, 12.30746, 12.47972, 12.65205, 
    12.82444, 12.99688, 13.16937, 13.34192, 13.51451, 13.68716, 13.85985, 
    14.03259, 14.20537, 14.3782, 14.55106, 14.72396, 14.8969, 15.06986, 
    15.24287, 15.4159, 15.58896, 15.76204, 15.93515, 16.10829, 16.28144, 
    16.45461, 16.6278, 16.80101, 16.97423, 17.14746, 17.32069, 17.49394, 
    17.66719, 17.84045, 18.0137, 18.18696, 18.36021, 18.53346, 18.70671, 
    18.87995, 19.05317, 19.22639, 19.39959, 19.57278, 19.74595, 19.9191, 
    20.09223, 20.26534, 20.43842, 20.61147, 20.7845, 20.9575, 21.13046, 
    21.30339, 21.47629, 21.64914, 21.82196, 21.99473, 22.16747, 22.34015, 
    22.51279, 22.68538, 22.85792, 23.03041, 23.20284, 23.37521, 23.54753, 
    23.71979, 23.89198, 24.06411, 24.23618, 24.40818, 24.5801, 24.75196, 
    24.92375, 25.09546, 25.2671, 25.43865, 25.61013, 25.78153, 25.95284, 
    26.12407, 26.29521, 26.46626, 26.63722, 26.80809, 26.97887, 27.14955, 
    27.32014, 27.49062, 27.66101, 27.83129, 28.00147, 28.17154, 28.34151, 
    28.51137, 28.68111, 28.85075, 29.02027, 29.18968, 29.35897, 29.52814, 
    29.69719, 29.86612, 30.03493, 30.20361, 30.37217, 30.5406, 30.7089, 
    30.87707, 31.0451, 31.21301, 31.38077, 31.5484, 31.71589, 31.88325, 
    32.05046, 32.21753, 32.38445, 32.55123, 32.71786, 32.88435, 33.05068, 
    33.21687, 33.3829, 33.54877, 33.7145, 33.88006, 34.04547, 34.21072, 
    34.3758, 34.54073, 34.7055, 34.8701, 35.03453, 35.1988, 35.3629, 
    35.52683, 35.69059, 35.85418, 36.01759, 36.18083, 36.3439, 36.50679, 
    36.6695, 36.83203, 36.99438, 37.15656, 37.31855, 37.48036, 37.64198, 
    37.80342, 37.96467, 38.12574, 38.28661, 38.4473, 38.60779, 38.7681, 
    38.92821, 39.08813, 39.24786, 39.40738, 39.56672, 39.72585, 39.88479, 
    40.04353, 40.20207, 40.36041, 40.51854, 40.67648, 40.83421, 40.99173, 
    41.14906, 41.30617, 41.46308, 41.61978, 41.77628, 41.93256, 42.08863, 
    42.2445, 42.40015, 42.55559, 42.71082, 42.86583, 43.02063, 43.17522, 
    43.32959, 43.48374, 43.63768, 43.7914, 43.9449, 44.09819, 44.25125, 
    44.40409, 44.55672, 44.70912, 44.8613, 45.01326, 45.165, 45.31651, 
    45.4678, 45.61887, 45.76971, 45.92033, 46.07072, 46.22088,
  -23.22191, -23.09334, -22.96453, -22.8355, -22.70623, -22.57673, -22.44699, 
    -22.31703, -22.18683, -22.05639, -21.92573, -21.79482, -21.66369, 
    -21.53232, -21.40072, -21.26888, -21.1368, -21.0045, -20.87195, 
    -20.73917, -20.60616, -20.4729, -20.33942, -20.20569, -20.07173, 
    -19.93754, -19.8031, -19.66843, -19.53353, -19.39838, -19.263, -19.12738, 
    -18.99153, -18.85543, -18.7191, -18.58253, -18.44573, -18.30869, 
    -18.1714, -18.03388, -17.89613, -17.75813, -17.6199, -17.48143, 
    -17.34272, -17.20377, -17.06458, -16.92516, -16.7855, -16.6456, 
    -16.50546, -16.36509, -16.22447, -16.08362, -15.94253, -15.80121, 
    -15.65964, -15.51784, -15.3758, -15.23353, -15.09101, -14.94826, 
    -14.80527, -14.66205, -14.51859, -14.37489, -14.23096, -14.08679, 
    -13.94238, -13.79774, -13.65286, -13.50775, -13.3624, -13.21682, -13.071, 
    -12.92495, -12.77866, -12.63214, -12.48539, -12.3384, -12.19118, 
    -12.04373, -11.89604, -11.74813, -11.59998, -11.4516, -11.30299, 
    -11.15414, -11.00507, -10.85577, -10.70624, -10.55648, -10.40649, 
    -10.25627, -10.10582, -9.955151, -9.804251, -9.653125, -9.501773, 
    -9.350195, -9.198393, -9.046366, -8.894115, -8.741641, -8.588943, 
    -8.436025, -8.282884, -8.129521, -7.975939, -7.822137, -7.668115, 
    -7.513875, -7.359416, -7.204741, -7.049848, -6.89474, -6.739416, 
    -6.583877, -6.428124, -6.272159, -6.11598, -5.95959, -5.802989, 
    -5.646177, -5.489156, -5.331926, -5.174489, -5.016844, -4.858993, 
    -4.700937, -4.542675, -4.384211, -4.225543, -4.066673, -3.907602, 
    -3.748331, -3.588861, -3.429192, -3.269325, -3.109263, -2.949004, 
    -2.788552, -2.627905, -2.467066, -2.306035, -2.144814, -1.983403, 
    -1.821804, -1.660017, -1.498044, -1.335886, -1.173543, -1.011018, 
    -0.8483099, -0.6854214, -0.5223531, -0.3591062, -0.1956819, -0.03208131, 
    0.1316944, 0.2956439, 0.4597662, 0.6240599, 0.7885239, 0.9531568, 
    1.117958, 1.282925, 1.448057, 1.613354, 1.778813, 1.944433, 2.110214, 
    2.276153, 2.44225, 2.608502, 2.774909, 2.94147, 3.108182, 3.275045, 
    3.442058, 3.609217, 3.776524, 3.943974, 4.111569, 4.279305, 4.447182, 
    4.615198, 4.783352, 4.951642, 5.120066, 5.288623, 5.457312, 5.62613, 
    5.795077, 5.964151, 6.133351, 6.302674, 6.472119, 6.641685, 6.81137, 
    6.981173, 7.151091, 7.321124, 7.491269, 7.661525, 7.83189, 8.002362, 
    8.172941, 8.343624, 8.51441, 8.685296, 8.856282, 9.027366, 9.198545, 
    9.369818, 9.541183, 9.712639, 9.884184, 10.05582, 10.22753, 10.39933, 
    10.57122, 10.74318, 10.91522, 11.08734, 11.25953, 11.4318, 11.60414, 
    11.77654, 11.94902, 12.12156, 12.29416, 12.46682, 12.63955, 12.81233, 
    12.98517, 13.15807, 13.33102, 13.50402, 13.67706, 13.85016, 14.0233, 
    14.19649, 14.36971, 14.54298, 14.71628, 14.88962, 15.06299, 15.2364, 
    15.40984, 15.5833, 15.75679, 15.93031, 16.10385, 16.27741, 16.45099, 
    16.62458, 16.79819, 16.97182, 17.14545, 17.3191, 17.49275, 17.66641, 
    17.84007, 18.01373, 18.1874, 18.36106, 18.53472, 18.70837, 18.88201, 
    19.05565, 19.22927, 19.40288, 19.57647, 19.75005, 19.9236, 20.09714, 
    20.27065, 20.44414, 20.6176, 20.79103, 20.96443, 21.1378, 21.31113, 
    21.48443, 21.65769, 21.83091, 22.00409, 22.17722, 22.35031, 22.52335, 
    22.69634, 22.86928, 23.04217, 23.215, 23.38778, 23.56049, 23.73315, 
    23.90574, 24.07827, 24.25073, 24.42313, 24.59546, 24.76771, 24.93989, 
    25.112, 25.28403, 25.45598, 25.62785, 25.79963, 25.97134, 26.14296, 
    26.31449, 26.48593, 26.65728, 26.82854, 26.9997, 27.17077, 27.34174, 
    27.51261, 27.68338, 27.85405, 28.02461, 28.19507, 28.36541, 28.53565, 
    28.70578, 28.8758, 29.04569, 29.21548, 29.38515, 29.55469, 29.72412, 
    29.89342, 30.0626, 30.23166, 30.40058, 30.56938, 30.73805, 30.90659, 
    31.07499, 31.24326, 31.41139, 31.57938, 31.74724, 31.91495, 32.08252, 
    32.24995, 32.41723, 32.58437, 32.75136, 32.9182, 33.08489, 33.25142, 
    33.41781, 33.58403, 33.75011, 33.91602, 34.08178, 34.24737, 34.4128, 
    34.57808, 34.74318, 34.90812, 35.0729, 35.2375, 35.40194, 35.56621, 
    35.7303, 35.89422, 36.05797, 36.22155, 36.38494, 36.54816, 36.7112, 
    36.87406, 37.03674, 37.19923, 37.36155, 37.52368, 37.68562, 37.84738, 
    38.00895, 38.17033, 38.33152, 38.49252, 38.65333, 38.81395, 38.97437, 
    39.13459, 39.29463, 39.45446, 39.6141, 39.77354, 39.93278, 40.09182, 
    40.25066, 40.40929, 40.56772, 40.72595, 40.88398, 41.04179, 41.19941, 
    41.35681, 41.51401, 41.671, 41.82777, 41.98434, 42.1407, 42.29684, 
    42.45278, 42.60849, 42.764, 42.91929, 43.07436, 43.22922, 43.38387, 
    43.53829, 43.69249, 43.84648, 44.00025, 44.1538, 44.30712, 44.46023, 
    44.61311, 44.76577, 44.91821, 45.07043, 45.22242, 45.37419, 45.52573, 
    45.67704, 45.82814, 45.979, 46.12964, 46.28004,
  -23.29825, -23.16955, -23.04062, -22.91145, -22.78205, -22.65242, 
    -22.52256, -22.39246, -22.26212, -22.13155, -22.00075, -21.86971, 
    -21.73844, -21.60693, -21.47518, -21.3432, -21.21098, -21.07853, 
    -20.94584, -20.81291, -20.67975, -20.54635, -20.41271, -20.27884, 
    -20.14472, -20.01037, -19.87578, -19.74096, -19.60589, -19.47059, 
    -19.33505, -19.19927, -19.06325, -18.927, -18.7905, -18.65376, -18.51679, 
    -18.37958, -18.24213, -18.10444, -17.96651, -17.82834, -17.68993, 
    -17.55128, -17.4124, -17.27327, -17.1339, -16.9943, -16.85446, -16.71437, 
    -16.57405, -16.43349, -16.29269, -16.15165, -16.01037, -15.86885, 
    -15.72709, -15.5851, -15.44286, -15.30039, -15.15768, -15.01472, 
    -14.87154, -14.72811, -14.58444, -14.44054, -14.2964, -14.15202, 
    -14.00741, -13.86256, -13.71747, -13.57214, -13.42658, -13.28078, 
    -13.13474, -12.98847, -12.84197, -12.69523, -12.54825, -12.40104, 
    -12.25359, -12.10591, -11.958, -11.80985, -11.66147, -11.51286, 
    -11.36401, -11.21494, -11.06563, -10.91609, -10.76632, -10.61631, 
    -10.46608, -10.31562, -10.16493, -10.01401, -9.862863, -9.711487, 
    -9.559884, -9.408054, -9.255998, -9.103716, -8.951208, -8.798476, 
    -8.64552, -8.49234, -8.338937, -8.185311, -8.031464, -7.877395, 
    -7.723105, -7.568595, -7.413867, -7.258918, -7.103752, -6.948369, 
    -6.792768, -6.636952, -6.48092, -6.324674, -6.168213, -6.01154, 
    -5.854654, -5.697556, -5.540248, -5.382729, -5.225001, -5.067065, 
    -4.90892, -4.750569, -4.592012, -4.43325, -4.274284, -4.115114, 
    -3.955742, -3.796168, -3.636393, -3.476419, -3.316246, -3.155874, 
    -2.995307, -2.834543, -2.673584, -2.512431, -2.351086, -2.189548, 
    -2.02782, -1.865902, -1.703795, -1.5415, -1.379019, -1.216352, -1.053501, 
    -0.8904669, -0.7272504, -0.5638528, -0.4002754, -0.2365193, -0.07258566, 
    0.09152431, 0.2558094, 0.4202685, 0.5849002, 0.7497034, 0.9146769, 
    1.079819, 1.245129, 1.410606, 1.576248, 1.742053, 1.908021, 2.074151, 
    2.24044, 2.406888, 2.573492, 2.740253, 2.907168, 3.074236, 3.241456, 
    3.408826, 3.576345, 3.744011, 3.911823, 4.07978, 4.247879, 4.416121, 
    4.584502, 4.753022, 4.921679, 5.090471, 5.259398, 5.428456, 5.597647, 
    5.766966, 5.936413, 6.105987, 6.275685, 6.445507, 6.615449, 6.785512, 
    6.955694, 7.125991, 7.296404, 7.466931, 7.637569, 7.808317, 7.979174, 
    8.150137, 8.321205, 8.492377, 8.663651, 8.835025, 9.006496, 9.178064, 
    9.349728, 9.521483, 9.693331, 9.865269, 10.03729, 10.2094, 10.3816, 
    10.55388, 10.72624, 10.89867, 11.07119, 11.24378, 11.41644, 11.58918, 
    11.76198, 11.93485, 12.10779, 12.2808, 12.45386, 12.62699, 12.80018, 
    12.97342, 13.14672, 13.32007, 13.49347, 13.66692, 13.84042, 14.01397, 
    14.18756, 14.36119, 14.53486, 14.70857, 14.88231, 15.05609, 15.22991, 
    15.40375, 15.57762, 15.75152, 15.92544, 16.09939, 16.27336, 16.44735, 
    16.62135, 16.79537, 16.9694, 17.14344, 17.3175, 17.49156, 17.66562, 
    17.83969, 18.01377, 18.18784, 18.36191, 18.53597, 18.71004, 18.88409, 
    19.05813, 19.23216, 19.40618, 19.58018, 19.75416, 19.92813, 20.10207, 
    20.27599, 20.44988, 20.62375, 20.79759, 20.9714, 21.14517, 21.31891, 
    21.49262, 21.66628, 21.83991, 22.01349, 22.18703, 22.36052, 22.53396, 
    22.70736, 22.8807, 23.05399, 23.22722, 23.4004, 23.57352, 23.74657, 
    23.91957, 24.0925, 24.26536, 24.43815, 24.61088, 24.78353, 24.95611, 
    25.12861, 25.30103, 25.47338, 25.64565, 25.81783, 25.98992, 26.16194, 
    26.33386, 26.50569, 26.67743, 26.84908, 27.02063, 27.19209, 27.36345, 
    27.53471, 27.70586, 27.87691, 28.04786, 28.2187, 28.38943, 28.56005, 
    28.73056, 28.90096, 29.07123, 29.2414, 29.41144, 29.58136, 29.75117, 
    29.92085, 30.0904, 30.25983, 30.42912, 30.5983, 30.76733, 30.93624, 
    31.10501, 31.27365, 31.44214, 31.6105, 31.77872, 31.9468, 32.11473, 
    32.28252, 32.45016, 32.61766, 32.78501, 32.9522, 33.11925, 33.28614, 
    33.45287, 33.61945, 33.78587, 33.95214, 34.11824, 34.28418, 34.44997, 
    34.61558, 34.78103, 34.94632, 35.11143, 35.27638, 35.44115, 35.60576, 
    35.77019, 35.93445, 36.09853, 36.26244, 36.42616, 36.58971, 36.75308, 
    36.91627, 37.07927, 37.2421, 37.40473, 37.56718, 37.72945, 37.89153, 
    38.05342, 38.21511, 38.37662, 38.53794, 38.69906, 38.85999, 39.02072, 
    39.18126, 39.34159, 39.50174, 39.66168, 39.82142, 39.98096, 40.1403, 
    40.29944, 40.45838, 40.61711, 40.77563, 40.93395, 41.09206, 41.24997, 
    41.40766, 41.56514, 41.72242, 41.87949, 42.03634, 42.19298, 42.3494, 
    42.50562, 42.66161, 42.8174, 42.97296, 43.12831, 43.28344, 43.43836, 
    43.59305, 43.74752, 43.90178, 44.05581, 44.20963, 44.36322, 44.51659, 
    44.66973, 44.82265, 44.97535, 45.12782, 45.28007, 45.43209, 45.58388, 
    45.73545, 45.88679, 46.0379, 46.18878, 46.33944,
  -23.37482, -23.246, -23.11694, -22.98764, -22.85812, -22.72835, -22.59835, 
    -22.46812, -22.33765, -22.20695, -22.07601, -21.94483, -21.81342, 
    -21.68177, -21.54988, -21.41776, -21.2854, -21.1528, -21.01997, 
    -20.88689, -20.75358, -20.62003, -20.48624, -20.35222, -20.21795, 
    -20.08345, -19.9487, -19.81372, -19.6785, -19.54304, -19.40734, -19.2714, 
    -19.13522, -18.99879, -18.86213, -18.72523, -18.58809, -18.45071, 
    -18.31309, -18.17523, -18.03713, -17.89878, -17.7602, -17.62138, 
    -17.48231, -17.34301, -17.20346, -17.06368, -16.92365, -16.78338, 
    -16.64288, -16.50213, -16.36114, -16.21991, -16.07844, -15.93673, 
    -15.79478, -15.65259, -15.51016, -15.36749, -15.22458, -15.08143, 
    -14.93804, -14.79441, -14.65054, -14.50643, -14.36208, -14.2175, 
    -14.07267, -13.92761, -13.78231, -13.63677, -13.49099, -13.34498, 
    -13.19873, -13.05224, -12.90551, -12.75855, -12.61135, -12.46391, 
    -12.31624, -12.16833, -12.02019, -11.87181, -11.7232, -11.57436, 
    -11.42528, -11.27596, -11.12642, -10.97664, -10.82663, -10.67638, 
    -10.52591, -10.3752, -10.22427, -10.0731, -9.921702, -9.770077, 
    -9.618222, -9.46614, -9.313829, -9.161291, -9.008527, -8.855536, 
    -8.70232, -8.548879, -8.395212, -8.241323, -8.08721, -7.932873, 
    -7.778316, -7.623536, -7.468535, -7.313314, -7.157874, -7.002215, 
    -6.846338, -6.690243, -6.533931, -6.377403, -6.22066, -6.063703, 
    -5.906531, -5.749146, -5.591549, -5.433741, -5.275722, -5.117493, 
    -4.959054, -4.800408, -4.641554, -4.482494, -4.323228, -4.163757, 
    -4.004083, -3.844205, -3.684125, -3.523844, -3.363364, -3.202683, 
    -3.041805, -2.880729, -2.719457, -2.55799, -2.396328, -2.234473, 
    -2.072427, -1.910188, -1.74776, -1.585143, -1.422338, -1.259346, 
    -1.096168, -0.9328061, -0.7692605, -0.6055325, -0.4416234, -0.2775343, 
    -0.1132664, 0.05117904, 0.2158009, 0.380598, 0.5455689, 0.7107127, 
    0.8760279, 1.041513, 1.207168, 1.372989, 1.538978, 1.705131, 1.871448, 
    2.037927, 2.204568, 2.371368, 2.538327, 2.705442, 2.872713, 3.040138, 
    3.207716, 3.375445, 3.543324, 3.711352, 3.879527, 4.047847, 4.216311, 
    4.384918, 4.553666, 4.722554, 4.89158, 5.060742, 5.23004, 5.39947, 
    5.569033, 5.738727, 5.908549, 6.078498, 6.248573, 6.418772, 6.589094, 
    6.759536, 6.930098, 7.100777, 7.271572, 7.442481, 7.613503, 7.784636, 
    7.955878, 8.127228, 8.298683, 8.470243, 8.641906, 8.813668, 8.985531, 
    9.15749, 9.329545, 9.501693, 9.673934, 9.846265, 10.01868, 10.19119, 
    10.36378, 10.53646, 10.70921, 10.88205, 11.05496, 11.22795, 11.40101, 
    11.57415, 11.74735, 11.92063, 12.09397, 12.26737, 12.44084, 12.61437, 
    12.78796, 12.96161, 13.13531, 13.30906, 13.48287, 13.65673, 13.83064, 
    14.00459, 14.17858, 14.35262, 14.5267, 14.70082, 14.87497, 15.04916, 
    15.22338, 15.39763, 15.57191, 15.74622, 15.92056, 16.09491, 16.26929, 
    16.44369, 16.6181, 16.79253, 16.96697, 17.14142, 17.31589, 17.49036, 
    17.66484, 17.83932, 18.0138, 18.18828, 18.36276, 18.53724, 18.71171, 
    18.88617, 19.06063, 19.23507, 19.40949, 19.5839, 19.7583, 19.93267, 
    20.10702, 20.28135, 20.45566, 20.62993, 20.80418, 20.9784, 21.15258, 
    21.32673, 21.50084, 21.67491, 21.84894, 22.02293, 22.19688, 22.37078, 
    22.54462, 22.71842, 22.89217, 23.06586, 23.2395, 23.41308, 23.5866, 
    23.76006, 23.93346, 24.10679, 24.28005, 24.45325, 24.62637, 24.79942, 
    24.9724, 25.1453, 25.31812, 25.49086, 25.66352, 25.8361, 26.0086, 26.181, 
    26.35332, 26.52554, 26.69768, 26.86972, 27.04166, 27.21351, 27.38526, 
    27.5569, 27.72845, 27.89988, 28.07122, 28.24244, 28.41356, 28.58456, 
    28.75545, 28.92623, 29.09689, 29.26743, 29.43786, 29.60816, 29.77834, 
    29.94839, 30.11832, 30.28812, 30.4578, 30.62734, 30.79675, 30.96603, 
    31.13517, 31.30417, 31.47304, 31.64176, 31.81035, 31.97879, 32.14709, 
    32.31524, 32.48324, 32.6511, 32.8188, 32.98635, 33.15376, 33.321, 
    33.48809, 33.65503, 33.8218, 33.98842, 34.15487, 34.32116, 34.48729, 
    34.65325, 34.81905, 34.98468, 35.15014, 35.31542, 35.48054, 35.64548, 
    35.81025, 35.97485, 36.13926, 36.3035, 36.46756, 36.63144, 36.79514, 
    36.95866, 37.12199, 37.28514, 37.4481, 37.61088, 37.77347, 37.93586, 
    38.09807, 38.26009, 38.42191, 38.58355, 38.74498, 38.90622, 39.06726, 
    39.22812, 39.38876, 39.54921, 39.70946, 39.86951, 40.02935, 40.189, 
    40.34843, 40.50767, 40.66669, 40.82552, 40.98413, 41.14254, 41.30073, 
    41.45872, 41.61649, 41.77406, 41.93141, 42.08855, 42.24547, 42.40218, 
    42.55867, 42.71495, 42.87101, 43.02685, 43.18248, 43.33788, 43.49307, 
    43.64803, 43.80278, 43.9573, 44.1116, 44.26568, 44.41954, 44.57317, 
    44.72657, 44.87975, 45.03271, 45.18544, 45.33794, 45.49021, 45.64226, 
    45.79408, 45.94567, 46.09703, 46.24816, 46.39906,
  -23.45163, -23.32268, -23.19349, -23.06407, -22.93441, -22.80452, 
    -22.67439, -22.54402, -22.41342, -22.28258, -22.1515, -22.02019, 
    -21.88864, -21.75685, -21.62482, -21.49256, -21.36005, -21.22731, 
    -21.09433, -20.96111, -20.82765, -20.69395, -20.56001, -20.42584, 
    -20.29142, -20.15676, -20.02186, -19.88672, -19.75134, -19.61572, 
    -19.47986, -19.34376, -19.20742, -19.07084, -18.93401, -18.79694, 
    -18.65964, -18.52209, -18.38429, -18.24626, -18.10799, -17.96947, 
    -17.83071, -17.69172, -17.55247, -17.41299, -17.27326, -17.1333, 
    -16.99309, -16.85264, -16.71194, -16.57101, -16.42983, -16.28841, 
    -16.14675, -16.00485, -15.86271, -15.72032, -15.5777, -15.43483, 
    -15.29172, -15.14837, -15.00478, -14.86095, -14.71687, -14.57256, 
    -14.42801, -14.28321, -14.13818, -13.9929, -13.84739, -13.70164, 
    -13.55565, -13.40941, -13.26294, -13.11623, -12.96929, -12.8221, 
    -12.67468, -12.52702, -12.37912, -12.23099, -12.08262, -11.93401, 
    -11.78516, -11.63609, -11.48677, -11.33722, -11.18744, -11.03742, 
    -10.88717, -10.73668, -10.58596, -10.43501, -10.28383, -10.13242, 
    -9.980772, -9.828896, -9.676789, -9.524453, -9.371888, -9.219094, 
    -9.066072, -8.912822, -8.759345, -8.605642, -8.451713, -8.297558, 
    -8.143178, -7.988575, -7.833747, -7.678697, -7.523425, -7.36793, 
    -7.212215, -7.05628, -6.900125, -6.743751, -6.587158, -6.430348, 
    -6.273322, -6.116079, -5.958622, -5.800949, -5.643063, -5.484964, 
    -5.326653, -5.16813, -5.009397, -4.850455, -4.691303, -4.531944, 
    -4.372377, -4.212605, -4.052627, -3.892445, -3.732059, -3.571471, 
    -3.410681, -3.249691, -3.0885, -2.927112, -2.765526, -2.603743, 
    -2.441764, -2.279591, -2.117224, -1.954665, -1.791915, -1.628974, 
    -1.465844, -1.302526, -1.13902, -0.975329, -0.8114531, -0.6473936, 
    -0.4831516, -0.3187284, -0.154125, 0.01065714, 0.175617, 0.3407533, 
    0.5060648, 0.6715503, 0.8372084, 1.003038, 1.169038, 1.335206, 1.501543, 
    1.668045, 1.834712, 2.001543, 2.168536, 2.33569, 2.503004, 2.670475, 
    2.838104, 3.005887, 3.173825, 3.341915, 3.510155, 3.678546, 3.847085, 
    4.01577, 4.184601, 4.353575, 4.522691, 4.691948, 4.861344, 5.030878, 
    5.200548, 5.370352, 5.540289, 5.710358, 5.880557, 6.050884, 6.221337, 
    6.391915, 6.562617, 6.73344, 6.904384, 7.075446, 7.246625, 7.417919, 
    7.589326, 7.760846, 7.932475, 8.104213, 8.276057, 8.448007, 8.620059, 
    8.792213, 8.964467, 9.13682, 9.309268, 9.481811, 9.654446, 9.827172, 
    9.999989, 10.17289, 10.34588, 10.51895, 10.69211, 10.86534, 11.03865, 
    11.21204, 11.38551, 11.55904, 11.73265, 11.90633, 12.08007, 12.25388, 
    12.42776, 12.60169, 12.77569, 12.94974, 13.12385, 13.29801, 13.47223, 
    13.64649, 13.8208, 13.99516, 14.16957, 14.34402, 14.5185, 14.69303, 
    14.86759, 15.04219, 15.21682, 15.39149, 15.56618, 15.7409, 15.91564, 
    16.09041, 16.2652, 16.44001, 16.61483, 16.78967, 16.96453, 17.13939, 
    17.31427, 17.48915, 17.66405, 17.83894, 18.01383, 18.18873, 18.36362, 
    18.53851, 18.71339, 18.88827, 19.06313, 19.23798, 19.41282, 19.58765, 
    19.76245, 19.93724, 20.112, 20.28674, 20.46146, 20.63614, 20.8108, 
    20.98543, 21.16002, 21.33458, 21.5091, 21.68358, 21.85802, 22.03242, 
    22.20677, 22.38108, 22.55534, 22.72954, 22.9037, 23.0778, 23.25184, 
    23.42583, 23.59975, 23.77361, 23.94741, 24.12115, 24.29481, 24.46841, 
    24.64194, 24.81539, 24.98877, 25.16207, 25.33529, 25.50843, 25.68149, 
    25.85447, 26.02735, 26.20016, 26.37287, 26.54549, 26.71802, 26.89045, 
    27.06279, 27.23503, 27.40716, 27.5792, 27.75113, 27.92296, 28.09468, 
    28.26629, 28.4378, 28.60918, 28.78046, 28.95162, 29.12267, 29.29359, 
    29.46439, 29.63508, 29.80563, 29.97607, 30.14637, 30.31655, 30.4866, 
    30.65652, 30.8263, 30.99595, 31.16546, 31.33484, 31.50407, 31.67316, 
    31.84212, 32.01092, 32.17958, 32.3481, 32.51647, 32.68468, 32.85275, 
    33.02066, 33.18842, 33.35603, 33.52347, 33.69076, 33.85789, 34.02486, 
    34.19166, 34.3583, 34.52478, 34.69109, 34.85723, 35.0232, 35.18901, 
    35.35464, 35.5201, 35.68538, 35.85049, 36.01542, 36.18018, 36.34475, 
    36.50914, 36.67336, 36.83739, 37.00124, 37.1649, 37.32837, 37.49166, 
    37.65476, 37.81767, 37.98039, 38.14292, 38.30526, 38.4674, 38.62935, 
    38.7911, 38.95266, 39.11401, 39.27517, 39.43613, 39.59689, 39.75744, 
    39.9178, 40.07795, 40.23789, 40.39763, 40.55717, 40.71649, 40.87561, 
    41.03452, 41.19322, 41.35171, 41.50999, 41.66805, 41.8259, 41.98354, 
    42.14097, 42.29818, 42.45517, 42.61194, 42.7685, 42.92484, 43.08096, 
    43.23686, 43.39254, 43.548, 43.70324, 43.85825, 44.01305, 44.16761, 
    44.32196, 44.47608, 44.62997, 44.78364, 44.93708, 45.09029, 45.24328, 
    45.39604, 45.54856, 45.70087, 45.85294, 46.00478, 46.15638, 46.30776, 
    46.45891,
  -23.52867, -23.3996, -23.27028, -23.14073, -23.01094, -22.88092, -22.75066, 
    -22.62016, -22.48942, -22.35845, -22.22724, -22.09579, -21.9641, 
    -21.83217, -21.7, -21.56759, -21.43495, -21.30206, -21.16893, -21.03557, 
    -20.90196, -20.76811, -20.63403, -20.4997, -20.36513, -20.23031, 
    -20.09526, -19.95997, -19.82443, -19.68865, -19.55263, -19.41637, 
    -19.27986, -19.14312, -19.00613, -18.86889, -18.73142, -18.5937, 
    -18.45574, -18.31754, -18.17909, -18.0404, -17.90147, -17.76229, 
    -17.62287, -17.48321, -17.34331, -17.20316, -17.06277, -16.92213, 
    -16.78125, -16.64013, -16.49877, -16.35716, -16.21531, -16.07321, 
    -15.93088, -15.7883, -15.64548, -15.50241, -15.3591, -15.21555, 
    -15.07176, -14.92773, -14.78345, -14.63893, -14.49417, -14.34917, 
    -14.20392, -14.05844, -13.91271, -13.76675, -13.62054, -13.47409, 
    -13.3274, -13.18047, -13.03331, -12.8859, -12.73825, -12.59037, 
    -12.44224, -12.29388, -12.14528, -11.99644, -11.84736, -11.69805, 
    -11.5485, -11.39872, -11.24869, -11.09844, -10.94794, -10.79722, 
    -10.64625, -10.49506, -10.34363, -10.19197, -10.04007, -9.887945, 
    -9.735586, -9.582996, -9.430176, -9.277125, -9.123845, -8.970336, 
    -8.816598, -8.662632, -8.508438, -8.354018, -8.199372, -8.044499, 
    -7.889403, -7.734081, -7.578536, -7.422768, -7.266777, -7.110565, 
    -6.954131, -6.797477, -6.640604, -6.483511, -6.3262, -6.168672, 
    -6.010927, -5.852966, -5.69479, -5.536399, -5.377795, -5.218979, 
    -5.05995, -4.90071, -4.741261, -4.581601, -4.421733, -4.261658, 
    -4.101376, -3.940888, -3.780195, -3.619299, -3.458199, -3.296898, 
    -3.135395, -2.973693, -2.811791, -2.649692, -2.487395, -2.324903, 
    -2.162215, -1.999334, -1.83626, -1.672994, -1.509538, -1.345893, 
    -1.182058, -1.018037, -0.8538297, -0.6894375, -0.5248615, -0.3601029, 
    -0.1951629, -0.03004281, 0.1352562, 0.300733, 0.4663863, 0.6322147, 
    0.7982172, 0.9643923, 1.130739, 1.297255, 1.463941, 1.630794, 1.797812, 
    1.964996, 2.132343, 2.299853, 2.467522, 2.635351, 2.803339, 2.971482, 
    3.139781, 3.308233, 3.476837, 3.645592, 3.814496, 3.983548, 4.152746, 
    4.322089, 4.491575, 4.661203, 4.830971, 5.000878, 5.170922, 5.341101, 
    5.511414, 5.68186, 5.852437, 6.023142, 6.193975, 6.364934, 6.536018, 
    6.707224, 6.878551, 7.049998, 7.221562, 7.393243, 7.565037, 7.736945, 
    7.908963, 8.081091, 8.253325, 8.425667, 8.598111, 8.770658, 8.943306, 
    9.116053, 9.288897, 9.461835, 9.634867, 9.807991, 9.981205, 10.15451, 
    10.3279, 10.50137, 10.67492, 10.84856, 11.02227, 11.19607, 11.36993, 
    11.54387, 11.71789, 11.89197, 12.06612, 12.24033, 12.41461, 12.58895, 
    12.76336, 12.93782, 13.11233, 13.2869, 13.46153, 13.6362, 13.81093, 
    13.9857, 14.16051, 14.33537, 14.51027, 14.68521, 14.86018, 15.03519, 
    15.21024, 15.38531, 15.56042, 15.73555, 15.91071, 16.08589, 16.26109, 
    16.43631, 16.61155, 16.78681, 16.96208, 17.13736, 17.31265, 17.48795, 
    17.66325, 17.83856, 18.01387, 18.18917, 18.36448, 18.53979, 18.71508, 
    18.89037, 19.06565, 19.24092, 19.41617, 19.59141, 19.76663, 19.94182, 
    20.117, 20.29216, 20.46728, 20.64238, 20.81745, 20.99249, 21.1675, 
    21.34247, 21.5174, 21.69229, 21.86714, 22.04195, 22.21671, 22.39143, 
    22.5661, 22.74071, 22.91528, 23.08978, 23.26423, 23.43863, 23.61296, 
    23.78723, 23.96144, 24.13557, 24.30964, 24.48365, 24.65758, 24.83143, 
    25.00521, 25.17891, 25.35254, 25.52608, 25.69954, 25.87291, 26.0462, 
    26.2194, 26.39251, 26.56553, 26.73845, 26.91128, 27.08401, 27.25664, 
    27.42917, 27.6016, 27.77393, 27.94614, 28.11826, 28.29026, 28.46214, 
    28.63392, 28.80558, 28.97713, 29.14856, 29.31987, 29.49105, 29.66212, 
    29.83306, 30.00387, 30.17455, 30.34511, 30.51554, 30.68583, 30.85599, 
    31.02601, 31.19589, 31.36564, 31.53524, 31.70471, 31.87403, 32.0432, 
    32.21223, 32.38111, 32.54984, 32.71843, 32.88685, 33.05513, 33.22324, 
    33.39121, 33.55901, 33.72665, 33.89414, 34.06146, 34.22862, 34.39561, 
    34.56244, 34.7291, 34.89558, 35.0619, 35.22805, 35.39403, 35.55983, 
    35.72546, 35.8909, 36.05618, 36.22127, 36.38618, 36.55091, 36.71545, 
    36.87982, 37.04399, 37.20799, 37.37179, 37.53541, 37.69883, 37.86207, 
    38.02511, 38.18796, 38.35062, 38.51308, 38.67535, 38.83741, 38.99929, 
    39.16096, 39.32243, 39.4837, 39.64476, 39.80563, 39.96629, 40.12674, 
    40.28699, 40.44704, 40.60687, 40.7665, 40.92591, 41.08512, 41.24411, 
    41.4029, 41.56147, 41.71983, 41.87797, 42.03589, 42.1936, 42.3511, 
    42.50837, 42.66543, 42.82227, 42.97889, 43.13529, 43.29147, 43.44742, 
    43.60316, 43.75867, 43.91395, 44.06901, 44.22385, 44.37846, 44.53284, 
    44.687, 44.84093, 44.99463, 45.14811, 45.30135, 45.45436, 45.60715, 
    45.7597, 45.91203, 46.06411, 46.21597, 46.3676, 46.51899,
  -23.60595, -23.47675, -23.34731, -23.21763, -23.08771, -22.95756, 
    -22.82717, -22.69654, -22.56566, -22.43456, -22.30321, -22.17162, 
    -22.03979, -21.90772, -21.77542, -21.64287, -21.51008, -21.37705, 
    -21.24378, -21.11027, -20.97651, -20.84252, -20.70828, -20.5738, 
    -20.43908, -20.30411, -20.1689, -20.03345, -19.89776, -19.76182, 
    -19.62564, -19.48922, -19.35255, -19.21564, -19.07849, -18.94109, 
    -18.80345, -18.66556, -18.52743, -18.38906, -18.25044, -18.11158, 
    -17.97247, -17.83312, -17.69352, -17.55368, -17.41359, -17.27326, 
    -17.13269, -16.99187, -16.85081, -16.7095, -16.56795, -16.42615, 
    -16.28411, -16.14182, -15.99929, -15.85652, -15.7135, -15.57024, 
    -15.42673, -15.28298, -15.13899, -14.99475, -14.85027, -14.70554, 
    -14.56057, -14.41536, -14.26991, -14.12421, -13.97828, -13.8321, 
    -13.68567, -13.53901, -13.3921, -13.24495, -13.09756, -12.94993, 
    -12.80206, -12.65395, -12.5056, -12.35701, -12.20818, -12.05911, 
    -11.9098, -11.76025, -11.61047, -11.46045, -11.31019, -11.15969, 
    -11.00896, -10.85798, -10.70678, -10.55534, -10.40366, -10.25175, 
    -10.09961, -9.947227, -9.794616, -9.641771, -9.488695, -9.335387, 
    -9.181848, -9.028078, -8.874079, -8.71985, -8.565392, -8.410706, 
    -8.255792, -8.100651, -7.945283, -7.78969, -7.633872, -7.477829, 
    -7.321561, -7.165071, -7.008358, -6.851424, -6.694268, -6.536892, 
    -6.379296, -6.221482, -6.063449, -5.905199, -5.746732, -5.588049, 
    -5.429152, -5.27004, -5.110714, -4.951177, -4.791428, -4.631467, 
    -4.471297, -4.310918, -4.150331, -3.989537, -3.828537, -3.667331, 
    -3.50592, -3.344307, -3.182491, -3.020473, -2.858256, -2.695838, 
    -2.533223, -2.37041, -2.207401, -2.044196, -1.880798, -1.717206, 
    -1.553423, -1.389448, -1.225284, -1.060932, -0.8963919, -0.7316657, 
    -0.5667545, -0.4016593, -0.2363815, -0.07092225, 0.09471726, 0.2605357, 
    0.426532, 0.5927048, 0.7590528, 0.9255747, 1.092269, 1.259135, 1.426171, 
    1.593376, 1.760747, 1.928285, 2.095988, 2.263854, 2.431881, 2.60007, 
    2.768417, 2.936921, 3.105582, 3.274398, 3.443367, 3.612488, 3.781759, 
    3.951179, 4.120746, 4.290459, 4.460317, 4.630317, 4.800458, 4.97074, 
    5.141159, 5.311715, 5.482406, 5.65323, 5.824186, 5.995273, 6.166488, 
    6.337829, 6.509296, 6.680887, 6.852599, 7.024432, 7.196383, 7.368452, 
    7.540636, 7.712933, 7.885342, 8.05786, 8.230488, 8.403222, 8.57606, 
    8.749002, 8.922046, 9.095188, 9.268429, 9.441766, 9.615196, 9.788719, 
    9.962333, 10.13604, 10.30982, 10.4837, 10.65766, 10.8317, 11.00582, 
    11.18001, 11.35428, 11.52863, 11.70305, 11.87754, 12.05209, 12.22672, 
    12.40141, 12.57616, 12.75097, 12.92584, 13.10076, 13.27575, 13.45078, 
    13.62587, 13.801, 13.97618, 14.15141, 14.32668, 14.502, 14.67735, 
    14.85274, 15.02816, 15.20362, 15.37911, 15.55463, 15.73018, 15.90575, 
    16.08134, 16.25696, 16.4326, 16.60826, 16.78393, 16.95961, 17.13531, 
    17.31101, 17.48673, 17.66245, 17.83817, 18.0139, 18.18962, 18.36535, 
    18.54107, 18.71678, 18.89248, 19.06818, 19.24386, 19.41953, 19.59518, 
    19.77082, 19.94643, 20.12203, 20.2976, 20.47314, 20.64865, 20.82414, 
    20.99959, 21.17501, 21.35039, 21.52574, 21.70105, 21.87631, 22.05153, 
    22.22671, 22.40183, 22.57691, 22.75194, 22.92691, 23.10183, 23.27669, 
    23.45149, 23.62623, 23.80091, 23.97552, 24.15007, 24.32455, 24.49895, 
    24.67329, 24.84755, 25.02173, 25.19584, 25.36987, 25.54381, 25.71767, 
    25.89145, 26.06514, 26.23874, 26.41224, 26.58566, 26.75898, 26.93221, 
    27.10533, 27.27836, 27.45129, 27.62411, 27.79683, 27.96944, 28.14194, 
    28.31433, 28.48661, 28.65877, 28.83082, 29.00276, 29.17457, 29.34626, 
    29.51784, 29.68928, 29.86061, 30.0318, 30.20287, 30.3738, 30.5446, 
    30.71527, 30.88581, 31.05621, 31.22647, 31.39658, 31.56656, 31.7364, 
    31.90609, 32.07563, 32.24503, 32.41428, 32.58337, 32.75232, 32.92111, 
    33.08974, 33.25822, 33.42654, 33.59471, 33.76271, 33.93055, 34.09823, 
    34.26574, 34.43309, 34.60026, 34.76727, 34.93411, 35.10078, 35.26727, 
    35.43359, 35.59974, 35.76571, 35.9315, 36.09711, 36.26254, 36.42779, 
    36.59285, 36.75774, 36.92243, 37.08694, 37.25127, 37.4154, 37.57934, 
    37.7431, 37.90666, 38.07003, 38.2332, 38.39618, 38.55896, 38.72154, 
    38.88393, 39.04612, 39.2081, 39.36988, 39.53147, 39.69284, 39.85402, 
    40.01498, 40.17575, 40.3363, 40.49665, 40.65678, 40.81671, 40.97643, 
    41.13593, 41.29522, 41.4543, 41.61316, 41.77181, 41.93024, 42.08846, 
    42.24646, 42.40424, 42.5618, 42.71914, 42.87626, 43.03316, 43.18984, 
    43.34629, 43.50253, 43.65854, 43.81432, 43.96988, 44.12521, 44.28031, 
    44.43519, 44.58984, 44.74426, 44.89845, 45.05242, 45.20615, 45.35965, 
    45.51292, 45.66597, 45.81877, 45.97135, 46.12369, 46.27579, 46.42767, 
    46.57931,
  -23.68347, -23.55414, -23.42457, -23.29477, -23.16472, -23.03444, 
    -22.90391, -22.77315, -22.64215, -22.5109, -22.37942, -22.2477, 
    -22.11573, -21.98352, -21.85108, -21.71839, -21.58546, -21.45228, 
    -21.31887, -21.18521, -21.05131, -20.91716, -20.78278, -20.64814, 
    -20.51327, -20.37815, -20.24279, -20.10718, -19.97133, -19.83524, 
    -19.6989, -19.56231, -19.42549, -19.28841, -19.15109, -19.01353, 
    -18.87572, -18.73767, -18.59937, -18.46082, -18.32203, -18.18299, 
    -18.04371, -17.90418, -17.76441, -17.62439, -17.48413, -17.34361, 
    -17.20286, -17.06186, -16.92061, -16.77911, -16.63737, -16.49538, 
    -16.35315, -16.21067, -16.06795, -15.92498, -15.78177, -15.63831, 
    -15.4946, -15.35065, -15.20646, -15.06202, -14.91733, -14.7724, 
    -14.62722, -14.4818, -14.33614, -14.19023, -14.04408, -13.89769, 
    -13.75105, -13.60417, -13.45704, -13.30967, -13.16206, -13.01421, 
    -12.86611, -12.71778, -12.5692, -12.42038, -12.27132, -12.12202, 
    -11.97248, -11.8227, -11.67268, -11.52242, -11.37192, -11.22118, 
    -11.0702, -10.91899, -10.76754, -10.61585, -10.46393, -10.31177, 
    -10.15937, -10.00674, -9.853878, -9.700779, -9.547446, -9.393881, 
    -9.240083, -9.086052, -8.93179, -8.777298, -8.622575, -8.467622, 
    -8.31244, -8.157029, -8.00139, -7.845525, -7.689433, -7.533114, -7.37657, 
    -7.219801, -7.062809, -6.905593, -6.748155, -6.590494, -6.432612, 
    -6.274511, -6.116189, -5.957649, -5.798891, -5.639915, -5.480723, 
    -5.321315, -5.161693, -5.001856, -4.841806, -4.681545, -4.521071, 
    -4.360388, -4.199495, -4.038393, -3.877084, -3.715568, -3.553846, 
    -3.391919, -3.229789, -3.067455, -2.90492, -2.742184, -2.579248, 
    -2.416114, -2.252782, -2.089253, -1.925529, -1.761611, -1.597499, 
    -1.433195, -1.2687, -1.104015, -0.939141, -0.7740797, -0.608832, 
    -0.4433991, -0.2777823, -0.1119826, 0.05399857, 0.2201601, 0.3865006, 
    0.5530189, 0.7197137, 0.8865837, 1.053628, 1.220844, 1.388232, 1.55579, 
    1.723516, 1.891409, 2.059469, 2.227692, 2.396079, 2.564628, 2.733336, 
    2.902204, 3.071229, 3.240409, 3.409745, 3.579233, 3.748872, 3.918662, 
    4.0886, 4.258685, 4.428915, 4.599289, 4.769806, 4.940464, 5.11126, 
    5.282194, 5.453264, 5.624469, 5.795806, 5.967274, 6.138872, 6.310598, 
    6.48245, 6.654427, 6.826527, 6.998747, 7.171088, 7.343545, 7.51612, 
    7.688808, 7.86161, 8.034522, 8.207543, 8.380672, 8.553906, 8.727245, 
    8.900685, 9.074226, 9.247866, 9.421601, 9.595433, 9.769357, 9.943373, 
    10.11748, 10.29167, 10.46595, 10.64031, 10.81475, 10.98928, 11.16388, 
    11.33856, 11.51331, 11.68814, 11.86304, 12.038, 12.21304, 12.38813, 
    12.5633, 12.73852, 12.9138, 13.08914, 13.26453, 13.43998, 13.61548, 
    13.79103, 13.96663, 14.14227, 14.31795, 14.49368, 14.66945, 14.84525, 
    15.02109, 15.19697, 15.37287, 15.54881, 15.72477, 15.90076, 16.07678, 
    16.25281, 16.42887, 16.60494, 16.78103, 16.95713, 17.13325, 17.30937, 
    17.48551, 17.66165, 17.83779, 18.01393, 18.19007, 18.36622, 18.54235, 
    18.71849, 18.89461, 19.07072, 19.24682, 19.42291, 19.59898, 19.77503, 
    19.95107, 20.12708, 20.30306, 20.47902, 20.65495, 20.83085, 21.00672, 
    21.18256, 21.35836, 21.53412, 21.70984, 21.88552, 22.06115, 22.23674, 
    22.41228, 22.58778, 22.76321, 22.9386, 23.11393, 23.2892, 23.46442, 
    23.63957, 23.81466, 23.98968, 24.16463, 24.33952, 24.51433, 24.68908, 
    24.86374, 25.03833, 25.21284, 25.38728, 25.56163, 25.73589, 25.91007, 
    26.08416, 26.25816, 26.43207, 26.60589, 26.77961, 26.95323, 27.12676, 
    27.30018, 27.4735, 27.64672, 27.81983, 27.99284, 28.16573, 28.33852, 
    28.51119, 28.68374, 28.85618, 29.0285, 29.2007, 29.37279, 29.54474, 
    29.71657, 29.88828, 30.05986, 30.23131, 30.40262, 30.5738, 30.74485, 
    30.91577, 31.08654, 31.25718, 31.42767, 31.59802, 31.76823, 31.93829, 
    32.10821, 32.27797, 32.44759, 32.61705, 32.78636, 32.95552, 33.12452, 
    33.29336, 33.46204, 33.63057, 33.79893, 33.96712, 34.13516, 34.30303, 
    34.47073, 34.63826, 34.80562, 34.97281, 35.13982, 35.30667, 35.47334, 
    35.63982, 35.80614, 35.97227, 36.13822, 36.30399, 36.46958, 36.63498, 
    36.8002, 36.96523, 37.13008, 37.29473, 37.4592, 37.62347, 37.78755, 
    37.95144, 38.11514, 38.27863, 38.44193, 38.60503, 38.76794, 38.93064, 
    39.09315, 39.25545, 39.41755, 39.57944, 39.74113, 39.90261, 40.06389, 
    40.22496, 40.38582, 40.54647, 40.70691, 40.86714, 41.02715, 41.18696, 
    41.34655, 41.50592, 41.66508, 41.82402, 41.98274, 42.14125, 42.29953, 
    42.4576, 42.61545, 42.77308, 42.93048, 43.08766, 43.24461, 43.40135, 
    43.55786, 43.71414, 43.8702, 44.02602, 44.18163, 44.337, 44.49215, 
    44.64706, 44.80175, 44.95621, 45.11043, 45.26443, 45.41819, 45.57172, 
    45.72501, 45.87807, 46.0309, 46.18349, 46.33585, 46.48798, 46.63986,
  -23.76123, -23.63177, -23.50208, -23.37214, -23.24197, -23.11156, -22.9809, 
    -22.85001, -22.71887, -22.5875, -22.45588, -22.32402, -22.19191, 
    -22.05957, -21.92698, -21.79415, -21.66108, -21.52776, -21.3942, 
    -21.2604, -21.12635, -20.99205, -20.85752, -20.72273, -20.58771, 
    -20.45244, -20.31692, -20.18116, -20.04515, -19.9089, -19.7724, 
    -19.63566, -19.49867, -19.36143, -19.22395, -19.08622, -18.94824, 
    -18.81002, -18.67155, -18.53283, -18.39387, -18.25466, -18.1152, 
    -17.9755, -17.83555, -17.69535, -17.5549, -17.41421, -17.27327, 
    -17.13209, -16.99065, -16.84897, -16.70704, -16.56487, -16.42244, 
    -16.27977, -16.13686, -15.99369, -15.85028, -15.70662, -15.56272, 
    -15.41857, -15.27417, -15.12953, -14.98464, -14.8395, -14.69412, 
    -14.54849, -14.40262, -14.2565, -14.11013, -13.96352, -13.81667, 
    -13.66957, -13.52223, -13.37464, -13.22681, -13.07873, -12.93041, 
    -12.78185, -12.63304, -12.48399, -12.3347, -12.18517, -12.0354, 
    -11.88538, -11.73512, -11.58462, -11.43389, -11.28291, -11.13169, 
    -10.98023, -10.82854, -10.67661, -10.52443, -10.37202, -10.21938, 
    -10.06649, -9.913376, -9.760022, -9.606432, -9.452608, -9.298551, 
    -9.144258, -8.989734, -8.834977, -8.679989, -8.524769, -8.369318, 
    -8.213637, -8.057727, -7.901588, -7.745221, -7.588626, -7.431805, 
    -7.274757, -7.117484, -6.959986, -6.802264, -6.644318, -6.48615, 
    -6.327761, -6.169149, -6.010318, -5.851268, -5.691998, -5.532511, 
    -5.372806, -5.212885, -5.052749, -4.892398, -4.731834, -4.571057, 
    -4.410068, -4.248868, -4.087458, -3.925839, -3.764011, -3.601977, 
    -3.439736, -3.27729, -3.11464, -2.951786, -2.788731, -2.625474, 
    -2.462017, -2.298361, -2.134507, -1.970456, -1.806209, -1.641768, 
    -1.477133, -1.312306, -1.147287, -0.9820786, -0.816681, -0.6510956, 
    -0.4853238, -0.3193666, -0.1532254, 0.01309873, 0.1796045, 0.3462905, 
    0.5131557, 0.6801986, 0.847418, 1.014813, 1.182381, 1.350122, 1.518034, 
    1.686116, 1.854367, 2.022784, 2.191367, 2.360115, 2.529025, 2.698097, 
    2.867328, 3.036719, 3.206266, 3.375969, 3.545825, 3.715835, 3.885996, 
    4.056306, 4.226764, 4.397369, 4.568119, 4.739012, 4.910047, 5.081223, 
    5.252536, 5.423987, 5.595573, 5.767293, 5.939146, 6.111129, 6.28324, 
    6.455479, 6.627843, 6.800332, 6.972942, 7.145673, 7.318522, 7.491489, 
    7.664571, 7.837766, 8.011073, 8.184491, 8.358016, 8.531648, 8.705385, 
    8.879225, 9.053165, 9.227205, 9.401342, 9.575576, 9.749903, 9.924321, 
    10.09883, 10.27343, 10.44811, 10.62288, 10.79773, 10.97266, 11.14767, 
    11.32276, 11.49793, 11.67316, 11.84847, 12.02385, 12.19929, 12.3748, 
    12.55037, 12.72601, 12.90171, 13.07746, 13.25327, 13.42913, 13.60504, 
    13.78101, 13.95702, 14.13308, 14.30918, 14.48533, 14.66151, 14.83773, 
    15.01399, 15.19029, 15.36661, 15.54296, 15.71935, 15.89576, 16.07219, 
    16.24865, 16.42512, 16.60161, 16.77812, 16.95465, 17.13118, 17.30773, 
    17.48428, 17.66084, 17.8374, 18.01397, 18.19053, 18.36709, 18.54365, 
    18.7202, 18.89675, 19.07328, 19.2498, 19.42631, 19.6028, 19.77927, 
    19.95572, 20.13215, 20.30856, 20.48493, 20.66128, 20.8376, 21.01389, 
    21.19014, 21.36636, 21.54254, 21.71868, 21.89477, 22.07082, 22.24683, 
    22.42278, 22.59869, 22.77455, 22.95035, 23.12609, 23.30178, 23.4774, 
    23.65297, 23.82847, 24.0039, 24.17927, 24.35456, 24.52979, 24.70494, 
    24.88001, 25.05501, 25.22993, 25.40477, 25.57952, 25.7542, 25.92878, 
    26.10328, 26.27768, 26.45199, 26.62621, 26.80033, 26.97436, 27.14828, 
    27.3221, 27.49582, 27.66944, 27.84295, 28.01635, 28.18964, 28.36282, 
    28.53588, 28.70883, 28.88166, 29.05437, 29.22696, 29.39943, 29.57178, 
    29.74399, 29.91608, 30.08805, 30.25988, 30.43158, 30.60314, 30.77457, 
    30.94586, 31.11702, 31.28803, 31.4589, 31.62963, 31.80021, 31.97064, 
    32.14093, 32.31107, 32.48105, 32.65089, 32.82056, 32.99009, 33.15945, 
    33.32866, 33.4977, 33.66659, 33.83531, 34.00387, 34.17226, 34.34048, 
    34.50854, 34.67642, 34.84414, 35.01168, 35.17905, 35.34624, 35.51325, 
    35.68009, 35.84674, 36.01322, 36.17952, 36.34563, 36.51156, 36.6773, 
    36.84286, 37.00822, 37.1734, 37.33839, 37.50319, 37.66779, 37.8322, 
    37.99642, 38.16044, 38.32426, 38.48788, 38.65131, 38.81454, 38.97756, 
    39.14038, 39.303, 39.46541, 39.62762, 39.78962, 39.95142, 40.113, 
    40.27438, 40.43555, 40.5965, 40.75725, 40.91778, 41.07809, 41.2382, 
    41.39808, 41.55775, 41.71721, 41.87644, 42.03546, 42.19426, 42.35283, 
    42.51118, 42.66932, 42.82723, 42.98491, 43.14238, 43.29961, 43.45663, 
    43.61341, 43.76997, 43.9263, 44.08241, 44.23828, 44.39392, 44.54934, 
    44.70452, 44.85947, 45.01419, 45.16868, 45.32294, 45.47696, 45.63074, 
    45.78429, 45.93761, 46.09069, 46.24354, 46.39615, 46.54852, 46.70065,
  -23.83922, -23.70964, -23.57982, -23.44976, -23.31946, -23.18892, 
    -23.05814, -22.92711, -22.79584, -22.66433, -22.53258, -22.40058, 
    -22.26834, -22.13585, -22.00313, -21.87016, -21.73694, -21.60348, 
    -21.46978, -21.33583, -21.20163, -21.06719, -20.9325, -20.79757, 
    -20.6624, -20.52697, -20.3913, -20.25538, -20.11922, -19.98281, 
    -19.84615, -19.70925, -19.57209, -19.43469, -19.29705, -19.15915, 
    -19.02101, -18.88262, -18.74398, -18.60509, -18.46596, -18.32658, 
    -18.18694, -18.04707, -17.90694, -17.76656, -17.62593, -17.48506, 
    -17.34394, -17.20257, -17.06095, -16.91908, -16.77696, -16.6346, 
    -16.49199, -16.34912, -16.20601, -16.06265, -15.91905, -15.77519, 
    -15.63109, -15.48674, -15.34214, -15.19729, -15.05219, -14.90685, 
    -14.76126, -14.61543, -14.46934, -14.32301, -14.17643, -14.02961, 
    -13.88254, -13.73522, -13.58766, -13.43985, -13.29179, -13.1435, 
    -12.99495, -12.84616, -12.69713, -12.54785, -12.39833, -12.24856, 
    -12.09856, -11.94831, -11.79781, -11.64708, -11.4961, -11.34488, 
    -11.19342, -11.04172, -10.88978, -10.7376, -10.58518, -10.43252, 
    -10.27962, -10.12648, -9.973111, -9.819501, -9.665654, -9.511571, 
    -9.357253, -9.2027, -9.047912, -8.89289, -8.737635, -8.582147, -8.426427, 
    -8.270475, -8.114293, -7.95788, -7.801238, -7.644366, -7.487267, 
    -7.329939, -7.172384, -7.014604, -6.856597, -6.698366, -6.539911, 
    -6.381233, -6.222332, -6.063209, -5.903865, -5.7443, -5.584517, 
    -5.424515, -5.264295, -5.103858, -4.943206, -4.782338, -4.621256, 
    -4.45996, -4.298452, -4.136733, -3.974803, -3.812664, -3.650315, 
    -3.487759, -3.324997, -3.162029, -2.998856, -2.835479, -2.6719, -2.50812, 
    -2.344139, -2.179958, -2.015579, -1.851004, -1.686232, -1.521265, 
    -1.356104, -1.190751, -1.025206, -0.859471, -0.6935469, -0.5274348, 
    -0.3611362, -0.1946521, -0.02798374, 0.1388675, 0.3059004, 0.4731137, 
    0.640506, 0.8080762, 0.9758228, 1.143745, 1.31184, 1.480108, 1.648547, 
    1.817156, 1.985933, 2.154877, 2.323987, 2.49326, 2.662696, 2.832293, 
    3.00205, 3.171966, 3.342038, 3.512265, 3.682646, 3.853179, 4.023863, 
    4.194696, 4.365677, 4.536804, 4.708076, 4.87949, 5.051045, 5.222741, 
    5.394574, 5.566544, 5.738648, 5.910886, 6.083255, 6.255754, 6.428382, 
    6.601136, 6.774014, 6.947016, 7.120139, 7.293382, 7.466743, 7.640219, 
    7.813811, 7.987514, 8.161329, 8.335253, 8.509284, 8.683421, 8.857661, 
    9.032004, 9.206447, 9.380987, 9.555624, 9.730356, 9.90518, 10.0801, 
    10.2551, 10.43019, 10.60537, 10.78063, 10.95597, 11.13139, 11.30689, 
    11.48246, 11.65811, 11.83383, 12.00962, 12.18548, 12.3614, 12.53739, 
    12.71344, 12.88955, 13.06572, 13.24195, 13.41823, 13.59456, 13.77094, 
    13.94737, 14.12385, 14.30037, 14.47693, 14.65354, 14.83018, 15.00686, 
    15.18357, 15.36032, 15.53709, 15.7139, 15.89073, 16.06758, 16.24446, 
    16.42135, 16.59827, 16.7752, 16.95214, 17.1291, 17.30607, 17.48305, 
    17.66003, 17.83701, 18.014, 18.19098, 18.36797, 18.54495, 18.72192, 
    18.89889, 19.07585, 19.25279, 19.42972, 19.60663, 19.78352, 19.9604, 
    20.13725, 20.31407, 20.49087, 20.66764, 20.84439, 21.02109, 21.19777, 
    21.3744, 21.551, 21.72756, 21.90407, 22.08054, 22.25696, 22.43334, 
    22.60966, 22.78593, 22.96215, 23.13831, 23.31441, 23.49045, 23.66643, 
    23.84234, 24.01819, 24.19397, 24.36968, 24.54531, 24.72088, 24.89636, 
    25.07177, 25.2471, 25.42235, 25.59751, 25.77259, 25.94758, 26.12248, 
    26.29729, 26.47201, 26.64663, 26.82115, 26.99558, 27.16991, 27.34413, 
    27.51825, 27.69227, 27.86617, 28.03997, 28.21366, 28.38723, 28.56069, 
    28.73403, 28.90725, 29.08036, 29.25334, 29.4262, 29.59893, 29.77154, 
    29.94402, 30.11637, 30.28859, 30.46067, 30.63262, 30.80443, 30.9761, 
    31.14763, 31.31903, 31.49027, 31.66138, 31.83234, 32.00315, 32.17381, 
    32.34431, 32.51467, 32.68488, 32.85492, 33.02481, 33.19455, 33.36412, 
    33.53353, 33.70277, 33.87186, 34.04078, 34.20953, 34.37811, 34.54652, 
    34.71476, 34.88283, 35.05072, 35.21844, 35.38599, 35.55335, 35.72054, 
    35.88754, 36.05436, 36.221, 36.38745, 36.55372, 36.71981, 36.8857, 
    37.05141, 37.21692, 37.38224, 37.54737, 37.71231, 37.87705, 38.0416, 
    38.20594, 38.37009, 38.53404, 38.69779, 38.86134, 39.02468, 39.18782, 
    39.35076, 39.51349, 39.67601, 39.83833, 40.00043, 40.16233, 40.32401, 
    40.48549, 40.64675, 40.8078, 40.96863, 41.12925, 41.28965, 41.44984, 
    41.60981, 41.76955, 41.92908, 42.08839, 42.24748, 42.40635, 42.56499, 
    42.72341, 42.88161, 43.03958, 43.19732, 43.35484, 43.51213, 43.6692, 
    43.82603, 43.98264, 44.13902, 44.29516, 44.45108, 44.60676, 44.76221, 
    44.91743, 45.07241, 45.22716, 45.38168, 45.53596, 45.69001, 45.84381, 
    45.99739, 46.15072, 46.30382, 46.45668, 46.6093, 46.76168,
  -23.91746, -23.78776, -23.65781, -23.52763, -23.3972, -23.26653, -23.13561, 
    -23.00445, -22.87305, -22.74141, -22.60952, -22.47739, -22.34501, 
    -22.21239, -22.07952, -21.94641, -21.81305, -21.67945, -21.5456, 
    -21.4115, -21.27716, -21.14258, -21.00774, -20.87266, -20.73733, 
    -20.60175, -20.46593, -20.32985, -20.19353, -20.05697, -19.92015, 
    -19.78308, -19.64577, -19.50821, -19.3704, -19.23234, -19.09403, 
    -18.95547, -18.81666, -18.6776, -18.5383, -18.39874, -18.25894, 
    -18.11888, -17.97857, -17.83802, -17.69721, -17.55616, -17.41485, 
    -17.2733, -17.13149, -16.98944, -16.84714, -16.70458, -16.56178, 
    -16.41872, -16.27542, -16.13186, -15.98806, -15.84401, -15.69971, 
    -15.55515, -15.41035, -15.2653, -15.12, -14.97445, -14.82866, -14.68261, 
    -14.53631, -14.38977, -14.24298, -14.09594, -13.94865, -13.80112, 
    -13.65334, -13.50531, -13.35703, -13.20851, -13.05974, -12.91072, 
    -12.76146, -12.61195, -12.4622, -12.3122, -12.16196, -12.01148, 
    -11.86074, -11.70977, -11.55855, -11.40709, -11.25539, -11.10345, 
    -10.95126, -10.79883, -10.64616, -10.49325, -10.3401, -10.18671, 
    -10.03308, -9.879218, -9.725114, -9.570771, -9.416192, -9.261376, 
    -9.106325, -8.951037, -8.795516, -8.639759, -8.483769, -8.327546, 
    -8.171091, -8.014403, -7.857485, -7.700336, -7.542958, -7.38535, 
    -7.227513, -7.069449, -6.911158, -6.75264, -6.593897, -6.434929, 
    -6.275737, -6.116322, -5.956684, -5.796824, -5.636744, -5.476443, 
    -5.315923, -5.155185, -4.994229, -4.833057, -4.671669, -4.510067, 
    -4.34825, -4.18622, -4.023978, -3.861526, -3.698863, -3.535991, 
    -3.372911, -3.209624, -3.04613, -2.882432, -2.71853, -2.554425, 
    -2.390117, -2.225609, -2.060902, -1.895995, -1.730892, -1.565592, 
    -1.400096, -1.234407, -1.068525, -0.9024514, -0.7361872, -0.5697338, 
    -0.4030923, -0.2362641, -0.06925032, 0.0979477, 0.2653287, 0.4328915, 
    0.6006346, 0.7685568, 0.9366568, 1.104933, 1.273385, 1.44201, 1.610807, 
    1.779776, 1.948914, 2.11822, 2.287693, 2.457331, 2.627133, 2.797098, 
    2.967223, 3.137508, 3.30795, 3.47855, 3.649304, 3.820211, 3.991271, 
    4.16248, 4.333838, 4.505344, 4.676995, 4.84879, 5.020728, 5.192806, 
    5.365024, 5.537378, 5.709869, 5.882494, 6.055252, 6.22814, 6.401157, 
    6.574302, 6.747573, 6.920968, 7.094485, 7.268123, 7.441879, 7.615753, 
    7.789742, 7.963844, 8.138058, 8.312383, 8.486814, 8.661353, 8.835997, 
    9.010742, 9.185589, 9.360535, 9.535578, 9.710716, 9.885947, 10.06127, 
    10.23668, 10.41218, 10.58777, 10.76344, 10.93919, 11.11503, 11.29094, 
    11.46693, 11.64299, 11.81912, 11.99533, 12.1716, 12.34794, 12.52435, 
    12.70081, 12.87734, 13.05393, 13.23057, 13.40727, 13.58402, 13.76082, 
    13.93767, 14.11457, 14.29151, 14.4685, 14.64552, 14.82259, 14.99969, 
    15.17682, 15.35399, 15.53119, 15.70842, 15.88567, 16.06295, 16.24025, 
    16.41757, 16.59491, 16.77226, 16.94963, 17.12701, 17.30441, 17.48181, 
    17.65921, 17.83662, 18.01403, 18.19144, 18.36885, 18.54626, 18.72366, 
    18.90105, 19.07843, 19.25579, 19.43315, 19.61048, 19.7878, 19.9651, 
    20.14237, 20.31962, 20.49684, 20.67404, 20.8512, 21.02833, 21.20542, 
    21.38248, 21.5595, 21.73648, 21.91341, 22.0903, 22.26715, 22.44394, 
    22.62068, 22.79737, 22.97401, 23.15059, 23.3271, 23.50356, 23.67996, 
    23.85629, 24.03255, 24.20874, 24.38487, 24.56092, 24.73689, 24.91279, 
    25.08861, 25.26435, 25.44001, 25.61558, 25.79107, 25.96647, 26.14178, 
    26.31699, 26.49212, 26.66714, 26.84208, 27.01691, 27.19164, 27.36626, 
    27.54078, 27.7152, 27.88951, 28.0637, 28.23779, 28.41176, 28.58561, 
    28.75935, 28.93297, 29.10647, 29.27984, 29.45309, 29.62622, 29.79922, 
    29.97208, 30.14482, 30.31742, 30.48989, 30.66223, 30.83442, 31.00648, 
    31.17839, 31.35017, 31.5218, 31.69328, 31.86461, 32.0358, 32.20683, 
    32.37772, 32.54845, 32.71902, 32.88944, 33.0597, 33.2298, 33.39974, 
    33.56952, 33.73912, 33.90857, 34.07785, 34.24696, 34.4159, 34.58467, 
    34.75327, 34.9217, 35.08995, 35.25802, 35.42591, 35.59363, 35.76116, 
    35.92851, 36.09568, 36.26266, 36.42947, 36.59608, 36.7625, 36.92873, 
    37.09478, 37.26063, 37.42629, 37.59175, 37.75702, 37.92209, 38.08697, 
    38.25164, 38.41612, 38.5804, 38.74447, 38.90834, 39.07201, 39.23547, 
    39.39872, 39.56177, 39.72461, 39.88724, 40.04966, 40.21186, 40.37386, 
    40.53564, 40.69721, 40.85857, 41.0197, 41.18063, 41.34133, 41.50182, 
    41.66208, 41.82212, 41.98195, 42.14155, 42.30093, 42.46009, 42.61902, 
    42.77773, 42.93621, 43.09447, 43.25249, 43.4103, 43.56787, 43.72521, 
    43.88232, 44.0392, 44.19585, 44.35227, 44.50846, 44.66441, 44.82013, 
    44.97562, 45.13087, 45.28588, 45.44066, 45.5952, 45.74951, 45.90357, 
    46.0574, 46.21099, 46.36435, 46.51746, 46.67033, 46.82296,
  -23.99595, -23.86612, -23.73605, -23.60573, -23.47518, -23.34438, 
    -23.21333, -23.08204, -22.95051, -22.81873, -22.68671, -22.55444, 
    -22.42193, -22.28917, -22.15616, -22.02291, -21.88941, -21.75567, 
    -21.62167, -21.48743, -21.35295, -21.21821, -21.08323, -20.94799, 
    -20.81251, -20.67678, -20.54081, -20.40458, -20.2681, -20.13138, 
    -19.9944, -19.85718, -19.7197, -19.58198, -19.444, -19.30577, -19.1673, 
    -19.02857, -18.8896, -18.75037, -18.61089, -18.47116, -18.33118, 
    -18.19095, -18.05046, -17.90973, -17.76875, -17.62751, -17.48602, 
    -17.34428, -17.20229, -17.06005, -16.91756, -16.77481, -16.63182, 
    -16.48857, -16.34508, -16.20133, -16.05733, -15.91308, -15.76857, 
    -15.62382, -15.47882, -15.33356, -15.18806, -15.0423, -14.8963, 
    -14.75004, -14.60354, -14.45678, -14.30978, -14.16252, -14.01502, 
    -13.86727, -13.71926, -13.57101, -13.42251, -13.27377, -13.12477, 
    -12.97553, -12.82604, -12.6763, -12.52632, -12.37609, -12.22561, 
    -12.07489, -11.92392, -11.77271, -11.62125, -11.46955, -11.31761, 
    -11.16541, -11.01298, -10.86031, -10.70739, -10.55423, -10.40083, 
    -10.24718, -10.0933, -9.939177, -9.784813, -9.630211, -9.47537, 
    -9.320292, -9.164975, -9.009422, -8.853633, -8.697607, -8.541347, 
    -8.384851, -8.228123, -8.07116, -7.913965, -7.756538, -7.59888, -7.44099, 
    -7.282871, -7.124523, -6.965946, -6.807141, -6.648109, -6.488851, 
    -6.329367, -6.169658, -6.009726, -5.84957, -5.689191, -5.528592, 
    -5.367771, -5.206731, -5.045471, -4.883994, -4.722299, -4.560388, 
    -4.398262, -4.235921, -4.073367, -3.910599, -3.747621, -3.584432, 
    -3.421033, -3.257426, -3.093612, -2.92959, -2.765364, -2.600933, 
    -2.436298, -2.271462, -2.106424, -1.941186, -1.77575, -1.610115, 
    -1.444284, -1.278258, -1.112037, -0.9456236, -0.7790182, -0.6122221, 
    -0.4452366, -0.278063, -0.1107025, 0.05684358, 0.224574, 0.3924875, 
    0.5605827, 0.7288583, 0.897313, 1.065945, 1.234754, 1.403738, 1.572895, 
    1.742225, 1.911726, 2.081395, 2.251233, 2.421237, 2.591407, 2.76174, 
    2.932235, 3.102891, 3.273706, 3.444678, 3.615807, 3.78709, 3.958526, 
    4.130114, 4.301852, 4.473737, 4.64577, 4.817947, 4.990268, 5.162731, 
    5.335334, 5.508076, 5.680954, 5.853969, 6.027116, 6.200395, 6.373805, 
    6.547342, 6.721007, 6.894796, 7.068709, 7.242743, 7.416898, 7.59117, 
    7.765558, 7.940061, 8.114676, 8.289402, 8.464237, 8.63918, 8.814228, 
    8.989379, 9.164632, 9.339985, 9.515435, 9.690982, 9.866623, 10.04236, 
    10.21818, 10.39409, 10.57009, 10.74617, 10.92234, 11.09859, 11.27491, 
    11.45131, 11.62779, 11.80434, 11.98097, 12.15766, 12.33441, 12.51124, 
    12.68812, 12.86507, 13.04208, 13.21914, 13.39626, 13.57343, 13.75066, 
    13.92793, 14.10525, 14.28261, 14.46002, 14.63747, 14.81496, 14.99248, 
    15.17004, 15.34764, 15.52526, 15.70291, 15.88059, 16.05829, 16.23602, 
    16.41376, 16.59153, 16.76931, 16.94711, 17.12491, 17.30273, 17.48056, 
    17.65839, 17.83623, 18.01406, 18.1919, 18.36974, 18.54757, 18.7254, 
    18.90321, 19.08102, 19.25881, 19.43659, 19.61435, 19.7921, 19.96982, 
    20.14752, 20.32519, 20.50284, 20.68046, 20.85805, 21.0356, 21.21312, 
    21.3906, 21.56804, 21.74545, 21.9228, 22.10011, 22.27738, 22.4546, 
    22.63176, 22.80887, 22.98592, 23.16292, 23.33986, 23.51674, 23.69355, 
    23.8703, 24.04698, 24.22359, 24.40013, 24.57659, 24.75299, 24.9293, 
    25.10553, 25.28168, 25.45776, 25.63374, 25.80964, 25.98545, 26.16117, 
    26.33679, 26.51233, 26.68776, 26.8631, 27.03833, 27.21347, 27.3885, 
    27.56343, 27.73824, 27.91295, 28.08755, 28.26204, 28.43641, 28.61066, 
    28.78479, 28.95881, 29.1327, 29.30647, 29.48012, 29.65364, 29.82702, 
    30.00028, 30.17341, 30.3464, 30.51926, 30.69198, 30.86456, 31.037, 
    31.2093, 31.38145, 31.55346, 31.72532, 31.89704, 32.0686, 32.24001, 
    32.41127, 32.58238, 32.75333, 32.92411, 33.09475, 33.26521, 33.43552, 
    33.60567, 33.77564, 33.94545, 34.1151, 34.28457, 34.45387, 34.623, 
    34.79196, 34.96074, 35.12934, 35.29777, 35.46602, 35.63409, 35.80197, 
    35.96967, 36.13719, 36.30452, 36.47166, 36.63862, 36.80539, 36.97196, 
    37.13834, 37.30453, 37.47053, 37.63633, 37.80193, 37.96734, 38.13254, 
    38.29755, 38.46235, 38.62696, 38.79136, 38.95555, 39.11954, 39.28332, 
    39.4469, 39.61026, 39.77341, 39.93636, 40.09909, 40.26162, 40.42392, 
    40.58601, 40.74789, 40.90955, 41.071, 41.23222, 41.39323, 41.55401, 
    41.71458, 41.87492, 42.03504, 42.19493, 42.35461, 42.51406, 42.67328, 
    42.83228, 42.99105, 43.14959, 43.3079, 43.46598, 43.62383, 43.78146, 
    43.93885, 44.096, 44.25293, 44.40962, 44.56608, 44.72231, 44.87829, 
    45.03404, 45.18956, 45.34484, 45.49988, 45.65468, 45.80925, 45.96357, 
    46.11766, 46.2715, 46.42511, 46.57847, 46.73159, 46.88447,
  -24.07468, -23.94472, -23.81453, -23.68409, -23.5534, -23.42248, -23.2913, 
    -23.15988, -23.02822, -22.89631, -22.76415, -22.63175, -22.4991, 
    -22.3662, -22.23306, -22.09966, -21.96602, -21.83213, -21.698, -21.56361, 
    -21.42898, -21.29409, -21.15896, -21.02358, -20.88795, -20.75207, 
    -20.61594, -20.47955, -20.34292, -20.20604, -20.0689, -19.93152, 
    -19.79388, -19.65599, -19.51785, -19.37947, -19.24082, -19.10193, 
    -18.96278, -18.82338, -18.68373, -18.54383, -18.40368, -18.26327, 
    -18.12261, -17.9817, -17.84053, -17.69911, -17.55744, -17.41552, 
    -17.27335, -17.13092, -16.98824, -16.8453, -16.70212, -16.55868, 
    -16.41499, -16.27104, -16.12685, -15.9824, -15.8377, -15.69274, 
    -15.54754, -15.40208, -15.25637, -15.11041, -14.96419, -14.81773, 
    -14.67101, -14.52404, -14.37683, -14.22936, -14.08164, -13.93366, 
    -13.78544, -13.63697, -13.48825, -13.33928, -13.19006, -13.04059, 
    -12.89087, -12.7409, -12.59069, -12.44022, -12.28951, -12.13856, 
    -11.98735, -11.8359, -11.6842, -11.53226, -11.38007, -11.22763, 
    -11.07495, -10.92203, -10.76886, -10.61545, -10.46179, -10.3079, 
    -10.15376, -9.999375, -9.844753, -9.689891, -9.534788, -9.379446, 
    -9.223865, -9.068045, -8.911987, -8.755692, -8.599161, -8.442393, 
    -8.28539, -8.128152, -7.970679, -7.812973, -7.655035, -7.496864, 
    -7.338461, -7.179828, -7.020964, -6.861871, -6.70255, -6.543001, 
    -6.383224, -6.223221, -6.062993, -5.90254, -5.741863, -5.580963, 
    -5.419841, -5.258497, -5.096933, -4.93515, -4.773147, -4.610927, 
    -4.44849, -4.285837, -4.122969, -3.959887, -3.796592, -3.633085, 
    -3.469367, -3.305438, -3.141301, -2.976956, -2.812404, -2.647646, 
    -2.482683, -2.317517, -2.152148, -1.986577, -1.820807, -1.654837, 
    -1.488669, -1.322304, -1.155744, -0.9889893, -0.8220413, -0.6549014, 
    -0.4875706, -0.3200504, -0.1523419, 0.01555362, 0.1836348, 0.3519003, 
    0.520349, 0.6889793, 0.8577901, 1.02678, 1.195947, 1.365291, 1.53481, 
    1.704502, 1.874366, 2.044401, 2.214606, 2.384978, 2.555516, 2.726219, 
    2.897085, 3.068114, 3.239302, 3.41065, 3.582155, 3.753815, 3.92563, 
    4.097597, 4.269715, 4.441983, 4.614398, 4.78696, 4.959666, 5.132515, 
    5.305506, 5.478636, 5.651904, 5.825308, 5.998847, 6.172519, 6.346322, 
    6.520255, 6.694314, 6.868501, 7.042811, 7.217244, 7.391798, 7.56647, 
    7.74126, 7.916164, 8.091183, 8.266313, 8.441553, 8.6169, 8.792355, 
    8.967913, 9.143574, 9.319336, 9.495195, 9.671153, 9.847205, 10.02335, 
    10.19959, 10.37591, 10.55232, 10.72882, 10.9054, 11.08207, 11.25881, 
    11.43563, 11.61252, 11.78949, 11.96653, 12.14364, 12.32082, 12.49807, 
    12.67537, 12.85274, 13.03017, 13.20766, 13.3852, 13.56279, 13.74044, 
    13.91814, 14.09588, 14.27367, 14.45151, 14.62938, 14.80729, 14.98524, 
    15.16323, 15.34125, 15.5193, 15.69738, 15.87548, 16.05362, 16.23177, 
    16.40994, 16.58814, 16.76635, 16.94457, 17.12281, 17.30105, 17.47931, 
    17.65757, 17.83583, 18.0141, 18.19237, 18.37063, 18.54889, 18.72714, 
    18.90539, 19.08362, 19.26184, 19.44005, 19.61824, 19.79641, 19.97456, 
    20.15269, 20.33079, 20.50887, 20.68691, 20.86493, 21.04291, 21.22085, 
    21.39876, 21.57663, 21.75445, 21.93224, 22.10997, 22.28766, 22.4653, 
    22.64289, 22.82042, 22.9979, 23.17532, 23.35268, 23.52998, 23.70721, 
    23.88438, 24.06148, 24.23851, 24.41546, 24.59235, 24.76916, 24.94588, 
    25.12253, 25.2991, 25.47559, 25.65199, 25.8283, 26.00452, 26.18065, 
    26.35669, 26.53263, 26.70847, 26.88422, 27.05986, 27.23541, 27.41084, 
    27.58617, 27.7614, 27.93651, 28.11151, 28.2864, 28.46117, 28.63582, 
    28.81036, 28.98477, 29.15906, 29.33323, 29.50727, 29.68118, 29.85496, 
    30.02861, 30.20213, 30.37551, 30.54876, 30.72187, 30.89484, 31.06766, 
    31.24035, 31.41289, 31.58528, 31.75752, 31.92962, 32.10156, 32.27335, 
    32.44498, 32.61647, 32.78779, 32.95895, 33.12996, 33.30079, 33.47147, 
    33.64198, 33.81233, 33.98251, 34.15252, 34.32235, 34.49202, 34.66151, 
    34.83083, 34.99996, 35.16893, 35.33771, 35.50631, 35.67473, 35.84296, 
    36.01102, 36.17888, 36.34656, 36.51405, 36.68135, 36.84846, 37.01538, 
    37.18211, 37.34863, 37.51497, 37.6811, 37.84704, 38.01278, 38.17832, 
    38.34366, 38.50879, 38.67372, 38.83845, 39.00297, 39.16728, 39.33138, 
    39.49528, 39.65896, 39.82244, 39.9857, 40.14875, 40.31158, 40.4742, 
    40.6366, 40.79879, 40.96075, 41.12251, 41.28403, 41.44534, 41.60643, 
    41.7673, 41.92794, 42.08835, 42.24855, 42.40851, 42.56825, 42.72777, 
    42.88705, 43.04611, 43.20494, 43.36353, 43.5219, 43.68003, 43.83794, 
    43.99561, 44.15304, 44.31024, 44.46721, 44.62394, 44.78043, 44.93669, 
    45.09271, 45.24849, 45.40403, 45.55934, 45.71441, 45.86923, 46.02381, 
    46.17815, 46.33226, 46.48611, 46.63973, 46.7931, 46.94623,
  -24.15365, -24.02357, -23.89326, -23.76269, -23.63188, -23.50082, 
    -23.36952, -23.23797, -23.10617, -22.97413, -22.84184, -22.7093, 
    -22.57651, -22.44348, -22.3102, -22.17666, -22.04288, -21.90885, 
    -21.77457, -21.64004, -21.50526, -21.37023, -21.23495, -21.09942, 
    -20.96364, -20.8276, -20.69132, -20.55478, -20.41799, -20.28095, 
    -20.14366, -20.00611, -19.86832, -19.73027, -19.59196, -19.45341, 
    -19.3146, -19.17554, -19.03622, -18.89665, -18.75683, -18.61676, 
    -18.47643, -18.33584, -18.19501, -18.05392, -17.91257, -17.77097, 
    -17.62912, -17.48701, -17.34465, -17.20204, -17.05917, -16.91605, 
    -16.77267, -16.62904, -16.48515, -16.34101, -16.19662, -16.05197, 
    -15.90707, -15.76192, -15.61651, -15.47085, -15.32493, -15.17877, 
    -15.03234, -14.88567, -14.73874, -14.59156, -14.44413, -14.29644, 
    -14.14851, -14.00032, -13.85187, -13.70318, -13.55424, -13.40504, 
    -13.2556, -13.1059, -12.95595, -12.80575, -12.65531, -12.50461, 
    -12.35366, -12.20247, -12.05103, -11.89933, -11.74739, -11.59521, 
    -11.44277, -11.29009, -11.13717, -10.98399, -10.83058, -10.67691, 
    -10.523, -10.36885, -10.21446, -10.05982, -9.904937, -9.749813, 
    -9.594448, -9.438842, -9.282995, -9.126908, -8.970582, -8.814016, 
    -8.657213, -8.500173, -8.342895, -8.18538, -8.027629, -7.869644, 
    -7.711424, -7.55297, -7.394284, -7.235365, -7.076214, -6.916832, 
    -6.757221, -6.59738, -6.43731, -6.277012, -6.116488, -5.955736, -5.79476, 
    -5.633559, -5.472134, -5.310486, -5.148617, -4.986526, -4.824215, 
    -4.661685, -4.498936, -4.33597, -4.172787, -4.009389, -3.845777, 
    -3.68195, -3.517911, -3.353661, -3.1892, -3.02453, -2.859652, -2.694566, 
    -2.529274, -2.363776, -2.198075, -2.032171, -1.866065, -1.699758, 
    -1.533252, -1.366548, -1.199647, -1.03255, -0.8652583, -0.6977732, 
    -0.5300959, -0.3622277, -0.1941699, -0.02592372, 0.1425095, 0.3111284, 
    0.4799318, 0.6489183, 0.8180864, 0.987435, 1.156963, 1.326668, 1.496549, 
    1.666605, 1.836835, 2.007236, 2.177809, 2.34855, 2.519458, 2.690533, 
    2.861772, 3.033175, 3.204738, 3.376462, 3.548345, 3.720384, 3.892579, 
    4.064927, 4.237428, 4.410079, 4.582879, 4.755826, 4.92892, 5.102157, 
    5.275537, 5.449057, 5.622716, 5.796513, 5.970445, 6.144511, 6.318709, 
    6.493038, 6.667495, 6.84208, 7.016789, 7.191623, 7.366577, 7.541652, 
    7.716845, 7.892153, 8.067576, 8.243113, 8.418758, 8.594514, 8.770376, 
    8.946344, 9.122415, 9.298587, 9.474858, 9.651228, 9.827693, 10.00425, 
    10.1809, 10.35764, 10.53447, 10.71139, 10.88838, 11.06546, 11.24263, 
    11.41986, 11.59718, 11.77457, 11.95203, 12.12956, 12.30716, 12.48483, 
    12.66256, 12.84035, 13.0182, 13.19612, 13.37408, 13.5521, 13.73018, 
    13.9083, 14.08647, 14.26469, 14.44295, 14.62125, 14.79959, 14.97797, 
    15.15638, 15.33483, 15.51331, 15.69182, 15.87035, 16.04892, 16.2275, 
    16.4061, 16.58473, 16.76336, 16.94202, 17.12069, 17.29936, 17.47805, 
    17.65674, 17.83544, 18.01413, 18.19283, 18.37153, 18.55022, 18.7289, 
    18.90758, 19.08624, 19.26489, 19.44353, 19.62215, 19.80075, 19.97933, 
    20.15789, 20.33642, 20.51492, 20.6934, 20.87184, 21.05025, 21.22862, 
    21.40696, 21.58525, 21.76351, 21.94172, 22.11988, 22.29799, 22.47606, 
    22.65407, 22.83203, 23.00993, 23.18778, 23.36556, 23.54328, 23.72093, 
    23.89852, 24.07605, 24.2535, 24.43087, 24.60818, 24.7854, 24.96255, 
    25.13962, 25.3166, 25.49351, 25.67032, 25.84705, 26.02368, 26.20023, 
    26.37668, 26.55303, 26.72929, 26.90544, 27.0815, 27.25745, 27.43329, 
    27.60903, 27.78466, 27.96018, 28.13559, 28.31088, 28.48605, 28.66111, 
    28.83604, 29.01085, 29.18554, 29.36011, 29.53455, 29.70885, 29.88303, 
    30.05708, 30.23099, 30.40476, 30.5784, 30.7519, 30.92526, 31.09847, 
    31.27154, 31.44447, 31.61724, 31.78987, 31.96235, 32.13467, 32.30684, 
    32.47886, 32.65071, 32.82241, 32.99395, 33.16533, 33.33654, 33.50759, 
    33.67847, 33.84919, 34.01973, 34.19011, 34.36031, 34.53033, 34.70019, 
    34.86987, 35.03936, 35.20869, 35.37783, 35.54678, 35.71556, 35.88415, 
    36.05255, 36.22077, 36.38879, 36.55663, 36.72428, 36.89174, 37.05899, 
    37.22606, 37.39293, 37.5596, 37.72608, 37.89235, 38.05843, 38.2243, 
    38.38997, 38.55544, 38.72069, 38.88575, 39.05059, 39.21523, 39.37966, 
    39.54387, 39.70788, 39.87167, 40.03525, 40.19862, 40.36176, 40.5247, 
    40.68741, 40.8499, 41.01218, 41.17424, 41.33607, 41.49768, 41.65907, 
    41.82024, 41.98118, 42.1419, 42.30238, 42.46265, 42.62268, 42.78248, 
    42.94206, 43.10141, 43.26052, 43.4194, 43.57805, 43.73647, 43.89465, 
    44.0526, 44.21031, 44.36779, 44.52503, 44.68203, 44.8388, 44.99533, 
    45.15162, 45.30766, 45.46347, 45.61904, 45.77437, 45.92945, 46.0843, 
    46.2389, 46.39325, 46.54737, 46.70124, 46.85486, 47.00824,
  -24.23287, -24.10267, -23.97223, -23.84154, -23.7106, -23.57942, -23.44798, 
    -23.31631, -23.18438, -23.0522, -22.91978, -22.78711, -22.65418, 
    -22.52101, -22.38759, -22.25392, -22.12, -21.98582, -21.8514, -21.71673, 
    -21.5818, -21.44662, -21.3112, -21.17551, -21.03958, -20.90339, 
    -20.76696, -20.63026, -20.49332, -20.35612, -20.21867, -20.08097, 
    -19.94301, -19.8048, -19.66633, -19.52761, -19.38864, -19.2494, 
    -19.10992, -18.97018, -18.83019, -18.68994, -18.54944, -18.40868, 
    -18.26766, -18.12639, -17.98487, -17.84309, -17.70106, -17.55877, 
    -17.41622, -17.27342, -17.13036, -16.98705, -16.84348, -16.69966, 
    -16.55558, -16.41124, -16.26665, -16.12181, -15.97671, -15.83135, 
    -15.68574, -15.53988, -15.39375, -15.24738, -15.10075, -14.95387, 
    -14.80673, -14.65933, -14.51169, -14.36379, -14.21563, -14.06722, 
    -13.91856, -13.76965, -13.62048, -13.47106, -13.32139, -13.17146, 
    -13.02129, -12.87086, -12.72018, -12.56925, -12.41807, -12.26663, 
    -12.11495, -11.96302, -11.81084, -11.65841, -11.50573, -11.35281, 
    -11.19963, -11.04621, -10.89254, -10.73862, -10.58446, -10.43006, 
    -10.2754, -10.12051, -9.965365, -9.80998, -9.654352, -9.498481, 
    -9.342368, -9.186013, -9.029418, -8.872581, -8.715506, -8.558191, 
    -8.400638, -8.242846, -8.084817, -7.926551, -7.76805, -7.609313, 
    -7.450341, -7.291136, -7.131697, -6.972026, -6.812123, -6.651989, 
    -6.491626, -6.331032, -6.17021, -6.009161, -5.847884, -5.686381, 
    -5.524652, -5.3627, -5.200524, -5.038125, -4.875504, -4.712663, 
    -4.549602, -4.386322, -4.222824, -4.059108, -3.895177, -3.73103, 
    -3.56667, -3.402097, -3.237311, -3.072315, -2.907109, -2.741694, 
    -2.576071, -2.410242, -2.244207, -2.077968, -1.911526, -1.744881, 
    -1.578036, -1.410991, -1.243748, -1.076307, -0.9086705, -0.740839, 
    -0.5728139, -0.4045965, -0.2361881, -0.06758997, 0.1011966, 0.2701703, 
    0.4393298, 0.6086737, 0.7782007, 0.9479094, 1.117798, 1.287866, 1.458112, 
    1.628534, 1.79913, 1.9699, 2.140841, 2.311953, 2.483233, 2.654681, 
    2.826294, 2.998072, 3.170013, 3.342115, 3.514377, 3.686796, 3.859373, 
    4.032104, 4.204988, 4.378025, 4.551211, 4.724546, 4.898028, 5.071654, 
    5.245425, 5.419337, 5.593389, 5.76758, 5.941907, 6.116369, 6.290965, 
    6.465692, 6.640548, 6.815533, 6.990644, 7.165878, 7.341236, 7.516715, 
    7.692312, 7.868027, 8.043857, 8.2198, 8.395855, 8.57202, 8.748292, 
    8.92467, 9.101153, 9.277738, 9.454423, 9.631207, 9.808086, 9.985061, 
    10.16213, 10.33929, 10.51653, 10.69386, 10.87128, 11.04878, 11.22636, 
    11.40403, 11.58176, 11.75957, 11.93746, 12.11541, 12.29344, 12.47153, 
    12.64968, 12.8279, 13.00618, 13.18452, 13.36291, 13.54136, 13.71986, 
    13.89841, 14.07701, 14.25566, 14.43435, 14.61308, 14.79185, 14.97066, 
    15.1495, 15.32838, 15.50729, 15.68623, 15.8652, 16.04419, 16.22321, 
    16.40224, 16.5813, 16.76037, 16.93946, 17.11856, 17.29767, 17.47679, 
    17.65591, 17.83504, 18.01417, 18.1933, 18.37243, 18.55155, 18.73067, 
    18.90977, 19.08887, 19.26796, 19.44703, 19.62608, 19.80511, 19.98412, 
    20.16311, 20.34208, 20.52101, 20.69991, 20.87879, 21.05763, 21.23643, 
    21.4152, 21.59392, 21.77261, 21.95124, 22.12984, 22.30838, 22.48687, 
    22.66531, 22.8437, 23.02202, 23.20029, 23.3785, 23.55665, 23.73473, 
    23.91274, 24.09068, 24.26856, 24.44636, 24.62408, 24.80173, 24.9793, 
    25.15679, 25.33419, 25.51151, 25.68874, 25.86589, 26.04294, 26.2199, 
    26.39676, 26.57353, 26.7502, 26.92677, 27.10324, 27.2796, 27.45585, 
    27.632, 27.80804, 27.98396, 28.15978, 28.33547, 28.51105, 28.68651, 
    28.86185, 29.03707, 29.21216, 29.38712, 29.56196, 29.73666, 29.91124, 
    30.08568, 30.25998, 30.43415, 30.60818, 30.78207, 30.95582, 31.12942, 
    31.30288, 31.47619, 31.64936, 31.82237, 31.99523, 32.16794, 32.34049, 
    32.51288, 32.68512, 32.8572, 33.02911, 33.20086, 33.37245, 33.54387, 
    33.71513, 33.88621, 34.05713, 34.22787, 34.39844, 34.56883, 34.73905, 
    34.90909, 35.07895, 35.24863, 35.41813, 35.58744, 35.75657, 35.92551, 
    36.09427, 36.26284, 36.43122, 36.59941, 36.7674, 36.9352, 37.10281, 
    37.27022, 37.43743, 37.60444, 37.77126, 37.93787, 38.10428, 38.27048, 
    38.43649, 38.60228, 38.76787, 38.93325, 39.09843, 39.26339, 39.42814, 
    39.59268, 39.75701, 39.92112, 40.08502, 40.2487, 40.41216, 40.57541, 
    40.73844, 40.90125, 41.06383, 41.22619, 41.38833, 41.55025, 41.71194, 
    41.87341, 42.03465, 42.19566, 42.35645, 42.51701, 42.67733, 42.83743, 
    42.9973, 43.15693, 43.31633, 43.4755, 43.63444, 43.79314, 43.9516, 
    44.10983, 44.26782, 44.42558, 44.58309, 44.74037, 44.89741, 45.0542, 
    45.21076, 45.36708, 45.52316, 45.67899, 45.83458, 45.98992, 46.14502, 
    46.29988, 46.4545, 46.60886, 46.76299, 46.91687, 47.0705,
  -24.31235, -24.18202, -24.05146, -23.92064, -23.78958, -23.65826, -23.5267, 
    -23.3949, -23.26284, -23.13053, -22.99797, -22.86516, -22.73211, 
    -22.5988, -22.46524, -22.33143, -22.19736, -22.06305, -21.92848, 
    -21.79366, -21.65859, -21.52327, -21.38769, -21.25186, -21.11578, 
    -20.97944, -20.84285, -20.70601, -20.5689, -20.43155, -20.29394, 
    -20.15608, -20.01796, -19.87958, -19.74095, -19.60207, -19.46293, 
    -19.32353, -19.18388, -19.04397, -18.9038, -18.76338, -18.62271, 
    -18.48177, -18.34058, -18.19913, -18.05743, -17.91547, -17.77325, 
    -17.63077, -17.48804, -17.34505, -17.20181, -17.05831, -16.91455, 
    -16.77053, -16.62626, -16.48173, -16.33694, -16.1919, -16.0466, 
    -15.90104, -15.75523, -15.60916, -15.46283, -15.31625, -15.16941, 
    -15.02232, -14.87497, -14.72736, -14.5795, -14.43139, -14.28301, 
    -14.13439, -13.9855, -13.83637, -13.68698, -13.53733, -13.38743, 
    -13.23728, -13.08687, -12.93621, -12.7853, -12.63414, -12.48272, 
    -12.33105, -12.17913, -12.02696, -11.87454, -11.72186, -11.56894, 
    -11.41577, -11.26235, -11.10868, -10.95475, -10.80059, -10.64617, 
    -10.49151, -10.3366, -10.18144, -10.02604, -9.870393, -9.714501, 
    -9.558365, -9.401985, -9.245362, -9.088497, -8.93139, -8.774041, 
    -8.616451, -8.458621, -8.300552, -8.142244, -7.983697, -7.824914, 
    -7.665893, -7.506636, -7.347143, -7.187416, -7.027454, -6.86726, 
    -6.706832, -6.546174, -6.385283, -6.224164, -6.062814, -5.901236, 
    -5.73943, -5.577398, -5.41514, -5.252656, -5.089949, -4.927017, 
    -4.763864, -4.600489, -4.436894, -4.273079, -4.109046, -3.944795, 
    -3.780327, -3.615644, -3.450747, -3.285635, -3.120312, -2.954777, 
    -2.789032, -2.623078, -2.456915, -2.290546, -2.123971, -1.957191, 
    -1.790207, -1.623022, -1.455635, -1.288048, -1.120263, -0.9522797, 
    -0.7841005, -0.6157264, -0.4471585, -0.2783981, -0.1094467, 0.05969459, 
    0.2290244, 0.3985413, 0.568244, 0.7381312, 0.9082015, 1.078453, 1.248886, 
    1.419497, 1.590285, 1.76125, 1.932389, 2.103701, 2.275185, 2.446839, 
    2.618661, 2.790651, 2.962806, 3.135125, 3.307606, 3.480249, 3.653051, 
    3.82601, 3.999126, 4.172396, 4.345819, 4.519393, 4.693117, 4.866989, 
    5.041007, 5.21517, 5.389476, 5.563922, 5.738509, 5.913233, 6.088093, 
    6.263087, 6.438214, 6.613472, 6.788858, 6.964372, 7.14001, 7.315773, 
    7.491657, 7.667662, 7.843784, 8.020022, 8.196375, 8.37284, 8.549417, 
    8.726101, 8.902892, 9.079788, 9.256788, 9.433888, 9.611088, 9.788384, 
    9.965776, 10.14326, 10.32084, 10.4985, 10.67626, 10.8541, 11.03202, 
    11.21002, 11.38811, 11.56627, 11.7445, 11.92281, 12.10119, 12.27964, 
    12.45816, 12.63674, 12.81539, 12.9941, 13.17286, 13.35169, 13.53056, 
    13.70949, 13.88848, 14.0675, 14.24658, 14.4257, 14.60487, 14.78407, 
    14.96331, 15.14259, 15.3219, 15.50124, 15.68062, 15.86002, 16.03944, 
    16.21889, 16.39837, 16.57785, 16.75736, 16.93688, 17.11642, 17.29596, 
    17.47551, 17.65507, 17.83464, 18.0142, 18.19377, 18.37333, 18.55289, 
    18.73244, 18.91198, 19.09152, 19.27103, 19.45054, 19.63003, 19.80949, 
    19.98894, 20.16836, 20.34776, 20.52713, 20.70646, 20.88577, 21.06504, 
    21.24428, 21.42348, 21.60263, 21.78175, 21.96082, 22.13984, 22.31881, 
    22.49774, 22.67661, 22.85542, 23.03418, 23.21287, 23.39151, 23.57008, 
    23.74859, 23.92703, 24.1054, 24.2837, 24.46192, 24.64007, 24.81814, 
    24.99613, 25.17404, 25.35187, 25.5296, 25.70726, 25.88482, 26.06229, 
    26.23967, 26.41695, 26.59413, 26.77122, 26.9482, 27.12508, 27.30186, 
    27.47852, 27.65508, 27.83153, 28.00786, 28.18408, 28.36019, 28.53617, 
    28.71204, 28.88778, 29.0634, 29.23889, 29.41426, 29.5895, 29.7646, 
    29.93958, 30.11441, 30.28912, 30.46368, 30.63811, 30.81239, 30.98653, 
    31.16052, 31.33437, 31.50807, 31.68162, 31.85502, 32.02827, 32.20136, 
    32.37429, 32.54707, 32.71969, 32.89214, 33.06444, 33.23656, 33.40853, 
    33.58033, 33.75195, 33.92341, 34.09469, 34.2658, 34.43674, 34.6075, 
    34.77809, 34.94849, 35.11871, 35.28875, 35.45861, 35.62828, 35.79778, 
    35.96707, 36.13618, 36.30511, 36.47383, 36.64237, 36.81072, 36.97887, 
    37.14682, 37.31457, 37.48212, 37.64948, 37.81664, 37.98359, 38.15033, 
    38.31688, 38.48321, 38.64934, 38.81527, 38.98098, 39.14648, 39.31177, 
    39.47684, 39.64171, 39.80636, 39.97079, 40.13501, 40.29901, 40.46279, 
    40.62635, 40.78969, 40.9528, 41.1157, 41.27837, 41.44082, 41.60304, 
    41.76504, 41.92681, 42.08835, 42.24966, 42.41075, 42.5716, 42.73222, 
    42.89262, 43.05277, 43.2127, 43.37239, 43.53184, 43.69106, 43.85005, 
    44.00879, 44.1673, 44.32557, 44.4836, 44.6414, 44.79895, 44.95626, 
    45.11333, 45.27015, 45.42674, 45.58308, 45.73918, 45.89503, 46.05064, 
    46.206, 46.36112, 46.51599, 46.67061, 46.82499, 46.97912, 47.133,
  -24.39207, -24.26163, -24.13093, -23.99999, -23.8688, -23.73736, -23.60567, 
    -23.47374, -23.34155, -23.20911, -23.07642, -22.94348, -22.81028, 
    -22.67684, -22.54314, -22.40919, -22.27499, -22.14053, -22.00582, 
    -21.87086, -21.73565, -21.60017, -21.46445, -21.32847, -21.19224, 
    -21.05575, -20.919, -20.782, -20.64475, -20.50724, -20.36947, -20.23145, 
    -20.09317, -19.95463, -19.81584, -19.67679, -19.53748, -19.39792, 
    -19.25809, -19.11802, -18.97768, -18.83708, -18.69623, -18.55512, 
    -18.41376, -18.27213, -18.13025, -17.9881, -17.8457, -17.70304, 
    -17.56013, -17.41695, -17.27352, -17.12983, -16.98588, -16.84167, 
    -16.6972, -16.55248, -16.40749, -16.26225, -16.11675, -15.97099, 
    -15.82498, -15.6787, -15.53217, -15.38538, -15.23834, -15.09103, 
    -14.94347, -14.79565, -14.64758, -14.49924, -14.35065, -14.20181, 
    -14.0527, -13.90335, -13.75373, -13.60386, -13.45374, -13.30336, 
    -13.15272, -13.00183, -12.85068, -12.69928, -12.54763, -12.39573, 
    -12.24357, -12.09115, -11.93849, -11.78557, -11.6324, -11.47898, 
    -11.32531, -11.17139, -11.01722, -10.8628, -10.70813, -10.55321, 
    -10.39804, -10.24263, -10.08696, -9.931054, -9.774898, -9.618496, 
    -9.461849, -9.304957, -9.147821, -8.990442, -8.83282, -8.674954, 
    -8.516849, -8.3585, -8.199912, -8.041084, -7.882017, -7.722712, 
    -7.563168, -7.403388, -7.243371, -7.083118, -6.922631, -6.76191, 
    -6.600955, -6.439768, -6.278349, -6.116699, -5.954819, -5.79271, 
    -5.630373, -5.467807, -5.305016, -5.141998, -4.978755, -4.815289, 
    -4.6516, -4.487689, -4.323556, -4.159204, -3.994632, -3.829842, 
    -3.664835, -3.499613, -3.334175, -3.168523, -3.002658, -2.836582, 
    -2.670295, -2.503798, -2.337093, -2.17018, -2.003062, -1.835738, 
    -1.668211, -1.500481, -1.332549, -1.164418, -0.9960875, -0.8275594, 
    -0.6588348, -0.4899151, -0.3208015, -0.1514954, 0.01800188, 0.1876891, 
    0.3575649, 0.5276278, 0.6978766, 0.8683098, 1.038926, 1.209724, 1.380702, 
    1.551859, 1.723193, 1.894703, 2.066388, 2.238245, 2.410274, 2.582472, 
    2.754839, 2.927373, 3.100072, 3.272935, 3.44596, 3.619145, 3.79249, 
    3.965991, 4.139649, 4.31346, 4.487424, 4.661539, 4.835803, 5.010214, 
    5.184771, 5.359471, 5.534315, 5.709299, 5.884421, 6.05968, 6.235075, 
    6.410604, 6.586264, 6.762054, 6.937973, 7.114017, 7.290187, 7.466479, 
    7.642891, 7.819423, 7.996072, 8.172836, 8.349713, 8.526703, 8.703801, 
    8.881007, 9.058319, 9.235735, 9.413253, 9.590871, 9.768586, 9.946398, 
    10.1243, 10.3023, 10.48039, 10.65857, 10.83683, 11.01517, 11.1936, 
    11.37211, 11.5507, 11.72936, 11.9081, 12.0869, 12.26578, 12.44473, 
    12.62374, 12.80282, 12.98195, 13.16115, 13.3404, 13.51971, 13.69908, 
    13.87849, 14.05795, 14.23746, 14.41702, 14.59661, 14.77625, 14.95593, 
    15.13564, 15.31539, 15.49517, 15.67498, 15.85481, 16.03467, 16.21456, 
    16.39447, 16.57439, 16.75434, 16.93429, 17.11427, 17.29425, 17.47424, 
    17.65423, 17.83423, 18.01424, 18.19424, 18.37424, 18.55424, 18.73422, 
    18.9142, 19.09417, 19.27413, 19.45407, 19.63399, 19.8139, 19.99378, 
    20.17364, 20.35347, 20.53327, 20.71305, 20.89279, 21.0725, 21.25217, 
    21.4318, 21.61139, 21.79094, 21.97044, 22.14989, 22.3293, 22.50865, 
    22.68796, 22.8672, 23.04639, 23.22552, 23.40458, 23.58358, 23.76252, 
    23.94139, 24.12018, 24.29891, 24.47756, 24.65613, 24.83463, 25.01304, 
    25.19138, 25.36963, 25.54779, 25.72586, 25.90384, 26.08174, 26.25953, 
    26.43723, 26.61483, 26.79234, 26.96974, 27.14703, 27.32422, 27.5013, 
    27.67827, 27.85513, 28.03188, 28.20851, 28.38502, 28.56142, 28.73769, 
    28.91384, 29.08986, 29.26576, 29.44153, 29.61717, 29.79268, 29.96805, 
    30.14329, 30.31839, 30.49335, 30.66817, 30.84285, 31.01739, 31.19177, 
    31.36601, 31.5401, 31.71404, 31.88783, 32.06146, 32.23494, 32.40826, 
    32.58142, 32.75442, 32.92726, 33.09993, 33.27244, 33.44478, 33.61695, 
    33.78895, 33.96078, 34.13244, 34.30392, 34.47523, 34.64635, 34.81731, 
    34.98808, 35.15866, 35.32907, 35.49929, 35.66932, 35.83916, 36.00882, 
    36.17829, 36.34756, 36.51665, 36.68554, 36.85423, 37.02273, 37.19103, 
    37.35913, 37.52703, 37.69473, 37.86222, 38.02951, 38.1966, 38.36348, 
    38.53015, 38.69661, 38.86287, 39.02891, 39.19474, 39.36036, 39.52576, 
    39.69095, 39.85592, 40.02068, 40.18521, 40.34953, 40.51363, 40.67751, 
    40.84116, 41.00459, 41.1678, 41.33078, 41.49354, 41.65607, 41.81837, 
    41.98044, 42.14228, 42.3039, 42.46528, 42.62643, 42.78735, 42.94803, 
    43.10848, 43.2687, 43.42868, 43.58842, 43.74793, 43.9072, 44.06622, 
    44.22501, 44.38356, 44.54187, 44.69994, 44.85777, 45.01535, 45.1727, 
    45.32979, 45.48664, 45.64325, 45.79961, 45.95573, 46.1116, 46.26723, 
    46.4226, 46.57773, 46.73261, 46.88724, 47.04163, 47.19576,
  -24.47204, -24.34148, -24.21066, -24.0796, -23.94828, -23.81672, -23.6849, 
    -23.55283, -23.42051, -23.28794, -23.15512, -23.02205, -22.88872, 
    -22.75513, -22.6213, -22.48721, -22.35287, -22.21827, -22.08342, 
    -21.94831, -21.81295, -21.67734, -21.54146, -21.40534, -21.26895, 
    -21.13231, -20.99541, -20.85826, -20.72085, -20.58318, -20.44526, 
    -20.30708, -20.16864, -20.02994, -19.89098, -19.75177, -19.61229, 
    -19.47256, -19.33257, -19.19232, -19.05182, -18.91105, -18.77002, 
    -18.62874, -18.48719, -18.34539, -18.20333, -18.061, -17.91842, 
    -17.77558, -17.63247, -17.48911, -17.34549, -17.20161, -17.05747, 
    -16.91307, -16.76841, -16.62349, -16.47831, -16.33287, -16.18717, 
    -16.04121, -15.89499, -15.74851, -15.60177, -15.45478, -15.30752, 
    -15.16001, -15.01223, -14.8642, -14.71591, -14.56736, -14.41855, 
    -14.26949, -14.12017, -13.97058, -13.82075, -13.67065, -13.5203, 
    -13.36969, -13.21882, -13.0677, -12.91632, -12.76469, -12.6128, 
    -12.46066, -12.30826, -12.1556, -12.0027, -11.84954, -11.69612, 
    -11.54245, -11.38853, -11.23436, -11.07994, -10.92526, -10.77034, 
    -10.61516, -10.45974, -10.30406, -10.14814, -9.991964, -9.835544, 
    -9.678876, -9.521961, -9.364799, -9.207393, -9.049741, -8.891844, 
    -8.733704, -8.575319, -8.416693, -8.257824, -8.098714, -7.939363, 
    -7.779771, -7.619941, -7.459872, -7.299565, -7.139021, -6.97824, 
    -6.817224, -6.655972, -6.494487, -6.332768, -6.170817, -6.008635, 
    -5.846221, -5.683577, -5.520704, -5.357604, -5.194275, -5.03072, 
    -4.86694, -4.702935, -4.538707, -4.374256, -4.209583, -4.04469, 
    -3.879577, -3.714245, -3.548696, -3.382931, -3.216949, -3.050754, 
    -2.884345, -2.717724, -2.550892, -2.38385, -2.216599, -2.04914, 
    -1.881475, -1.713605, -1.545531, -1.377254, -1.208775, -1.040095, 
    -0.8712171, -0.7021408, -0.532868, -0.3633999, -0.1937378, -0.02388312, 
    0.1461629, 0.3163989, 0.4868234, 0.6574352, 0.8282328, 0.9992148, 
    1.17038, 1.341726, 1.513253, 1.684958, 1.856841, 2.028899, 2.201132, 
    2.373537, 2.546113, 2.718859, 2.891773, 3.064854, 3.238099, 3.411508, 
    3.585079, 3.75881, 3.932699, 4.106746, 4.280947, 4.455302, 4.629809, 
    4.804467, 4.979273, 5.154226, 5.329323, 5.504565, 5.679948, 5.855471, 
    6.031132, 6.206929, 6.382861, 6.558926, 6.735121, 6.911446, 7.087899, 
    7.264476, 7.441178, 7.618001, 7.794944, 7.972005, 8.149182, 8.326474, 
    8.503879, 8.681393, 8.859016, 9.036746, 9.21458, 9.392517, 9.570555, 
    9.748691, 9.926925, 10.10525, 10.28367, 10.46218, 10.64079, 10.81947, 
    10.99825, 11.1771, 11.35604, 11.53505, 11.71414, 11.89331, 12.07255, 
    12.25185, 12.43123, 12.61067, 12.79018, 12.96975, 13.14938, 13.32907, 
    13.50881, 13.68861, 13.86845, 14.04835, 14.2283, 14.40829, 14.58832, 
    14.76839, 14.94851, 15.12866, 15.30884, 15.48906, 15.6693, 15.84958, 
    16.02988, 16.2102, 16.39055, 16.57092, 16.7513, 16.93169, 17.1121, 
    17.29252, 17.47295, 17.65339, 17.83383, 18.01427, 18.19471, 18.37515, 
    18.55559, 18.73602, 18.91644, 19.09684, 19.27724, 19.45762, 19.63798, 
    19.81832, 19.99864, 20.17894, 20.35921, 20.53945, 20.71966, 20.89984, 
    21.07998, 21.26009, 21.44016, 21.62019, 21.80017, 21.98011, 22.16, 
    22.33984, 22.51963, 22.69936, 22.87904, 23.05866, 23.23822, 23.41772, 
    23.59715, 23.77652, 23.95581, 24.13504, 24.31419, 24.49327, 24.67227, 
    24.8512, 25.03004, 25.2088, 25.38747, 25.56606, 25.74456, 25.92296, 
    26.10128, 26.27949, 26.45761, 26.63564, 26.81356, 26.99137, 27.16909, 
    27.34669, 27.52419, 27.70158, 27.87885, 28.05601, 28.23305, 28.40998, 
    28.58678, 28.76346, 28.94002, 29.11645, 29.29276, 29.46893, 29.64498, 
    29.82089, 29.99666, 30.1723, 30.34781, 30.52316, 30.69838, 30.87346, 
    31.04839, 31.22317, 31.3978, 31.57229, 31.74662, 31.9208, 32.09482, 
    32.26868, 32.44239, 32.61593, 32.78931, 32.96254, 33.13559, 33.30848, 
    33.4812, 33.65375, 33.82613, 33.99833, 34.17036, 34.34221, 34.51389, 
    34.68539, 34.85671, 35.02784, 35.1988, 35.36956, 35.54015, 35.71054, 
    35.88075, 36.05077, 36.22059, 36.39022, 36.55966, 36.7289, 36.89795, 
    37.06679, 37.23544, 37.40388, 37.57213, 37.74017, 37.90801, 38.07564, 
    38.24307, 38.41029, 38.5773, 38.74409, 38.91068, 39.07706, 39.24322, 
    39.40917, 39.5749, 39.74041, 39.90571, 40.07079, 40.23565, 40.40028, 
    40.5647, 40.72889, 40.89286, 41.05661, 41.22013, 41.38342, 41.54648, 
    41.70932, 41.87193, 42.03431, 42.19645, 42.35836, 42.52005, 42.6815, 
    42.84271, 43.00369, 43.16443, 43.32494, 43.48521, 43.64524, 43.80503, 
    43.96458, 44.1239, 44.28297, 44.4418, 44.60039, 44.75874, 44.91684, 
    45.0747, 45.23231, 45.38968, 45.5468, 45.70367, 45.8603, 46.01669, 
    46.17282, 46.3287, 46.48434, 46.63972, 46.79486, 46.94975, 47.10438, 
    47.25877,
  -24.55227, -24.42159, -24.29065, -24.15946, -24.02802, -23.89633, 
    -23.76438, -23.63219, -23.49974, -23.36703, -23.23408, -23.10087, 
    -22.96741, -22.83369, -22.69972, -22.56549, -22.43101, -22.29627, 
    -22.16128, -22.02603, -21.89052, -21.75476, -21.61874, -21.48246, 
    -21.34593, -21.20914, -21.07209, -20.93478, -20.79722, -20.65939, 
    -20.52131, -20.38297, -20.24437, -20.10551, -19.96639, -19.82701, 
    -19.68737, -19.54747, -19.40731, -19.2669, -19.12621, -18.98528, 
    -18.84408, -18.70262, -18.56089, -18.41891, -18.27667, -18.13416, 
    -17.9914, -17.84837, -17.70509, -17.56154, -17.41773, -17.27366, 
    -17.12932, -16.98473, -16.83988, -16.69476, -16.54938, -16.40374, 
    -16.25784, -16.11168, -15.96526, -15.81858, -15.67164, -15.52443, 
    -15.37697, -15.22924, -15.08126, -14.93301, -14.78451, -14.63574, 
    -14.48672, -14.33743, -14.18789, -14.03808, -13.88802, -13.7377, 
    -13.58712, -13.43628, -13.28519, -13.13383, -12.98222, -12.83035, 
    -12.67823, -12.52584, -12.37321, -12.22031, -12.06716, -11.91376, 
    -11.7601, -11.60618, -11.45201, -11.29759, -11.14291, -10.98798, 
    -10.8328, -10.67737, -10.52169, -10.36575, -10.20956, -10.05313, 
    -9.896441, -9.739506, -9.582323, -9.424891, -9.267213, -9.109287, 
    -8.951116, -8.792699, -8.634037, -8.47513, -8.31598, -8.156587, 
    -7.996952, -7.837074, -7.676956, -7.516598, -7.356, -7.195163, -7.034088, 
    -6.872776, -6.711227, -6.549443, -6.387424, -6.225171, -6.062684, 
    -5.899965, -5.737014, -5.573833, -5.410422, -5.246782, -5.082914, 
    -4.918818, -4.754498, -4.589951, -4.42518, -4.260187, -4.094971, 
    -3.929533, -3.763876, -3.598, -3.431905, -3.265593, -3.099066, -2.932323, 
    -2.765367, -2.598199, -2.430818, -2.263228, -2.095428, -1.927421, 
    -1.759206, -1.590786, -1.422162, -1.253335, -1.084305, -0.9150753, 
    -0.7456461, -0.5760188, -0.4061949, -0.2361755, -0.06596201, 0.1044442, 
    0.2750418, 0.4458293, 0.6168055, 0.7879689, 0.9593181, 1.130852, 
    1.302568, 1.474466, 1.646544, 1.818801, 1.991234, 2.163843, 2.336627, 
    2.509582, 2.682709, 2.856005, 3.029469, 3.203098, 3.376893, 3.550851, 
    3.72497, 3.899248, 4.073685, 4.248279, 4.423027, 4.597928, 4.772981, 
    4.948183, 5.123534, 5.29903, 5.474671, 5.650455, 5.82638, 6.002444, 
    6.178646, 6.354983, 6.531455, 6.708057, 6.884791, 7.061653, 7.238641, 
    7.415753, 7.592989, 7.770346, 7.947821, 8.125414, 8.303122, 8.480943, 
    8.658875, 8.836916, 9.015065, 9.19332, 9.371678, 9.550138, 9.728698, 
    9.907354, 10.08611, 10.26495, 10.44389, 10.62292, 10.80203, 10.98123, 
    11.16052, 11.33988, 11.51933, 11.69885, 11.87844, 12.05811, 12.23785, 
    12.41766, 12.59754, 12.77748, 12.95749, 13.13755, 13.31767, 13.49785, 
    13.67808, 13.85837, 14.0387, 14.21909, 14.39951, 14.57999, 14.7605, 
    14.94105, 15.12164, 15.30226, 15.48292, 15.66361, 15.84432, 16.02506, 
    16.20583, 16.38661, 16.56742, 16.74824, 16.92908, 17.10993, 17.29079, 
    17.47166, 17.65254, 17.83342, 18.01431, 18.19519, 18.37607, 18.55695, 
    18.73782, 18.91868, 19.09953, 19.28036, 19.46118, 19.64199, 19.82277, 
    20.00353, 20.18427, 20.36498, 20.54566, 20.72631, 20.90693, 21.08751, 
    21.26806, 21.44856, 21.62903, 21.80945, 21.98983, 22.17015, 22.35043, 
    22.53065, 22.71082, 22.89094, 23.07099, 23.25099, 23.43092, 23.61078, 
    23.79058, 23.97031, 24.14997, 24.32956, 24.50907, 24.6885, 24.86785, 
    25.04712, 25.22631, 25.40541, 25.58442, 25.76334, 25.94217, 26.12091, 
    26.29955, 26.4781, 26.65654, 26.83488, 27.01312, 27.19125, 27.36928, 
    27.54719, 27.725, 27.90269, 28.08026, 28.25772, 28.43505, 28.61227, 
    28.78936, 28.96633, 29.14317, 29.31989, 29.49647, 29.67292, 29.84924, 
    30.02542, 30.20146, 30.37736, 30.55312, 30.72874, 30.90421, 31.07954, 
    31.25472, 31.42975, 31.60463, 31.77935, 31.95392, 32.12833, 32.30259, 
    32.47668, 32.65061, 32.82438, 32.99798, 33.17142, 33.34469, 33.51779, 
    33.69072, 33.86347, 34.03605, 34.20846, 34.38069, 34.55274, 34.72461, 
    34.89629, 35.0678, 35.23912, 35.41025, 35.5812, 35.75196, 35.92252, 
    36.0929, 36.26308, 36.43307, 36.60286, 36.77246, 36.94186, 37.11106, 
    37.28005, 37.44885, 37.61744, 37.78583, 37.95401, 38.12199, 38.28975, 
    38.45731, 38.62466, 38.79179, 38.95871, 39.12542, 39.29192, 39.45819, 
    39.62425, 39.7901, 39.95572, 40.12112, 40.2863, 40.45126, 40.61599, 
    40.78051, 40.94479, 41.10885, 41.27268, 41.43629, 41.59966, 41.76281, 
    41.92572, 42.0884, 42.25085, 42.41307, 42.57505, 42.7368, 42.89831, 
    43.05958, 43.22062, 43.38142, 43.54198, 43.7023, 43.86238, 44.02222, 
    44.18182, 44.34117, 44.50028, 44.65915, 44.81778, 44.97615, 45.13428, 
    45.29217, 45.44981, 45.6072, 45.76435, 45.92124, 46.07789, 46.23429, 
    46.39043, 46.54633, 46.70197, 46.85737, 47.01251, 47.1674, 47.32203,
  -24.63276, -24.50195, -24.37089, -24.23958, -24.10801, -23.97619, 
    -23.84412, -23.7118, -23.57922, -23.44638, -23.3133, -23.17995, 
    -23.04636, -22.9125, -22.77839, -22.64403, -22.50941, -22.37453, 
    -22.2394, -22.104, -21.96835, -21.83244, -21.69628, -21.55985, -21.42317, 
    -21.28623, -21.14902, -21.01156, -20.87384, -20.73586, -20.59762, 
    -20.45912, -20.32036, -20.18134, -20.04206, -19.90252, -19.76271, 
    -19.62265, -19.48232, -19.34173, -19.20088, -19.05977, -18.9184, 
    -18.77676, -18.63486, -18.4927, -18.35028, -18.20759, -18.06465, 
    -17.92144, -17.77796, -17.63423, -17.49023, -17.34597, -17.20144, 
    -17.05666, -16.91161, -16.7663, -16.62073, -16.47489, -16.32879, 
    -16.18243, -16.0358, -15.88892, -15.74177, -15.59436, -15.44668, 
    -15.29875, -15.15055, -15.00209, -14.85337, -14.70439, -14.55514, 
    -14.40564, -14.25587, -14.10585, -13.95556, -13.80501, -13.65421, 
    -13.50314, -13.35181, -13.20023, -13.04838, -12.89628, -12.74391, 
    -12.59129, -12.43841, -12.28528, -12.13189, -11.97824, -11.82433, 
    -11.67017, -11.51575, -11.36107, -11.20614, -11.05096, -10.89552, 
    -10.73983, -10.58389, -10.42769, -10.27124, -10.11454, -9.957591, 
    -9.800388, -9.642937, -9.485234, -9.327284, -9.169085, -9.010637, 
    -8.851943, -8.693002, -8.533815, -8.374383, -8.214706, -8.054786, 
    -7.894622, -7.734215, -7.573567, -7.412677, -7.251547, -7.090177, 
    -6.928569, -6.766722, -6.604638, -6.442317, -6.279761, -6.11697, 
    -5.953944, -5.790686, -5.627195, -5.463473, -5.29952, -5.135338, 
    -4.970927, -4.806288, -4.641423, -4.476332, -4.311016, -4.145476, 
    -3.979713, -3.813729, -3.647524, -3.4811, -3.314456, -3.147596, 
    -2.980519, -2.813226, -2.64572, -2.478, -2.310069, -2.141927, -1.973576, 
    -1.805016, -1.636249, -1.467276, -1.298099, -1.128718, -0.9591358, 
    -0.7893522, -0.6193693, -0.4491881, -0.27881, -0.1082364, 0.06253137, 
    0.2334919, 0.4046439, 0.575986, 0.7475166, 0.9192345, 1.091138, 1.263226, 
    1.435497, 1.607949, 1.780581, 1.953391, 2.126379, 2.299541, 2.472878, 
    2.646387, 2.820066, 2.993914, 3.16793, 3.342112, 3.516459, 3.690967, 
    3.865637, 4.040466, 4.215453, 4.390596, 4.565893, 4.741343, 4.916944, 
    5.092693, 5.26859, 5.444633, 5.62082, 5.797149, 5.973618, 6.150226, 
    6.32697, 6.50385, 6.680861, 6.858005, 7.035278, 7.212678, 7.390205, 
    7.567854, 7.745626, 7.923518, 8.101527, 8.279654, 8.457893, 8.636246, 
    8.814708, 8.993279, 9.171956, 9.350738, 9.529621, 9.708605, 9.887688, 
    10.06687, 10.24614, 10.42551, 10.60496, 10.78451, 10.96414, 11.14385, 
    11.32365, 11.50352, 11.68348, 11.86351, 12.04361, 12.22379, 12.40403, 
    12.58434, 12.76472, 12.94516, 13.12566, 13.30622, 13.48684, 13.66751, 
    13.84823, 14.02901, 14.20983, 14.3907, 14.57161, 14.75256, 14.93356, 
    15.11459, 15.29565, 15.47675, 15.65788, 15.83904, 16.02022, 16.20143, 
    16.38266, 16.5639, 16.74517, 16.92645, 17.10775, 17.28905, 17.47037, 
    17.65169, 17.83301, 18.01434, 18.19567, 18.37699, 18.55831, 18.73963, 
    18.92093, 19.10222, 19.2835, 19.46477, 19.64601, 19.82724, 20.00844, 
    20.18962, 20.37078, 20.5519, 20.73299, 20.91405, 21.09508, 21.27606, 
    21.45701, 21.63791, 21.81878, 21.99959, 22.18036, 22.36107, 22.54174, 
    22.72235, 22.90289, 23.08339, 23.26382, 23.44419, 23.62449, 23.80472, 
    23.98488, 24.16498, 24.34499, 24.52494, 24.7048, 24.88458, 25.06429, 
    25.2439, 25.42343, 25.60287, 25.78222, 25.96148, 26.14065, 26.31971, 
    26.49868, 26.67755, 26.85632, 27.03498, 27.21353, 27.39197, 27.57031, 
    27.74853, 27.92664, 28.10463, 28.2825, 28.46025, 28.63789, 28.81539, 
    28.99277, 29.17002, 29.34715, 29.52414, 29.701, 29.87772, 30.05431, 
    30.23075, 30.40706, 30.58322, 30.75924, 30.93512, 31.11084, 31.28642, 
    31.46185, 31.63712, 31.81224, 31.9872, 32.162, 32.33665, 32.51113, 
    32.68545, 32.85961, 33.0336, 33.20742, 33.38107, 33.55455, 33.72786, 
    33.901, 34.07396, 34.24674, 34.41934, 34.59177, 34.76401, 34.93607, 
    35.10794, 35.27963, 35.45113, 35.62244, 35.79356, 35.96449, 36.13523, 
    36.30577, 36.47612, 36.64627, 36.81622, 36.98597, 37.15553, 37.32487, 
    37.49402, 37.66296, 37.83169, 38.00022, 38.16854, 38.33665, 38.50454, 
    38.67223, 38.8397, 39.00696, 39.174, 39.34083, 39.50744, 39.67383, 39.84, 
    40.00595, 40.17168, 40.33718, 40.50246, 40.66752, 40.83235, 40.99695, 
    41.16132, 41.32547, 41.48939, 41.65307, 41.81652, 41.97975, 42.14273, 
    42.30549, 42.46801, 42.63029, 42.79234, 42.95415, 43.11572, 43.27705, 
    43.43814, 43.599, 43.75961, 43.91998, 44.0801, 44.23998, 44.39962, 
    44.55901, 44.71816, 44.87706, 45.03572, 45.19413, 45.35229, 45.5102, 
    45.66786, 45.82527, 45.98243, 46.13935, 46.29601, 46.45242, 46.60857, 
    46.76448, 46.92013, 47.07553, 47.23067, 47.38556,
  -24.7135, -24.58257, -24.45139, -24.31995, -24.18826, -24.05632, -23.92412, 
    -23.79167, -23.65896, -23.526, -23.39278, -23.2593, -23.12557, -22.99158, 
    -22.85733, -22.72283, -22.58807, -22.45305, -22.31778, -22.18224, 
    -22.04645, -21.91039, -21.77408, -21.63751, -21.50067, -21.36358, 
    -21.22623, -21.08861, -20.95074, -20.8126, -20.6742, -20.53555, 
    -20.39663, -20.25744, -20.118, -19.97829, -19.83832, -19.69809, 
    -19.55759, -19.41684, -19.27581, -19.13453, -18.99298, -18.85117, 
    -18.7091, -18.56676, -18.42416, -18.28129, -18.13816, -17.99477, 
    -17.85111, -17.70719, -17.563, -17.41855, -17.27383, -17.12886, 
    -16.98361, -16.83811, -16.69234, -16.5463, -16.4, -16.25344, -16.10661, 
    -15.95952, -15.81216, -15.66455, -15.51666, -15.36852, -15.22011, 
    -15.07143, -14.9225, -14.7733, -14.62384, -14.47411, -14.32413, 
    -14.17388, -14.02337, -13.87259, -13.72156, -13.57026, -13.4187, 
    -13.26688, -13.1148, -12.96246, -12.80986, -12.65701, -12.50389, 
    -12.35051, -12.19687, -12.04298, -11.88882, -11.73441, -11.57974, 
    -11.42482, -11.26963, -11.1142, -10.9585, -10.80255, -10.64635, 
    -10.48989, -10.33318, -10.17621, -10.019, -9.861526, -9.703804, 
    -9.545831, -9.387607, -9.229134, -9.07041, -8.911438, -8.752218, 
    -8.59275, -8.433035, -8.273074, -8.112867, -7.952416, -7.79172, 
    -7.630781, -7.469599, -7.308175, -7.146509, -6.984603, -6.822457, 
    -6.660072, -6.497449, -6.334589, -6.171493, -6.00816, -5.844593, 
    -5.680792, -5.516758, -5.352491, -5.187994, -5.023266, -4.858309, 
    -4.693124, -4.527711, -4.362072, -4.196208, -4.030118, -3.863806, 
    -3.697272, -3.530516, -3.36354, -3.196345, -3.028933, -2.861303, 
    -2.693458, -2.525398, -2.357124, -2.188639, -2.019942, -1.851036, 
    -1.681921, -1.512599, -1.34307, -1.173337, -1.0034, -0.833261, 
    -0.6629209, -0.4923811, -0.321643, -0.1507079, 0.0204228, 0.1917478, 
    0.3632656, 0.5349749, 0.7068742, 0.8789622, 1.051237, 1.223698, 1.396343, 
    1.569171, 1.74218, 1.915369, 2.088736, 2.26228, 2.435999, 2.609891, 
    2.783956, 2.95819, 3.132594, 3.307165, 3.481901, 3.656801, 3.831864, 
    4.007087, 4.182469, 4.358008, 4.533703, 4.709552, 4.885552, 5.061703, 
    5.238003, 5.414449, 5.59104, 5.767775, 5.944651, 6.121666, 6.29882, 
    6.476109, 6.653533, 6.831089, 7.008775, 7.186589, 7.364531, 7.542596, 
    7.720785, 7.899095, 8.077524, 8.256069, 8.434731, 8.613504, 8.79239, 
    8.971384, 9.150485, 9.329692, 9.509002, 9.688413, 9.867924, 10.04753, 
    10.22723, 10.40703, 10.58692, 10.76689, 10.94695, 11.1271, 11.30733, 
    11.48764, 11.66803, 11.84849, 12.02903, 12.20965, 12.39033, 12.57108, 
    12.75189, 12.93277, 13.11371, 13.29471, 13.47577, 13.65688, 13.83805, 
    14.01926, 14.20053, 14.38184, 14.56319, 14.74459, 14.92602, 15.1075, 
    15.28901, 15.47055, 15.65212, 15.83372, 16.01535, 16.197, 16.37868, 
    16.56037, 16.74208, 16.92381, 17.10555, 17.28731, 17.46906, 17.65083, 
    17.8326, 18.01438, 18.19615, 18.37792, 18.55969, 18.74145, 18.92319, 
    19.10493, 19.28666, 19.46837, 19.65006, 19.83173, 20.01338, 20.19501, 
    20.3766, 20.55817, 20.73971, 20.92121, 21.10268, 21.28411, 21.4655, 
    21.64685, 21.82815, 22.00941, 22.19061, 22.37177, 22.55287, 22.73392, 
    22.91491, 23.09584, 23.27671, 23.45752, 23.63826, 23.81893, 23.99953, 
    24.18006, 24.36051, 24.54089, 24.72119, 24.9014, 25.08154, 25.26158, 
    25.44155, 25.62142, 25.8012, 25.98089, 26.16048, 26.33997, 26.51937, 
    26.69866, 26.87785, 27.05694, 27.23591, 27.41478, 27.59354, 27.77218, 
    27.95071, 28.12912, 28.30741, 28.48558, 28.66363, 28.84155, 29.01934, 
    29.19701, 29.37454, 29.55194, 29.72921, 29.90634, 30.08334, 30.26019, 
    30.4369, 30.61347, 30.78989, 30.96617, 31.1423, 31.31828, 31.4941, 
    31.66977, 31.84528, 32.02064, 32.19584, 32.37088, 32.54575, 32.72046, 
    32.895, 33.06938, 33.24359, 33.41763, 33.59149, 33.76518, 33.9387, 
    34.11204, 34.2852, 34.45818, 34.63098, 34.8036, 34.97602, 35.14827, 
    35.32033, 35.4922, 35.66388, 35.83537, 36.00666, 36.17776, 36.34866, 
    36.51937, 36.68988, 36.86019, 37.0303, 37.2002, 37.3699, 37.5394, 
    37.70869, 37.87777, 38.04664, 38.21531, 38.38375, 38.55199, 38.72002, 
    38.88783, 39.05543, 39.22281, 39.38997, 39.55691, 39.72363, 39.89013, 
    40.05641, 40.22246, 40.38829, 40.55389, 40.71927, 40.88442, 41.04934, 
    41.21403, 41.37849, 41.54272, 41.70672, 41.87048, 42.03401, 42.19731, 
    42.36037, 42.52319, 42.68578, 42.84812, 43.01023, 43.1721, 43.33372, 
    43.49511, 43.65625, 43.81716, 43.97781, 44.13823, 44.29839, 44.45832, 
    44.61799, 44.77742, 44.9366, 45.09554, 45.25422, 45.41265, 45.57084, 
    45.72877, 45.88645, 46.04388, 46.20106, 46.35799, 46.51466, 46.67107, 
    46.82724, 46.98315, 47.1388, 47.2942, 47.44934,
  -24.7945, -24.66345, -24.53214, -24.40059, -24.26877, -24.1367, -24.00438, 
    -23.8718, -23.73896, -23.60587, -23.47252, -23.33891, -23.20504, 
    -23.07092, -22.93654, -22.8019, -22.667, -22.53184, -22.39642, -22.26074, 
    -22.1248, -21.98861, -21.85215, -21.71543, -21.57844, -21.4412, 
    -21.30369, -21.16593, -21.0279, -20.88961, -20.75105, -20.61223, 
    -20.47315, -20.33381, -20.1942, -20.05433, -19.9142, -19.7738, -19.63313, 
    -19.49221, -19.35102, -19.20956, -19.06784, -18.92585, -18.7836, 
    -18.64108, -18.4983, -18.35526, -18.21194, -18.06837, -17.92452, 
    -17.78041, -17.63604, -17.4914, -17.34649, -17.20132, -17.05589, 
    -16.91018, -16.76422, -16.61798, -16.47148, -16.32472, -16.17769, 
    -16.03039, -15.88283, -15.735, -15.58691, -15.43855, -15.28993, 
    -15.14105, -14.99189, -14.84248, -14.6928, -14.54285, -14.39264, 
    -14.24217, -14.09144, -13.94044, -13.78917, -13.63765, -13.48586, 
    -13.33381, -13.18149, -13.02892, -12.87608, -12.72298, -12.56962, 
    -12.416, -12.26212, -12.10798, -11.95358, -11.79892, -11.644, -11.48882, 
    -11.33338, -11.17769, -11.02174, -10.86553, -10.70907, -10.55235, 
    -10.39537, -10.23814, -10.08066, -9.922919, -9.764927, -9.606682, 
    -9.448185, -9.289436, -9.130436, -8.971186, -8.811686, -8.651936, 
    -8.491938, -8.331692, -8.171199, -8.010459, -7.849473, -7.688242, 
    -7.526767, -7.365047, -7.203085, -7.040882, -6.878436, -6.71575, 
    -6.552824, -6.389658, -6.226255, -6.062615, -5.898738, -5.734626, 
    -5.570279, -5.405698, -5.240884, -5.075839, -4.910563, -4.745056, 
    -4.579321, -4.413358, -4.247167, -4.080751, -3.91411, -3.747245, 
    -3.580157, -3.412847, -3.245317, -3.077567, -2.909599, -2.741413, 
    -2.573012, -2.404395, -2.235565, -2.066522, -1.897268, -1.727804, 
    -1.55813, -1.38825, -1.218162, -1.04787, -0.877374, -0.7066754, 
    -0.5357757, -0.3646762, -0.1933782, -0.02188314, 0.1498076, 0.3216927, 
    0.4937707, 0.6660402, 0.8384997, 1.011148, 1.183983, 1.357004, 1.530209, 
    1.703597, 1.877165, 2.050914, 2.22484, 2.398943, 2.573221, 2.747672, 
    2.922295, 3.097088, 3.272049, 3.447177, 3.622471, 3.797928, 3.973547, 
    4.149326, 4.325263, 4.501357, 4.677606, 4.854009, 5.030562, 5.207266, 
    5.384118, 5.561115, 5.738257, 5.915542, 6.092968, 6.270532, 6.448233, 
    6.62607, 6.804039, 6.982141, 7.160371, 7.338729, 7.517214, 7.695822, 
    7.874551, 8.053401, 8.232369, 8.411452, 8.590651, 8.76996, 8.94938, 
    9.128908, 9.308542, 9.48828, 9.66812, 9.848061, 10.0281, 10.20823, 
    10.38846, 10.56878, 10.74919, 10.92968, 11.11027, 11.29093, 11.47168, 
    11.6525, 11.83341, 12.01439, 12.19544, 12.37656, 12.55775, 12.739, 
    12.92032, 13.1017, 13.28315, 13.46465, 13.6462, 13.82781, 14.00947, 
    14.19118, 14.37293, 14.55473, 14.73657, 14.91845, 15.10037, 15.28233, 
    15.46432, 15.64634, 15.82838, 16.01046, 16.19256, 16.37468, 16.55682, 
    16.73898, 16.92116, 17.10335, 17.28555, 17.46776, 17.64997, 17.83219, 
    18.01441, 18.19663, 18.37885, 18.56107, 18.74327, 18.92547, 19.10766, 
    19.28983, 19.47199, 19.65413, 19.83625, 20.01834, 20.20041, 20.38246, 
    20.56447, 20.74646, 20.92841, 21.11032, 21.2922, 21.47403, 21.65582, 
    21.83757, 22.01927, 22.20092, 22.38252, 22.56407, 22.74556, 22.92699, 
    23.10836, 23.28967, 23.47092, 23.6521, 23.83321, 24.01425, 24.19521, 
    24.3761, 24.55692, 24.73765, 24.9183, 25.09887, 25.27936, 25.45975, 
    25.64005, 25.82027, 26.00039, 26.18041, 26.36033, 26.54016, 26.71988, 
    26.8995, 27.07901, 27.25841, 27.4377, 27.61688, 27.79595, 27.9749, 
    28.15373, 28.33244, 28.51103, 28.68949, 28.86783, 29.04604, 29.22412, 
    29.40207, 29.57989, 29.75756, 29.93511, 30.11251, 30.28977, 30.46689, 
    30.64387, 30.8207, 30.99738, 31.17391, 31.35028, 31.52651, 31.70258, 
    31.87849, 32.05424, 32.22984, 32.40527, 32.58054, 32.75564, 32.93057, 
    33.10534, 33.27993, 33.45436, 33.62861, 33.80268, 33.97658, 34.1503, 
    34.32384, 34.4972, 34.67038, 34.84337, 35.01617, 35.18879, 35.36122, 
    35.53346, 35.70551, 35.87737, 36.04902, 36.22049, 36.39175, 36.56282, 
    36.73369, 36.90436, 37.07482, 37.24508, 37.41513, 37.58498, 37.75462, 
    37.92406, 38.09328, 38.26229, 38.43108, 38.59966, 38.76803, 38.93618, 
    39.10412, 39.27183, 39.43933, 39.6066, 39.77365, 39.94048, 40.10709, 
    40.27347, 40.43962, 40.60555, 40.77125, 40.93672, 41.10196, 41.26697, 
    41.43175, 41.59629, 41.7606, 41.92467, 42.08852, 42.25212, 42.41549, 
    42.57861, 42.7415, 42.90415, 43.06656, 43.22872, 43.39064, 43.55233, 
    43.71376, 43.87495, 44.0359, 44.1966, 44.35706, 44.51727, 44.67722, 
    44.83693, 44.99639, 45.15561, 45.31456, 45.47327, 45.63173, 45.78994, 
    45.94789, 46.10559, 46.26303, 46.42022, 46.57716, 46.73384, 46.89026, 
    47.04642, 47.20234, 47.35799, 47.51339,
  -24.87576, -24.74459, -24.61316, -24.48148, -24.34954, -24.21735, -24.0849, 
    -23.95219, -23.81923, -23.686, -23.55252, -23.41878, -23.28478, 
    -23.15052, -23.016, -22.88123, -22.74619, -22.61089, -22.47533, 
    -22.33951, -22.20343, -22.06709, -21.93048, -21.79361, -21.65648, 
    -21.51909, -21.38143, -21.24351, -21.10533, -20.96688, -20.82817, 
    -20.68919, -20.54995, -20.41045, -20.27068, -20.13064, -19.99034, 
    -19.84978, -19.70895, -19.56785, -19.42649, -19.28486, -19.14296, 
    -19.0008, -18.85837, -18.71568, -18.57272, -18.42949, -18.286, -18.14223, 
    -17.99821, -17.85391, -17.70935, -17.56452, -17.41942, -17.27406, 
    -17.12843, -16.98253, -16.83636, -16.68993, -16.54323, -16.39627, 
    -16.24903, -16.10153, -15.95376, -15.80573, -15.65743, -15.50886, 
    -15.36003, -15.21093, -15.06156, -14.91193, -14.76203, -14.61186, 
    -14.46143, -14.31074, -14.15978, -14.00855, -13.85706, -13.7053, 
    -13.55328, -13.401, -13.24845, -13.09564, -12.94256, -12.78922, 
    -12.63562, -12.48176, -12.32763, -12.17325, -12.0186, -11.86369, 
    -11.70852, -11.55309, -11.3974, -11.24145, -11.08524, -10.92877, 
    -10.77205, -10.61507, -10.45783, -10.30033, -10.14258, -9.984571, 
    -9.826307, -9.66779, -9.509019, -9.349995, -9.190717, -9.031188, 
    -8.871407, -8.711375, -8.551093, -8.390561, -8.22978, -8.068751, 
    -7.907475, -7.745952, -7.584183, -7.422168, -7.259909, -7.097405, 
    -6.934659, -6.771671, -6.608441, -6.444971, -6.28126, -6.117311, 
    -5.953124, -5.788699, -5.624038, -5.459142, -5.294011, -5.128647, 
    -4.96305, -4.797222, -4.631163, -4.464874, -4.298357, -4.131612, 
    -3.964641, -3.797444, -3.630023, -3.462378, -3.294511, -3.126423, 
    -2.958116, -2.789589, -2.620844, -2.451884, -2.282707, -2.113317, 
    -1.943714, -1.773899, -1.603873, -1.433639, -1.263196, -1.092547, 
    -0.9216929, -0.7506346, -0.5793735, -0.4079112, -0.236249, -0.06438813, 
    0.1076699, 0.2799237, 0.4523718, 0.6250129, 0.7978455, 0.9708681, 
    1.144079, 1.317477, 1.491061, 1.664829, 1.838779, 2.012911, 2.187221, 
    2.36171, 2.536375, 2.711214, 2.886226, 3.06141, 3.236764, 3.412286, 
    3.587974, 3.763827, 3.939843, 4.116021, 4.292358, 4.468853, 4.645505, 
    4.822311, 4.999269, 5.176379, 5.353638, 5.531044, 5.708595, 5.88629, 
    6.064127, 6.242104, 6.420219, 6.598471, 6.776856, 6.955375, 7.134023, 
    7.312801, 7.491705, 7.670734, 7.849886, 8.029159, 8.20855, 8.388059, 
    8.567683, 8.747419, 8.927267, 9.107224, 9.287287, 9.467455, 9.647726, 
    9.828098, 10.00857, 10.18914, 10.3698, 10.55055, 10.7314, 10.91233, 
    11.09335, 11.27445, 11.45564, 11.6369, 11.81824, 11.99966, 12.18115, 
    12.36272, 12.54435, 12.72605, 12.90781, 13.08963, 13.27152, 13.45346, 
    13.63546, 13.81752, 13.99962, 14.18178, 14.36398, 14.54623, 14.72851, 
    14.91084, 15.09321, 15.27562, 15.45805, 15.64052, 15.82302, 16.00554, 
    16.18809, 16.37066, 16.55326, 16.73587, 16.91849, 17.10113, 17.28378, 
    17.46644, 17.64911, 17.83178, 18.01445, 18.19712, 18.37979, 18.56245, 
    18.74511, 18.92776, 19.1104, 19.29302, 19.47563, 19.65822, 19.84079, 
    20.02333, 20.20585, 20.38834, 20.57081, 20.75324, 20.93564, 21.118, 
    21.30032, 21.4826, 21.66484, 21.84704, 22.02919, 22.21128, 22.39333, 
    22.57532, 22.75726, 22.93913, 23.12095, 23.3027, 23.48439, 23.66601, 
    23.84756, 24.02904, 24.21045, 24.39178, 24.57303, 24.7542, 24.93529, 
    25.1163, 25.29722, 25.47805, 25.65879, 25.83943, 26.01999, 26.20044, 
    26.3808, 26.56105, 26.7412, 26.92125, 27.10119, 27.28102, 27.46074, 
    27.64034, 27.81983, 27.99921, 28.17846, 28.35759, 28.5366, 28.71549, 
    28.89425, 29.07287, 29.25137, 29.42974, 29.60797, 29.78606, 29.96401, 
    30.14183, 30.3195, 30.49703, 30.67441, 30.85165, 31.02873, 31.20567, 
    31.38245, 31.55908, 31.73555, 31.91186, 32.08801, 32.264, 32.43983, 
    32.61549, 32.79099, 32.96631, 33.14147, 33.31646, 33.49127, 33.6659, 
    33.84036, 34.01464, 34.18875, 34.36267, 34.53641, 34.70996, 34.88333, 
    35.05651, 35.22951, 35.40231, 35.57492, 35.74734, 35.91956, 36.09159, 
    36.26342, 36.43505, 36.60648, 36.77771, 36.94873, 37.11956, 37.29017, 
    37.46058, 37.63078, 37.80077, 37.97056, 38.14013, 38.30948, 38.47863, 
    38.64755, 38.81626, 38.98475, 39.15303, 39.32108, 39.48891, 39.65652, 
    39.82391, 39.99107, 40.158, 40.32471, 40.49119, 40.65744, 40.82347, 
    40.98926, 41.15482, 41.32015, 41.48524, 41.6501, 41.81472, 41.97911, 
    42.14326, 42.30717, 42.47084, 42.63428, 42.79747, 42.96042, 43.12313, 
    43.28559, 43.44781, 43.60979, 43.77152, 43.933, 44.09424, 44.25523, 
    44.41597, 44.57646, 44.73671, 44.8967, 45.05644, 45.21593, 45.37517, 
    45.53415, 45.69288, 45.85136, 46.00958, 46.16755, 46.32526, 46.48272, 
    46.63992, 46.79686, 46.95354, 47.10997, 47.26614, 47.42204, 47.57769,
  -24.95728, -24.82599, -24.69444, -24.56264, -24.43058, -24.29826, 
    -24.16568, -24.03285, -23.89975, -23.7664, -23.63279, -23.49892, 
    -23.36478, -23.23039, -23.09574, -22.96082, -22.82565, -22.69021, 
    -22.55451, -22.41855, -22.28232, -22.14583, -22.00908, -21.87207, 
    -21.73479, -21.59724, -21.45943, -21.32136, -21.18303, -21.04442, 
    -20.90555, -20.76642, -20.62702, -20.48736, -20.34742, -20.20723, 
    -20.06676, -19.92603, -19.78503, -19.64376, -19.50223, -19.36043, 
    -19.21836, -19.07603, -18.93342, -18.79055, -18.64741, -18.504, 
    -18.36032, -18.21638, -18.07217, -17.92768, -17.78293, -17.63791, 
    -17.49263, -17.34707, -17.20124, -17.05515, -16.90879, -16.76216, 
    -16.61526, -16.46809, -16.32065, -16.17295, -16.02497, -15.87673, 
    -15.72822, -15.57944, -15.4304, -15.28108, -15.1315, -14.98165, 
    -14.83153, -14.68114, -14.53049, -14.37957, -14.22839, -14.07693, 
    -13.92521, -13.77323, -13.62097, -13.46846, -13.31567, -13.16263, 
    -13.00931, -12.85573, -12.70189, -12.54778, -12.39341, -12.23878, 
    -12.08388, -11.92873, -11.7733, -11.61762, -11.46168, -11.30547, -11.149, 
    -10.99228, -10.83529, -10.67805, -10.52054, -10.36278, -10.20476, 
    -10.04648, -9.887948, -9.729157, -9.570111, -9.41081, -9.251255, 
    -9.091446, -8.931384, -8.77107, -8.610502, -8.449684, -8.288616, 
    -8.127297, -7.965729, -7.803913, -7.641849, -7.479538, -7.31698, 
    -7.154178, -6.99113, -6.827838, -6.664303, -6.500526, -6.336508, 
    -6.172249, -6.00775, -5.843012, -5.678037, -5.512824, -5.347375, 
    -5.181692, -5.015773, -4.849622, -4.683239, -4.516623, -4.349778, 
    -4.182704, -4.015401, -3.847872, -3.680116, -3.512136, -3.343931, 
    -3.175504, -3.006855, -2.837986, -2.668898, -2.499591, -2.330068, 
    -2.160329, -1.990375, -1.820208, -1.649829, -1.47924, -1.308441, 
    -1.137434, -0.9662195, -0.7948, -0.6231763, -0.4513498, -0.2793218, 
    -0.1070938, 0.06533285, 0.2379568, 0.4107766, 0.5837908, 0.7569979, 
    0.9303964, 1.103985, 1.277762, 1.451726, 1.625876, 1.800209, 1.974725, 
    2.149421, 2.324297, 2.499351, 2.67458, 2.849984, 3.02556, 3.201308, 
    3.377225, 3.55331, 3.729561, 3.905976, 4.082554, 4.259293, 4.436191, 
    4.613246, 4.790458, 4.967823, 5.14534, 5.323008, 5.500823, 5.678786, 
    5.856894, 6.035144, 6.213536, 6.392067, 6.570735, 6.749539, 6.928476, 
    7.107545, 7.286743, 7.46607, 7.645522, 7.825098, 8.004795, 8.184613, 
    8.364549, 8.5446, 8.724766, 8.905043, 9.085429, 9.265924, 9.446525, 
    9.627229, 9.808035, 9.98894, 10.16994, 10.35104, 10.53223, 10.71352, 
    10.89489, 11.07634, 11.25789, 11.43951, 11.62122, 11.803, 11.98486, 
    12.1668, 12.34881, 12.53088, 12.71302, 12.89523, 13.0775, 13.25984, 
    13.44223, 13.62467, 13.80718, 13.98973, 14.17233, 14.35498, 14.53768, 
    14.72042, 14.9032, 15.08601, 15.26887, 15.45176, 15.63468, 15.81763, 
    16.0006, 16.1836, 16.36663, 16.54967, 16.73273, 16.91581, 17.0989, 
    17.28201, 17.46512, 17.64824, 17.83136, 18.01448, 18.19761, 18.38073, 
    18.56385, 18.74696, 18.93006, 19.11315, 19.29622, 19.47928, 19.66233, 
    19.84535, 20.02834, 20.21132, 20.39426, 20.57718, 20.76006, 20.94291, 
    21.12572, 21.30849, 21.49122, 21.67391, 21.85656, 22.03915, 22.2217, 
    22.40419, 22.58663, 22.76901, 22.95133, 23.13359, 23.31579, 23.49792, 
    23.67999, 23.86198, 24.04391, 24.22576, 24.40753, 24.58922, 24.77084, 
    24.95236, 25.13381, 25.31517, 25.49644, 25.67761, 25.8587, 26.03968, 
    26.22057, 26.40136, 26.58205, 26.76263, 26.94311, 27.12348, 27.30374, 
    27.48389, 27.66392, 27.84384, 28.02364, 28.20332, 28.38287, 28.56231, 
    28.74161, 28.92079, 29.09984, 29.27875, 29.45754, 29.63618, 29.81469, 
    29.99306, 30.17129, 30.34937, 30.52731, 30.70511, 30.88275, 31.06024, 
    31.23759, 31.41477, 31.5918, 31.76867, 31.94539, 32.12194, 32.29833, 
    32.47456, 32.65061, 32.8265, 33.00222, 33.17777, 33.35315, 33.52835, 
    33.70338, 33.87822, 34.05289, 34.22738, 34.40168, 34.57581, 34.74974, 
    34.92348, 35.09705, 35.27041, 35.44359, 35.61657, 35.78936, 35.96196, 
    36.13435, 36.30655, 36.47854, 36.65034, 36.82193, 36.99332, 37.1645, 
    37.33547, 37.50624, 37.6768, 37.84714, 38.01727, 38.18719, 38.3569, 
    38.52639, 38.69566, 38.86471, 39.03355, 39.20216, 39.37055, 39.53872, 
    39.70667, 39.87439, 40.04188, 40.20915, 40.37619, 40.543, 40.70957, 
    40.87592, 41.04203, 41.20792, 41.37356, 41.53897, 41.70415, 41.86909, 
    42.03379, 42.19825, 42.36247, 42.52645, 42.69019, 42.85368, 43.01694, 
    43.17995, 43.34271, 43.50523, 43.6675, 43.82952, 43.9913, 44.15283, 
    44.31411, 44.47514, 44.63592, 44.79644, 44.95672, 45.11674, 45.27651, 
    45.43603, 45.59529, 45.75429, 45.91304, 46.07154, 46.22977, 46.38775, 
    46.54548, 46.70294, 46.86014, 47.01709, 47.17377, 47.3302, 47.48636, 
    47.64227,
  -25.03907, -24.90766, -24.77599, -24.64406, -24.51188, -24.37943, 
    -24.24673, -24.11377, -23.98055, -23.84707, -23.71333, -23.57932, 
    -23.44506, -23.31053, -23.17574, -23.04069, -22.90537, -22.7698, 
    -22.63396, -22.49785, -22.36148, -22.22485, -22.08795, -21.95079, 
    -21.81336, -21.67567, -21.53771, -21.39949, -21.261, -21.12224, 
    -20.98321, -20.84392, -20.70436, -20.56454, -20.42444, -20.28408, 
    -20.14345, -20.00255, -19.86139, -19.71995, -19.57825, -19.43628, 
    -19.29403, -19.15152, -19.00874, -18.86569, -18.72237, -18.57878, 
    -18.43493, -18.2908, -18.1464, -18.00173, -17.85679, -17.71158, -17.5661, 
    -17.42035, -17.27434, -17.12805, -16.98149, -16.83466, -16.68756, 
    -16.54019, -16.39255, -16.24464, -16.09646, -15.94801, -15.79929, 
    -15.6503, -15.50104, -15.35151, -15.20171, -15.05164, -14.90131, 
    -14.7507, -14.59982, -14.44868, -14.29727, -14.14559, -13.99364, 
    -13.84142, -13.68894, -13.53619, -13.38317, -13.22988, -13.07633, 
    -12.92251, -12.76843, -12.61408, -12.45947, -12.30458, -12.14944, 
    -11.99403, -11.83836, -11.68242, -11.52622, -11.36976, -11.21303, 
    -11.05605, -10.8988, -10.74129, -10.58352, -10.42549, -10.2672, 
    -10.10865, -9.949849, -9.790786, -9.631464, -9.471887, -9.312053, 
    -9.151963, -8.991619, -8.83102, -8.670169, -8.509064, -8.347706, 
    -8.186097, -8.024237, -7.862127, -7.699767, -7.537159, -7.374302, 
    -7.211199, -7.047849, -6.884254, -6.720413, -6.556329, -6.392001, 
    -6.227432, -6.062621, -5.897569, -5.732277, -5.566748, -5.40098, 
    -5.234975, -5.068735, -4.902259, -4.73555, -4.568607, -4.401433, 
    -4.234028, -4.066394, -3.89853, -3.730439, -3.562121, -3.393578, 
    -3.22481, -3.05582, -2.886607, -2.717173, -2.54752, -2.377648, -2.207559, 
    -2.037254, -1.866733, -1.696, -1.525054, -1.353897, -1.182531, -1.010955, 
    -0.8391734, -0.6671857, -0.4949936, -0.3225986, -0.150002, 0.02279485, 
    0.1957904, 0.3689833, 0.542372, 0.7159552, 0.8897313, 1.063699, 1.237856, 
    1.412202, 1.586735, 1.761453, 1.936355, 2.111439, 2.286704, 2.462147, 
    2.637768, 2.813565, 2.989536, 3.165679, 3.341993, 3.518476, 3.695127, 
    3.871943, 4.048923, 4.226065, 4.403368, 4.58083, 4.758448, 4.936222, 
    5.114148, 5.292227, 5.470455, 5.64883, 5.827352, 6.006018, 6.184826, 
    6.363775, 6.542861, 6.722085, 6.901443, 7.080934, 7.260556, 7.440306, 
    7.620183, 7.800185, 7.98031, 8.160556, 8.34092, 8.521401, 8.701998, 
    8.882707, 9.063526, 9.244454, 9.425489, 9.606629, 9.78787, 9.969213, 
    10.15065, 10.33219, 10.51382, 10.69554, 10.87735, 11.05925, 11.24124, 
    11.42331, 11.60546, 11.78769, 11.96999, 12.15237, 12.33482, 12.51735, 
    12.69994, 12.88259, 13.06531, 13.24809, 13.43093, 13.61383, 13.79678, 
    13.97978, 14.16284, 14.34594, 14.52909, 14.71228, 14.89551, 15.07878, 
    15.26209, 15.44543, 15.6288, 15.8122, 15.99564, 16.17909, 16.36257, 
    16.54607, 16.72958, 16.91312, 17.09666, 17.28022, 17.46379, 17.64736, 
    17.83094, 18.01452, 18.1981, 18.38168, 18.56525, 18.74882, 18.93237, 
    19.11592, 19.29945, 19.48296, 19.66646, 19.84993, 20.03338, 20.21681, 
    20.40021, 20.58358, 20.76691, 20.95021, 21.13348, 21.3167, 21.49989, 
    21.68303, 21.86612, 22.04917, 22.23216, 22.41511, 22.59799, 22.78082, 
    22.9636, 23.14631, 23.32895, 23.51153, 23.69404, 23.87648, 24.05885, 
    24.24114, 24.42336, 24.6055, 24.78755, 24.96952, 25.15141, 25.33321, 
    25.51492, 25.69653, 25.87805, 26.05948, 26.2408, 26.42203, 26.60316, 
    26.78417, 26.96508, 27.14589, 27.32658, 27.50715, 27.68762, 27.86796, 
    28.04819, 28.2283, 28.40828, 28.58814, 28.76787, 28.94747, 29.12694, 
    29.30627, 29.48548, 29.66454, 29.84347, 30.02225, 30.2009, 30.3794, 
    30.55775, 30.73595, 30.91401, 31.09191, 31.26966, 31.44725, 31.62469, 
    31.80197, 31.97908, 32.15604, 32.33283, 32.50945, 32.68591, 32.86219, 
    33.03831, 33.21426, 33.39002, 33.56562, 33.74103, 33.91627, 34.09132, 
    34.2662, 34.44089, 34.61539, 34.7897, 34.96383, 35.13777, 35.31152, 
    35.48507, 35.65842, 35.83159, 36.00455, 36.17732, 36.34988, 36.52224, 
    36.6944, 36.86636, 37.03811, 37.20965, 37.38099, 37.55211, 37.72302, 
    37.89372, 38.06421, 38.23448, 38.40453, 38.57437, 38.74399, 38.91339, 
    39.08257, 39.25152, 39.42025, 39.58876, 39.75704, 39.9251, 40.09293, 
    40.26052, 40.42789, 40.59503, 40.76194, 40.92861, 41.09505, 41.26125, 
    41.42722, 41.59295, 41.75844, 41.92369, 42.08871, 42.25348, 42.41801, 
    42.5823, 42.74635, 42.91015, 43.0737, 43.23701, 43.40008, 43.5629, 
    43.72547, 43.88779, 44.04986, 44.21168, 44.37325, 44.53456, 44.69563, 
    44.85644, 45.017, 45.1773, 45.33735, 45.49715, 45.65668, 45.81596, 
    45.97499, 46.13375, 46.29226, 46.45051, 46.60849, 46.76622, 46.92369, 
    47.0809, 47.23784, 47.39453, 47.55095, 47.7071,
  -25.12111, -24.98959, -24.8578, -24.72575, -24.59344, -24.46088, -24.32805, 
    -24.19496, -24.06161, -23.928, -23.79413, -23.65999, -23.5256, -23.39094, 
    -23.25601, -23.12082, -22.98537, -22.84966, -22.71367, -22.57743, 
    -22.44092, -22.30414, -22.1671, -22.02979, -21.89221, -21.75437, 
    -21.61626, -21.47788, -21.33924, -21.20033, -21.06115, -20.9217, 
    -20.78198, -20.64199, -20.50174, -20.36121, -20.22042, -20.07935, 
    -19.93802, -19.79642, -19.65454, -19.5124, -19.36998, -19.2273, 
    -19.08434, -18.94111, -18.79762, -18.65384, -18.5098, -18.36549, 
    -18.22091, -18.07605, -17.93093, -17.78553, -17.63986, -17.49392, 
    -17.3477, -17.20122, -17.05446, -16.90743, -16.76013, -16.61256, 
    -16.46472, -16.3166, -16.16822, -16.01956, -15.87063, -15.72143, 
    -15.57196, -15.42221, -15.2722, -15.12191, -14.97136, -14.82053, 
    -14.66943, -14.51806, -14.36643, -14.21452, -14.06234, -13.90989, 
    -13.75718, -13.60419, -13.45094, -13.29742, -13.14363, -12.98957, 
    -12.83524, -12.68065, -12.52579, -12.37066, -12.21526, -12.0596, 
    -11.90368, -11.74749, -11.59103, -11.43431, -11.27733, -11.12008, 
    -10.96257, -10.8048, -10.64677, -10.48847, -10.32991, -10.17109, 
    -10.01201, -9.852676, -9.69308, -9.533224, -9.373111, -9.212741, 
    -9.052114, -8.891231, -8.730093, -8.5687, -8.407053, -8.245152, -8.083, 
    -7.920595, -7.757939, -7.595033, -7.431877, -7.268472, -7.104819, 
    -6.940919, -6.776772, -6.61238, -6.447742, -6.282861, -6.117736, 
    -5.95237, -5.786762, -5.620914, -5.454825, -5.288499, -5.121935, 
    -4.955135, -4.788099, -4.620828, -4.453324, -4.285587, -4.11762, 
    -3.949421, -3.780993, -3.612337, -3.443454, -3.274345, -3.105011, 
    -2.935453, -2.765673, -2.595671, -2.42545, -2.255009, -2.084351, 
    -1.913477, -1.742387, -1.571084, -1.399567, -1.22784, -1.055903, 
    -0.8837567, -0.7114035, -0.5388445, -0.3660809, -0.1931142, -0.01994582, 
    0.1534228, 0.3269903, 0.5007551, 0.6747158, 0.8488709, 1.023219, 
    1.197758, 1.372488, 1.547405, 1.72251, 1.897799, 2.073272, 2.248927, 
    2.424763, 2.600777, 2.776969, 2.953336, 3.129876, 3.306589, 3.483472, 
    3.660524, 3.837743, 4.015127, 4.192674, 4.370384, 4.548253, 4.72628, 
    4.904464, 5.082802, 5.261293, 5.439935, 5.618726, 5.797664, 5.976747, 
    6.155973, 6.335341, 6.514849, 6.694494, 6.874275, 7.05419, 7.234237, 
    7.414413, 7.594718, 7.775147, 7.955701, 8.136377, 8.317173, 8.498086, 
    8.679115, 8.860258, 9.041512, 9.222877, 9.404347, 9.585924, 9.767605, 
    9.949386, 10.13127, 10.31324, 10.49531, 10.67748, 10.85973, 11.04208, 
    11.22451, 11.40702, 11.58962, 11.77229, 11.95504, 12.13787, 12.32077, 
    12.50374, 12.68678, 12.86989, 13.05306, 13.23629, 13.41958, 13.60293, 
    13.78633, 13.96979, 14.1533, 14.33685, 14.52045, 14.7041, 14.88778, 
    15.07151, 15.25527, 15.43907, 15.6229, 15.80676, 15.99064, 16.17455, 
    16.35849, 16.54244, 16.72642, 16.91041, 17.09441, 17.27843, 17.46245, 
    17.64648, 17.83052, 18.01455, 18.19859, 18.38263, 18.56666, 18.75068, 
    18.93469, 19.1187, 19.30268, 19.48666, 19.67061, 19.85454, 20.03845, 
    20.22233, 20.40618, 20.59001, 20.7738, 20.95756, 21.14128, 21.32495, 
    21.50859, 21.69219, 21.87574, 22.05923, 22.24268, 22.42608, 22.60942, 
    22.7927, 22.97592, 23.15908, 23.34218, 23.52521, 23.70817, 23.89106, 
    24.07387, 24.25661, 24.43927, 24.62186, 24.80436, 24.98677, 25.1691, 
    25.35134, 25.53349, 25.71555, 25.89751, 26.07938, 26.26114, 26.4428, 
    26.62436, 26.80582, 26.98717, 27.1684, 27.34953, 27.53054, 27.71143, 
    27.89221, 28.07287, 28.2534, 28.43381, 28.6141, 28.79425, 28.97428, 
    29.15417, 29.33393, 29.51356, 29.69304, 29.87239, 30.05159, 30.23065, 
    30.40957, 30.58833, 30.76695, 30.94542, 31.12373, 31.30189, 31.47989, 
    31.65774, 31.83542, 32.01294, 32.1903, 32.36749, 32.54452, 32.72137, 
    32.89806, 33.07457, 33.25092, 33.42708, 33.60306, 33.77887, 33.9545, 
    34.12994, 34.3052, 34.48028, 34.65516, 34.82986, 35.00437, 35.17869, 
    35.35281, 35.52674, 35.70048, 35.87402, 36.04735, 36.22049, 36.39342, 
    36.56615, 36.73868, 36.911, 37.08311, 37.25502, 37.42671, 37.59819, 
    37.76947, 37.94052, 38.11136, 38.28199, 38.45239, 38.62258, 38.79255, 
    38.96229, 39.13181, 39.30111, 39.47018, 39.63903, 39.80765, 39.97604, 
    40.1442, 40.31214, 40.47984, 40.6473, 40.81454, 40.98154, 41.1483, 
    41.31483, 41.48111, 41.64716, 41.81297, 41.97854, 42.14387, 42.30896, 
    42.4738, 42.6384, 42.80275, 42.96686, 43.13072, 43.29434, 43.4577, 
    43.62082, 43.78369, 43.9463, 44.10867, 44.27078, 44.43264, 44.59425, 
    44.7556, 44.9167, 45.07754, 45.23812, 45.39846, 45.55853, 45.71834, 
    45.8779, 46.0372, 46.19623, 46.35501, 46.51353, 46.67178, 46.82978, 
    46.98751, 47.14497, 47.30218, 47.45912, 47.6158, 47.77221,
  -25.20343, -25.07178, -24.93987, -24.8077, -24.67528, -24.54259, -24.40963, 
    -24.27642, -24.14294, -24.0092, -23.8752, -23.74094, -23.60641, 
    -23.47161, -23.33655, -23.20123, -23.06564, -22.92979, -22.79367, 
    -22.65728, -22.52063, -22.38371, -22.24652, -22.10906, -21.97134, 
    -21.83335, -21.69509, -21.55656, -21.41776, -21.27869, -21.13935, 
    -20.99975, -20.85987, -20.71972, -20.57931, -20.43862, -20.29766, 
    -20.15643, -20.01493, -19.87316, -19.73111, -19.5888, -19.44621, 
    -19.30335, -19.16022, -19.01681, -18.87313, -18.72918, -18.58496, 
    -18.44047, -18.2957, -18.15066, -18.00534, -17.85975, -17.71389, 
    -17.56776, -17.42135, -17.27467, -17.12772, -16.98049, -16.83299, 
    -16.68521, -16.53717, -16.38885, -16.24026, -16.09139, -15.94225, 
    -15.79284, -15.64315, -15.49319, -15.34296, -15.19246, -15.04168, 
    -14.89064, -14.73932, -14.58772, -14.43586, -14.28372, -14.13132, 
    -13.97864, -13.82569, -13.67247, -13.51898, -13.36522, -13.21119, 
    -13.05689, -12.90232, -12.74749, -12.59238, -12.43701, -12.28136, 
    -12.12545, -11.96927, -11.81283, -11.65612, -11.49914, -11.3419, 
    -11.18439, -11.02662, -10.86858, -10.71028, -10.55171, -10.39289, 
    -10.2338, -10.07444, -9.914832, -9.754959, -9.594826, -9.434433, 
    -9.273781, -9.11287, -8.951702, -8.790277, -8.628596, -8.46666, 
    -8.304467, -8.14202, -7.979321, -7.816368, -7.653162, -7.489706, 
    -7.325999, -7.162042, -6.997836, -6.833382, -6.66868, -6.503732, 
    -6.338538, -6.1731, -6.007417, -5.841492, -5.675324, -5.508915, 
    -5.342266, -5.175378, -5.008252, -4.840888, -4.673288, -4.505453, 
    -4.337383, -4.16908, -4.000546, -3.83178, -3.662785, -3.49356, -3.324108, 
    -3.15443, -2.984526, -2.814399, -2.644048, -2.473475, -2.302682, 
    -2.13167, -1.96044, -1.788993, -1.61733, -1.445453, -1.273364, -1.101063, 
    -0.9285516, -0.7558315, -0.582904, -0.4097705, -0.2364323, -0.06289089, 
    0.1108523, 0.2847958, 0.4589382, 0.633278, 0.8078137, 0.9825438, 
    1.157467, 1.332581, 1.507885, 1.683377, 1.859056, 2.03492, 2.210967, 
    2.387196, 2.563606, 2.740193, 2.916958, 3.093898, 3.271011, 3.448296, 
    3.625751, 3.803374, 3.981164, 4.159118, 4.337236, 4.515515, 4.693953, 
    4.872549, 5.0513, 5.230206, 5.409263, 5.588471, 5.767827, 5.94733, 
    6.126976, 6.306766, 6.486696, 6.666765, 6.846971, 7.027312, 7.207786, 
    7.38839, 7.569123, 7.749983, 7.930969, 8.112077, 8.293305, 8.474652, 
    8.656116, 8.837695, 9.019386, 9.201188, 9.383099, 9.565114, 9.747235, 
    9.929458, 10.11178, 10.2942, 10.47672, 10.65932, 10.84202, 11.02481, 
    11.20769, 11.39065, 11.57369, 11.75682, 11.94002, 12.12329, 12.30664, 
    12.49007, 12.67356, 12.85712, 13.04074, 13.22442, 13.40817, 13.59197, 
    13.77583, 13.95974, 14.1437, 14.32771, 14.51177, 14.69587, 14.88002, 
    15.0642, 15.24842, 15.43267, 15.61696, 15.80128, 15.98562, 16.16999, 
    16.35439, 16.5388, 16.72324, 16.90769, 17.09215, 17.27662, 17.46111, 
    17.6456, 17.8301, 18.01459, 18.19909, 18.38358, 18.56808, 18.75256, 
    18.93703, 19.12149, 19.30594, 19.49037, 19.67478, 19.85917, 20.04354, 
    20.22788, 20.41219, 20.59647, 20.78072, 20.96494, 21.14911, 21.33325, 
    21.51735, 21.7014, 21.8854, 22.06935, 22.25326, 22.43711, 22.6209, 
    22.80464, 22.98831, 23.17192, 23.35547, 23.53895, 23.72236, 23.9057, 
    24.08897, 24.27216, 24.45527, 24.6383, 24.82125, 25.00411, 25.18688, 
    25.36957, 25.55216, 25.73466, 25.91707, 26.09937, 26.28158, 26.46368, 
    26.64568, 26.82758, 27.00936, 27.19103, 27.37259, 27.55404, 27.73537, 
    27.91658, 28.09767, 28.27863, 28.45947, 28.64019, 28.82077, 29.00122, 
    29.18154, 29.36173, 29.54177, 29.72168, 29.90145, 30.08108, 30.26055, 
    30.43989, 30.61907, 30.79811, 30.97699, 31.15571, 31.33428, 31.5127, 
    31.69095, 31.86904, 32.04697, 32.22474, 32.40233, 32.57976, 32.75702, 
    32.9341, 33.11102, 33.28775, 33.46431, 33.64069, 33.81689, 33.99291, 
    34.16875, 34.34439, 34.51986, 34.69513, 34.87022, 35.04511, 35.21981, 
    35.39431, 35.56862, 35.74273, 35.91665, 36.09035, 36.26387, 36.43717, 
    36.61027, 36.78316, 36.95585, 37.12833, 37.3006, 37.47266, 37.6445, 
    37.81613, 37.98754, 38.15874, 38.32971, 38.50047, 38.67101, 38.84132, 
    39.01142, 39.18129, 39.35093, 39.52034, 39.68953, 39.85849, 40.02722, 
    40.19572, 40.36398, 40.53202, 40.69981, 40.86738, 41.0347, 41.20179, 
    41.36864, 41.53526, 41.70163, 41.86776, 42.03364, 42.19929, 42.36469, 
    42.52984, 42.69475, 42.85941, 43.02383, 43.188, 43.35191, 43.51558, 
    43.679, 43.84216, 44.00507, 44.16773, 44.33014, 44.49229, 44.65419, 
    44.81583, 44.97721, 45.13834, 45.29921, 45.45982, 45.62017, 45.78027, 
    45.9401, 46.09967, 46.25898, 46.41803, 46.57681, 46.73534, 46.8936, 
    47.05159, 47.20932, 47.36679, 47.52399, 47.68092, 47.83759,
  -25.28601, -25.15425, -25.02222, -24.88993, -24.75738, -24.62457, 
    -24.49149, -24.35815, -24.22455, -24.09068, -23.95655, -23.82215, 
    -23.68749, -23.55256, -23.41737, -23.28191, -23.14618, -23.01019, 
    -22.87393, -22.7374, -22.60061, -22.46354, -22.32621, -22.18861, 
    -22.05074, -21.9126, -21.77419, -21.63551, -21.49656, -21.35733, 
    -21.21784, -21.07808, -20.93804, -20.79774, -20.65716, -20.51631, 
    -20.37518, -20.23379, -20.09212, -19.95018, -19.80796, -19.66548, 
    -19.52271, -19.37968, -19.23637, -19.09279, -18.94893, -18.8048, 
    -18.6604, -18.51572, -18.37077, -18.22554, -18.08004, -17.93426, 
    -17.78821, -17.64188, -17.49528, -17.3484, -17.20125, -17.05383, 
    -16.90612, -16.75815, -16.6099, -16.46137, -16.31257, -16.1635, 
    -16.01415, -15.86453, -15.71463, -15.56445, -15.41401, -15.26329, 
    -15.11229, -14.96102, -14.80948, -14.65766, -14.50557, -14.35321, 
    -14.20057, -14.04766, -13.89448, -13.74103, -13.5873, -13.43331, 
    -13.27904, -13.1245, -12.96968, -12.8146, -12.65925, -12.50363, 
    -12.34773, -12.19157, -12.03514, -11.87844, -11.72147, -11.56424, 
    -11.40674, -11.24897, -11.09093, -10.93263, -10.77406, -10.61523, 
    -10.45613, -10.29677, -10.13714, -9.977255, -9.817104, -9.656693, 
    -9.496019, -9.335085, -9.173891, -9.012437, -8.850725, -8.688754, 
    -8.526526, -8.364041, -8.201301, -8.038304, -7.875054, -7.711549, 
    -7.547791, -7.383781, -7.21952, -7.055007, -6.890245, -6.725234, 
    -6.559974, -6.394466, -6.228713, -6.062713, -5.896469, -5.729981, 
    -5.563251, -5.396278, -5.229064, -5.061611, -4.893918, -4.725987, 
    -4.55782, -4.389417, -4.220778, -4.051907, -3.882802, -3.713466, -3.5439, 
    -3.374104, -3.20408, -3.033829, -2.863352, -2.692651, -2.521726, 
    -2.350579, -2.179211, -2.007624, -1.835818, -1.663795, -1.491557, 
    -1.319104, -1.146438, -0.9735597, -0.8004714, -0.6271741, -0.4536691, 
    -0.279958, -0.1060421, 0.06807715, 0.2423982, 0.4169197, 0.5916401, 
    0.7665579, 0.9416716, 1.11698, 1.29248, 1.468173, 1.644054, 1.820124, 
    1.99638, 2.172822, 2.349446, 2.526252, 2.703238, 2.880402, 3.057742, 
    3.235257, 3.412946, 3.590806, 3.768835, 3.947032, 4.125396, 4.303924, 
    4.482614, 4.661465, 4.840474, 5.019641, 5.198963, 5.378438, 5.558064, 
    5.737841, 5.917764, 6.097834, 6.278047, 6.458402, 6.638896, 6.81953, 
    7.000298, 7.181201, 7.362235, 7.5434, 7.724692, 7.90611, 8.087652, 
    8.269317, 8.4511, 8.633001, 8.815018, 8.997149, 9.17939, 9.36174, 
    9.544198, 9.726761, 9.909427, 10.09219, 10.27506, 10.45802, 10.64108, 
    10.82422, 11.00746, 11.19078, 11.37419, 11.55769, 11.74126, 11.92491, 
    12.10864, 12.29245, 12.47632, 12.66027, 12.84428, 13.02836, 13.2125, 
    13.3967, 13.58096, 13.76527, 13.94964, 14.13406, 14.31853, 14.50305, 
    14.68761, 14.87221, 15.05685, 15.24153, 15.42625, 15.611, 15.79577, 
    15.98058, 16.16541, 16.35027, 16.53514, 16.72004, 16.90495, 17.08987, 
    17.27481, 17.45976, 17.64471, 17.82967, 18.01463, 18.19959, 18.38455, 
    18.5695, 18.75444, 18.93938, 19.1243, 19.30921, 19.4941, 19.67898, 
    19.86383, 20.04865, 20.23346, 20.41823, 20.60297, 20.78768, 20.97236, 
    21.15699, 21.34159, 21.52614, 21.71065, 21.89511, 22.07952, 22.26389, 
    22.44819, 22.63244, 22.81664, 23.00076, 23.18483, 23.36884, 23.55277, 
    23.73663, 23.92043, 24.10414, 24.28778, 24.47134, 24.65482, 24.83822, 
    25.02153, 25.20476, 25.38789, 25.57093, 25.75387, 25.93672, 26.11947, 
    26.30212, 26.48467, 26.66711, 26.84945, 27.03167, 27.21378, 27.39578, 
    27.57766, 27.75943, 27.94107, 28.12259, 28.30399, 28.48527, 28.66641, 
    28.84742, 29.02831, 29.20905, 29.38966, 29.57014, 29.75047, 29.93066, 
    30.11071, 30.29061, 30.47036, 30.64996, 30.82941, 31.00871, 31.18785, 
    31.36684, 31.54566, 31.72433, 31.90283, 32.08117, 32.25934, 32.43734, 
    32.61517, 32.79284, 32.97032, 33.14764, 33.32477, 33.50173, 33.6785, 
    33.8551, 34.03151, 34.20774, 34.38378, 34.55963, 34.73529, 34.91076, 
    35.08604, 35.26112, 35.43601, 35.6107, 35.78519, 35.95948, 36.13357, 
    36.30745, 36.48113, 36.6546, 36.82787, 37.00092, 37.17376, 37.3464, 
    37.51882, 37.69102, 37.86301, 38.03478, 38.20633, 38.37767, 38.54878, 
    38.71967, 38.89034, 39.06078, 39.23099, 39.40098, 39.57074, 39.74027, 
    39.90957, 40.07864, 40.24747, 40.41607, 40.58444, 40.75257, 40.92046, 
    41.08812, 41.25553, 41.42271, 41.58964, 41.75633, 41.92278, 42.08899, 
    42.25495, 42.42066, 42.58613, 42.75135, 42.91632, 43.08105, 43.24552, 
    43.40974, 43.57371, 43.73743, 43.90089, 44.06411, 44.22706, 44.38976, 
    44.5522, 44.71439, 44.87632, 45.03799, 45.19941, 45.36056, 45.52145, 
    45.68208, 45.84246, 46.00256, 46.16241, 46.32199, 46.48132, 46.64037, 
    46.79916, 46.95769, 47.11595, 47.27394, 47.43167, 47.58913, 47.74632, 
    47.90325,
  -25.36886, -25.23698, -25.10483, -24.97242, -24.83975, -24.70681, 
    -24.57361, -24.44015, -24.30642, -24.17243, -24.03817, -23.90364, 
    -23.76885, -23.63379, -23.49846, -23.36287, -23.227, -23.09087, 
    -22.95447, -22.8178, -22.68087, -22.54366, -22.40618, -22.26843, 
    -22.13041, -21.99213, -21.85357, -21.71473, -21.57563, -21.43625, 
    -21.29661, -21.15668, -21.01649, -20.87602, -20.73528, -20.59427, 
    -20.45298, -20.31142, -20.16959, -20.02748, -19.8851, -19.74244, 
    -19.5995, -19.45629, -19.31281, -19.16905, -19.02501, -18.8807, 
    -18.73612, -18.59126, -18.44612, -18.3007, -18.15501, -18.00905, 
    -17.8628, -17.71628, -17.56949, -17.42242, -17.27507, -17.12744, 
    -16.97954, -16.83137, -16.68291, -16.53418, -16.38517, -16.23589, 
    -16.08633, -15.9365, -15.78638, -15.636, -15.48533, -15.33439, -15.18318, 
    -15.03169, -14.87992, -14.72788, -14.57557, -14.42297, -14.27011, 
    -14.11697, -13.96355, -13.80986, -13.6559, -13.50167, -13.34716, 
    -13.19238, -13.03732, -12.88199, -12.72639, -12.57052, -12.41438, 
    -12.25797, -12.10128, -11.94433, -11.7871, -11.62961, -11.47185, 
    -11.31382, -11.15552, -10.99695, -10.83811, -10.67901, -10.51964, 
    -10.36001, -10.20011, -10.03995, -9.879519, -9.718827, -9.557873, 
    -9.396656, -9.235177, -9.073437, -8.911436, -8.749176, -8.586657, 
    -8.423879, -8.260842, -8.097549, -7.934, -7.770195, -7.606135, -7.441822, 
    -7.277254, -7.112434, -6.947363, -6.782041, -6.616468, -6.450647, 
    -6.284577, -6.11826, -5.951696, -5.784887, -5.617834, -5.450536, 
    -5.282996, -5.115214, -4.947192, -4.77893, -4.610429, -4.441691, 
    -4.272716, -4.103506, -3.934061, -3.764383, -3.594473, -3.424332, 
    -3.253962, -3.083362, -2.912535, -2.741482, -2.570204, -2.398702, 
    -2.226978, -2.055032, -1.882866, -1.710482, -1.53788, -1.365062, 
    -1.192029, -1.018783, -0.845325, -0.6716564, -0.4977786, -0.3236931, 
    -0.1494012, 0.0250956, 0.1997958, 0.3746979, 0.5498005, 0.7251019, 
    0.9006008, 1.076295, 1.252185, 1.428266, 1.604539, 1.781002, 1.957652, 
    2.134489, 2.31151, 2.488714, 2.6661, 2.843665, 3.021408, 3.199327, 
    3.377421, 3.555687, 3.734125, 3.912732, 4.091506, 4.270445, 4.449549, 
    4.628814, 4.808239, 4.987823, 5.167563, 5.347458, 5.527505, 5.707704, 
    5.888051, 6.068544, 6.249183, 6.429965, 6.610887, 6.791949, 6.973147, 
    7.154481, 7.335948, 7.517546, 7.699272, 7.881126, 8.063105, 8.245205, 
    8.427427, 8.609768, 8.792225, 8.974796, 9.157479, 9.340273, 9.523175, 
    9.706182, 9.889294, 10.07251, 10.25582, 10.43923, 10.62273, 10.80633, 
    10.99002, 11.17379, 11.35765, 11.5416, 11.72563, 11.90973, 12.09392, 
    12.27818, 12.46251, 12.64691, 12.83138, 13.01591, 13.20051, 13.38517, 
    13.56989, 13.75466, 13.93949, 14.12437, 14.3093, 14.49428, 14.6793, 
    14.86436, 15.04947, 15.23461, 15.41979, 15.605, 15.79024, 15.97551, 
    16.1608, 16.34612, 16.53146, 16.71682, 16.9022, 17.08759, 17.27299, 
    17.4584, 17.64382, 17.82924, 18.01467, 18.20009, 18.38551, 18.57093, 
    18.75634, 18.94174, 19.12712, 19.3125, 19.49785, 19.68319, 19.86851, 
    20.0538, 20.23907, 20.4243, 20.60951, 20.79468, 20.97981, 21.16491, 
    21.34997, 21.53499, 21.71996, 21.90488, 22.08975, 22.27457, 22.45934, 
    22.64404, 22.8287, 23.01328, 23.19781, 23.38227, 23.56666, 23.75098, 
    23.93522, 24.11939, 24.30349, 24.4875, 24.67144, 24.85528, 25.03905, 
    25.22272, 25.4063, 25.58979, 25.77319, 25.95648, 26.13968, 26.32277, 
    26.50576, 26.68865, 26.87143, 27.05409, 27.23664, 27.41908, 27.60141, 
    27.78361, 27.96569, 28.14765, 28.32948, 28.51119, 28.69277, 28.87421, 
    29.05552, 29.2367, 29.41774, 29.59864, 29.7794, 29.96002, 30.14049, 
    30.32081, 30.50098, 30.68101, 30.86088, 31.04059, 31.22015, 31.39955, 
    31.57879, 31.75787, 31.93678, 32.11553, 32.29411, 32.47252, 32.65076, 
    32.82883, 33.00672, 33.18444, 33.36197, 33.53933, 33.7165, 33.8935, 
    34.0703, 34.24693, 34.42336, 34.5996, 34.77565, 34.95151, 35.12717, 
    35.30264, 35.47791, 35.65298, 35.82785, 36.00252, 36.17699, 36.35125, 
    36.5253, 36.69914, 36.87278, 37.0462, 37.21941, 37.39241, 37.5652, 
    37.73777, 37.91011, 38.08224, 38.25416, 38.42585, 38.59731, 38.76855, 
    38.93957, 39.11036, 39.28093, 39.45126, 39.62136, 39.79124, 39.96088, 
    40.13029, 40.29946, 40.4684, 40.6371, 40.80556, 40.97379, 41.14177, 
    41.30951, 41.47702, 41.64428, 41.81129, 41.97806, 42.14458, 42.31086, 
    42.47689, 42.64268, 42.80821, 42.97349, 43.13852, 43.3033, 43.46783, 
    43.6321, 43.79612, 43.95989, 44.1234, 44.28665, 44.44965, 44.61238, 
    44.77486, 44.93708, 45.09904, 45.26074, 45.42218, 45.58335, 45.74426, 
    45.90491, 46.0653, 46.22542, 46.38528, 46.54487, 46.7042, 46.86325, 
    47.02205, 47.18058, 47.33883, 47.49682, 47.65454, 47.81199, 47.96917,
  -25.45198, -25.31998, -25.18772, -25.05519, -24.9224, -24.78934, -24.65601, 
    -24.52242, -24.38857, -24.25445, -24.12006, -23.9854, -23.85048, 
    -23.71529, -23.57983, -23.4441, -23.3081, -23.17183, -23.03529, 
    -22.89848, -22.7614, -22.62405, -22.48643, -22.34854, -22.21037, 
    -22.07193, -21.93322, -21.79424, -21.65499, -21.51546, -21.37565, 
    -21.23557, -21.09522, -20.9546, -20.8137, -20.67252, -20.53107, 
    -20.38934, -20.24734, -20.10506, -19.96251, -19.81968, -19.67657, 
    -19.53319, -19.38953, -19.24559, -19.10138, -18.95689, -18.81212, 
    -18.66708, -18.52175, -18.37615, -18.23027, -18.08412, -17.93769, 
    -17.79097, -17.64398, -17.49672, -17.34917, -17.20135, -17.05325, 
    -16.90487, -16.75621, -16.60727, -16.45806, -16.30857, -16.1588, 
    -16.00875, -15.85843, -15.70782, -15.55694, -15.40579, -15.25435, 
    -15.10264, -14.95065, -14.79838, -14.64584, -14.49302, -14.33993, 
    -14.18655, -14.03291, -13.87898, -13.72478, -13.57031, -13.41556, 
    -13.26054, -13.10524, -12.94967, -12.79382, -12.6377, -12.48131, 
    -12.32464, -12.1677, -12.01049, -11.85301, -11.69526, -11.53724, 
    -11.37894, -11.22038, -11.06154, -10.90244, -10.74307, -10.58343, 
    -10.42352, -10.26335, -10.10291, -9.942204, -9.781232, -9.619995, 
    -9.458495, -9.296731, -9.134704, -8.972415, -8.809864, -8.647052, 
    -8.48398, -8.320648, -8.157058, -7.993209, -7.829103, -7.66474, 
    -7.500121, -7.335248, -7.17012, -7.004738, -6.839104, -6.673218, 
    -6.507082, -6.340695, -6.174059, -6.007175, -5.840044, -5.672666, 
    -5.505043, -5.337175, -5.169065, -5.000711, -4.832117, -4.663281, 
    -4.494207, -4.324895, -4.155345, -3.985559, -3.815538, -3.645284, 
    -3.474797, -3.304078, -3.133129, -2.96195, -2.790544, -2.618911, 
    -2.447053, -2.27497, -2.102665, -1.930138, -1.75739, -1.584424, 
    -1.411239, -1.237839, -1.064223, -0.8903942, -0.7163529, -0.5421007, 
    -0.3676393, -0.1929699, -0.01809411, 0.1569867, 0.332271, 0.5077572, 
    0.683444, 0.8593296, 1.035413, 1.211691, 1.388164, 1.56483, 1.741687, 
    1.918733, 2.095967, 2.273386, 2.450991, 2.628778, 2.806746, 2.984894, 
    3.163218, 3.341719, 3.520394, 3.699242, 3.878259, 4.057446, 4.236799, 
    4.416318, 4.596, 4.775843, 4.955846, 5.136006, 5.316322, 5.496792, 
    5.677414, 5.858186, 6.039106, 6.220172, 6.401383, 6.582736, 6.764228, 
    6.945858, 7.127625, 7.309526, 7.49156, 7.673723, 7.856013, 8.03843, 
    8.220971, 8.403633, 8.586415, 8.769315, 8.952329, 9.135457, 9.318696, 
    9.502044, 9.685498, 9.869057, 10.05272, 10.23648, 10.42034, 10.60429, 
    10.78834, 10.97248, 11.15671, 11.34103, 11.52543, 11.70991, 11.89447, 
    12.07911, 12.26383, 12.44862, 12.63348, 12.81841, 13.0034, 13.18846, 
    13.37358, 13.55876, 13.74399, 13.92929, 14.11463, 14.30002, 14.48546, 
    14.67095, 14.85648, 15.04204, 15.22765, 15.41329, 15.59897, 15.78468, 
    15.97041, 16.15617, 16.34196, 16.52777, 16.71359, 16.89943, 17.08529, 
    17.27116, 17.45704, 17.64292, 17.82881, 18.0147, 18.20059, 18.38648, 
    18.57237, 18.75824, 18.94411, 19.12996, 19.3158, 19.50163, 19.68743, 
    19.87321, 20.05897, 20.2447, 20.4304, 20.61607, 20.80171, 20.98731, 
    21.17287, 21.3584, 21.54387, 21.72931, 21.91469, 22.10003, 22.28531, 
    22.47054, 22.65571, 22.84082, 23.02587, 23.21085, 23.39577, 23.58062, 
    23.76539, 23.9501, 24.13473, 24.31928, 24.50375, 24.68813, 24.87244, 
    25.05665, 25.24078, 25.42481, 25.60875, 25.79259, 25.97634, 26.15999, 
    26.34353, 26.52697, 26.7103, 26.89352, 27.07663, 27.25962, 27.44251, 
    27.62527, 27.80791, 27.99043, 28.17283, 28.3551, 28.53724, 28.71926, 
    28.90114, 29.08288, 29.26449, 29.44596, 29.62729, 29.80848, 29.98952, 
    30.17042, 30.35117, 30.53176, 30.71221, 30.8925, 31.07264, 31.25261, 
    31.43243, 31.61209, 31.79158, 31.97091, 32.15007, 32.32906, 32.50788, 
    32.68653, 32.865, 33.0433, 33.22142, 33.39936, 33.57711, 33.75469, 
    33.93208, 34.10929, 34.2863, 34.46313, 34.63976, 34.81621, 34.99245, 
    35.16851, 35.34436, 35.52002, 35.69547, 35.87072, 36.04577, 36.22062, 
    36.39525, 36.56968, 36.7439, 36.9179, 37.0917, 37.26528, 37.43865, 
    37.6118, 37.78473, 37.95744, 38.12994, 38.3022, 38.47425, 38.64608, 
    38.81767, 38.98904, 39.16019, 39.3311, 39.50178, 39.67223, 39.84245, 
    40.01243, 40.18218, 40.35169, 40.52097, 40.69001, 40.8588, 41.02736, 
    41.19567, 41.36375, 41.53157, 41.69916, 41.8665, 42.03359, 42.20044, 
    42.36703, 42.53338, 42.69947, 42.86532, 43.03091, 43.19626, 43.36134, 
    43.52618, 43.69076, 43.85508, 44.01915, 44.18295, 44.3465, 44.50979, 
    44.67282, 44.83559, 44.9981, 45.16035, 45.32234, 45.48406, 45.64552, 
    45.80671, 45.96764, 46.12831, 46.2887, 46.44884, 46.6087, 46.7683, 
    46.92763, 47.08669, 47.24548, 47.404, 47.56225, 47.72023, 47.87794, 
    48.03538,
  -25.53538, -25.40326, -25.27088, -25.13823, -25.00532, -24.87214, 
    -24.73869, -24.60497, -24.47099, -24.33674, -24.20223, -24.06744, 
    -23.93239, -23.79706, -23.66147, -23.52561, -23.38947, -23.25307, 
    -23.11639, -22.97944, -22.84222, -22.70473, -22.56696, -22.42892, 
    -22.29061, -22.15203, -22.01316, -21.87403, -21.73462, -21.59494, 
    -21.45498, -21.31475, -21.17424, -21.03345, -20.89239, -20.75105, 
    -20.60944, -20.46755, -20.32538, -20.18293, -20.04021, -19.89721, 
    -19.75393, -19.61037, -19.46654, -19.32242, -19.17803, -19.03336, 
    -18.88841, -18.74318, -18.59767, -18.45189, -18.30582, -18.15948, 
    -18.01285, -17.86595, -17.71876, -17.5713, -17.42356, -17.27554, 
    -17.12723, -16.97865, -16.82979, -16.68065, -16.53123, -16.38153, 
    -16.23155, -16.08129, -15.93075, -15.77993, -15.62884, -15.47746, 
    -15.32581, -15.17387, -15.02166, -14.86917, -14.7164, -14.56335, 
    -14.41003, -14.25642, -14.10254, -13.94838, -13.79395, -13.63923, 
    -13.48425, -13.32898, -13.17344, -13.01762, -12.86153, -12.70516, 
    -12.54851, -12.3916, -12.2344, -12.07694, -11.9192, -11.76119, -11.6029, 
    -11.44434, -11.28551, -11.12642, -10.96704, -10.8074, -10.64749, 
    -10.48731, -10.32686, -10.16615, -10.00516, -9.843908, -9.682389, 
    -9.520605, -9.358555, -9.19624, -9.033662, -8.870819, -8.707714, 
    -8.544348, -8.380719, -8.21683, -8.052681, -7.888273, -7.723607, 
    -7.558682, -7.393502, -7.228065, -7.062373, -6.896426, -6.730226, 
    -6.563773, -6.397069, -6.230113, -6.062907, -5.895453, -5.72775, 
    -5.559801, -5.391605, -5.223164, -5.054478, -4.88555, -4.71638, 
    -4.546968, -4.377316, -4.207426, -4.037298, -3.866933, -3.696332, 
    -3.525498, -3.35443, -3.18313, -3.011599, -2.839838, -2.667849, 
    -2.495633, -2.323191, -2.150525, -1.977635, -1.804523, -1.631191, 
    -1.457639, -1.283869, -1.109882, -0.9356807, -0.7612652, -0.5866373, 
    -0.4117985, -0.2367502, -0.06149377, 0.1139692, 0.2896371, 0.4655087, 
    0.6415823, 0.8178563, 0.9943292, 1.170999, 1.347865, 1.524925, 1.702178, 
    1.879622, 2.057254, 2.235075, 2.413081, 2.591271, 2.769644, 2.948197, 
    3.12693, 3.30584, 3.484925, 3.664184, 3.843615, 4.023215, 4.202985, 
    4.38292, 4.56302, 4.743283, 4.923707, 5.10429, 5.285029, 5.465924, 
    5.646972, 5.828171, 6.009519, 6.191015, 6.372656, 6.55444, 6.736366, 
    6.918431, 7.100633, 7.28297, 7.46544, 7.648042, 7.830772, 8.01363, 
    8.196612, 8.379717, 8.562943, 8.746286, 8.929747, 9.11332, 9.297007, 
    9.480803, 9.664706, 9.848716, 10.03283, 10.21704, 10.40135, 10.58576, 
    10.77026, 10.95486, 11.13954, 11.32432, 11.50917, 11.69411, 11.87913, 
    12.06423, 12.24941, 12.43466, 12.61998, 12.80537, 12.99082, 13.17635, 
    13.36193, 13.54757, 13.73327, 13.91903, 14.10484, 14.29069, 14.4766, 
    14.66255, 14.84855, 15.03458, 15.22066, 15.40677, 15.59291, 15.77908, 
    15.96529, 16.15152, 16.33777, 16.52405, 16.71034, 16.89665, 17.08298, 
    17.26932, 17.45567, 17.64202, 17.82838, 18.01474, 18.2011, 18.38746, 
    18.57381, 18.76016, 18.9465, 19.13282, 19.31913, 19.50542, 19.69169, 
    19.87794, 20.06417, 20.25037, 20.43654, 20.62267, 20.80878, 20.99485, 
    21.18088, 21.36687, 21.55281, 21.73871, 21.92456, 22.11036, 22.29611, 
    22.4818, 22.66743, 22.853, 23.03852, 23.22396, 23.40934, 23.59465, 
    23.77989, 23.96505, 24.15014, 24.33515, 24.52007, 24.70492, 24.88968, 
    25.07435, 25.25893, 25.44341, 25.62781, 25.81211, 25.9963, 26.1804, 
    26.36439, 26.54828, 26.73206, 26.91573, 27.09928, 27.28272, 27.46605, 
    27.64926, 27.83234, 28.0153, 28.19814, 28.38085, 28.56343, 28.74588, 
    28.9282, 29.11038, 29.29242, 29.47433, 29.65609, 29.8377, 30.01918, 
    30.2005, 30.38168, 30.5627, 30.74357, 30.92429, 31.10484, 31.28524, 
    31.46548, 31.64555, 31.82546, 32.00521, 32.18478, 32.36419, 32.54342, 
    32.72247, 32.90136, 33.08006, 33.25858, 33.43693, 33.61509, 33.79307, 
    33.97086, 34.14846, 34.32587, 34.50309, 34.68013, 34.85696, 35.0336, 
    35.21004, 35.38628, 35.56232, 35.73816, 35.9138, 36.08923, 36.26445, 
    36.43947, 36.61427, 36.78887, 36.96325, 37.13742, 37.31137, 37.48511, 
    37.65862, 37.83192, 38.005, 38.17785, 38.35048, 38.52289, 38.69507, 
    38.86702, 39.03875, 39.21024, 39.3815, 39.55254, 39.72334, 39.8939, 
    40.06422, 40.23431, 40.40417, 40.57378, 40.74316, 40.91229, 41.08118, 
    41.24982, 41.41823, 41.58638, 41.7543, 41.92196, 42.08937, 42.25654, 
    42.42345, 42.59012, 42.75653, 42.92269, 43.0886, 43.25425, 43.41965, 
    43.58479, 43.74967, 43.9143, 44.07866, 44.24277, 44.40662, 44.57021, 
    44.73353, 44.8966, 45.05939, 45.22193, 45.3842, 45.54622, 45.70796, 
    45.86943, 46.03064, 46.19159, 46.35226, 46.51267, 46.67281, 46.83267, 
    46.99227, 47.1516, 47.31066, 47.46944, 47.62796, 47.7862, 47.94417, 
    48.10186,
  -25.61905, -25.48681, -25.35431, -25.22154, -25.08851, -24.95521, 
    -24.82164, -24.6878, -24.5537, -24.41932, -24.28468, -24.14976, 
    -24.01458, -23.87912, -23.74339, -23.6074, -23.47112, -23.33458, 
    -23.19777, -23.06068, -22.92332, -22.78568, -22.64777, -22.50959, 
    -22.37113, -22.2324, -22.09339, -21.95411, -21.81454, -21.67471, 
    -21.5346, -21.39421, -21.25354, -21.11259, -20.97137, -20.82987, 
    -20.68809, -20.54604, -20.4037, -20.26109, -20.11819, -19.97502, 
    -19.83157, -19.68784, -19.54383, -19.39954, -19.25497, -19.11012, 
    -18.96499, -18.81958, -18.67388, -18.52791, -18.38166, -18.23512, 
    -18.08831, -17.94121, -17.79383, -17.64617, -17.49823, -17.35001, 
    -17.20151, -17.05273, -16.90366, -16.75432, -16.60469, -16.45478, 
    -16.30459, -16.15412, -16.00337, -15.85233, -15.70102, -15.54943, 
    -15.39755, -15.2454, -15.09296, -14.94024, -14.78725, -14.63397, 
    -14.48041, -14.32658, -14.17246, -14.01807, -13.8634, -13.70844, 
    -13.55322, -13.39771, -13.24192, -13.08586, -12.92952, -12.7729, -12.616, 
    -12.45883, -12.30139, -12.14366, -11.98567, -11.82739, -11.66885, 
    -11.51003, -11.35093, -11.19157, -11.03193, -10.87201, -10.71183, 
    -10.55138, -10.39065, -10.22966, -10.06839, -9.906858, -9.745057, 
    -9.582987, -9.42065, -9.258048, -9.095179, -8.932045, -8.768646, 
    -8.604983, -8.441058, -8.27687, -8.11242, -7.947709, -7.782738, 
    -7.617508, -7.452019, -7.286272, -7.120268, -6.954008, -6.787493, 
    -6.620723, -6.453699, -6.286423, -6.118896, -5.951117, -5.783088, 
    -5.614811, -5.446285, -5.277513, -5.108495, -4.939232, -4.769725, 
    -4.599975, -4.429983, -4.259751, -4.089279, -3.918569, -3.747622, 
    -3.576438, -3.40502, -3.233368, -3.061483, -2.889367, -2.717021, 
    -2.544446, -2.371643, -2.198614, -2.02536, -1.851882, -1.678183, 
    -1.504262, -1.330121, -1.155762, -0.9811865, -0.8063954, -0.6313902, 
    -0.4561725, -0.2807437, -0.1051052, 0.07074143, 0.2467947, 0.4230531, 
    0.599515, 0.776179, 0.9530434, 1.130107, 1.307367, 1.484823, 1.662474, 
    1.840316, 2.01835, 2.196572, 2.374982, 2.553577, 2.732356, 2.911318, 
    3.090459, 3.26978, 3.449277, 3.62895, 3.808795, 3.988812, 4.168999, 
    4.349354, 4.529874, 4.710559, 4.891405, 5.072412, 5.253577, 5.434898, 
    5.616374, 5.798003, 5.979781, 6.161708, 6.343782, 6.526, 6.708361, 
    6.890862, 7.073502, 7.256277, 7.439187, 7.62223, 7.805401, 7.988702, 
    8.172128, 8.355678, 8.539349, 8.723139, 8.907047, 9.09107, 9.275206, 
    9.459453, 9.643807, 9.828268, 10.01283, 10.1975, 10.38227, 10.56713, 
    10.75209, 10.93714, 11.12229, 11.30752, 11.49283, 11.67823, 11.86372, 
    12.04928, 12.23491, 12.42062, 12.60641, 12.79226, 12.97818, 13.16417, 
    13.35022, 13.53633, 13.72249, 13.90872, 14.09499, 14.28132, 14.46769, 
    14.65411, 14.84058, 15.02708, 15.21362, 15.4002, 15.58682, 15.77346, 
    15.96014, 16.14684, 16.33356, 16.52031, 16.70708, 16.89386, 17.08066, 
    17.26747, 17.45429, 17.64111, 17.82794, 18.01478, 18.20161, 18.38844, 
    18.57527, 18.76208, 18.94889, 19.13569, 19.32247, 19.50923, 19.69597, 
    19.8827, 20.06939, 20.25606, 20.4427, 20.62931, 20.81589, 21.00242, 
    21.18892, 21.37538, 21.56179, 21.74816, 21.93448, 22.12075, 22.30696, 
    22.49312, 22.67922, 22.86526, 23.05123, 23.23714, 23.42298, 23.60876, 
    23.79446, 23.98008, 24.16563, 24.3511, 24.53649, 24.72179, 24.90701, 
    25.09213, 25.27717, 25.46212, 25.64697, 25.83172, 26.01637, 26.20092, 
    26.38536, 26.5697, 26.75393, 26.93805, 27.12205, 27.30594, 27.48971, 
    27.67336, 27.8569, 28.0403, 28.22358, 28.40673, 28.58975, 28.77264, 
    28.9554, 29.13802, 29.3205, 29.50283, 29.68503, 29.86708, 30.04898, 
    30.23074, 30.41234, 30.59379, 30.77509, 30.95623, 31.13721, 31.31803, 
    31.49869, 31.67919, 31.85951, 32.03967, 32.21967, 32.39948, 32.57913, 
    32.7586, 32.93789, 33.117, 33.29594, 33.47469, 33.65325, 33.83163, 
    34.00983, 34.18783, 34.36564, 34.54326, 34.72068, 34.89791, 35.07495, 
    35.25178, 35.42841, 35.60484, 35.78107, 35.95709, 36.1329, 36.30851, 
    36.4839, 36.65909, 36.83406, 37.00882, 37.18336, 37.35768, 37.53179, 
    37.70567, 37.87934, 38.05278, 38.226, 38.39899, 38.57176, 38.7443, 
    38.91661, 39.08869, 39.26054, 39.43215, 39.60353, 39.77468, 39.94559, 
    40.11626, 40.28669, 40.45689, 40.62684, 40.79655, 40.96602, 41.13525, 
    41.30423, 41.47296, 41.64145, 41.80968, 41.97767, 42.14541, 42.3129, 
    42.48014, 42.64712, 42.81385, 42.98032, 43.14655, 43.31251, 43.47821, 
    43.64366, 43.80885, 43.97378, 44.13845, 44.30286, 44.46701, 44.63089, 
    44.79451, 44.95787, 45.12096, 45.28379, 45.44635, 45.60864, 45.77067, 
    45.93243, 46.09392, 46.25514, 46.41609, 46.57677, 46.73719, 46.89733, 
    47.0572, 47.21679, 47.37612, 47.53517, 47.69394, 47.85245, 48.01068, 
    48.16863,
  -25.70299, -25.57064, -25.43802, -25.30514, -25.17198, -25.03856, 
    -24.90487, -24.77091, -24.63668, -24.50217, -24.3674, -24.23236, 
    -24.09705, -23.96146, -23.8256, -23.68947, -23.55306, -23.41638, 
    -23.27943, -23.1422, -23.0047, -22.86692, -22.72887, -22.59054, 
    -22.45194, -22.31306, -22.1739, -22.03446, -21.89475, -21.75476, 
    -21.61449, -21.47395, -21.33312, -21.19202, -21.05064, -20.90898, 
    -20.76703, -20.62481, -20.48231, -20.33953, -20.19647, -20.05313, 
    -19.9095, -19.7656, -19.62141, -19.47695, -19.3322, -19.18717, -19.04185, 
    -18.89626, -18.75038, -18.60422, -18.45778, -18.31106, -18.16405, 
    -18.01676, -17.86919, -17.72134, -17.5732, -17.42478, -17.27608, 
    -17.12709, -16.97782, -16.82827, -16.67844, -16.52832, -16.37792, 
    -16.22724, -16.07627, -15.92502, -15.77349, -15.62168, -15.46958, 
    -15.31721, -15.16455, -15.01161, -14.85838, -14.70488, -14.55109, 
    -14.39702, -14.24267, -14.08804, -13.93313, -13.77794, -13.62247, 
    -13.46672, -13.31069, -13.15438, -12.99779, -12.84092, -12.68378, 
    -12.52635, -12.36865, -12.21067, -12.05242, -11.89388, -11.73507, 
    -11.57599, -11.41663, -11.257, -11.09709, -10.9369, -10.77645, -10.61572, 
    -10.45472, -10.29344, -10.1319, -9.970085, -9.808, -9.645644, -9.483021, 
    -9.320128, -9.156969, -8.993543, -8.829849, -8.665891, -8.501667, 
    -8.337178, -8.172427, -8.007413, -7.842136, -7.676599, -7.510801, 
    -7.344743, -7.178427, -7.011853, -6.845021, -6.677933, -6.51059, 
    -6.342992, -6.175141, -6.007038, -5.838682, -5.670076, -5.50122, 
    -5.332115, -5.162763, -4.993164, -4.823319, -4.65323, -4.482897, 
    -4.312322, -4.141506, -3.970449, -3.799154, -3.62762, -3.45585, 
    -3.283844, -3.111604, -2.939131, -2.766427, -2.593491, -2.420327, 
    -2.246934, -2.073315, -1.89947, -1.725401, -1.55111, -1.376597, 
    -1.201865, -1.026913, -0.8517452, -0.6763613, -0.5007631, -0.3249523, 
    -0.1489302, 0.02730167, 0.2037418, 0.3803886, 0.5572405, 0.7342961, 
    0.9115537, 1.089012, 1.266669, 1.444523, 1.622572, 1.800815, 1.979251, 
    2.157877, 2.336692, 2.515694, 2.694882, 2.874253, 3.053806, 3.233539, 
    3.41345, 3.593538, 3.7738, 3.954236, 4.134842, 4.315618, 4.49656, 
    4.677668, 4.858939, 5.040372, 5.221965, 5.403715, 5.58562, 5.76768, 
    5.949891, 6.132252, 6.31476, 6.497415, 6.680212, 6.863152, 7.046231, 
    7.229447, 7.412798, 7.596283, 7.7799, 7.963645, 8.147516, 8.331513, 
    8.515632, 8.699872, 8.88423, 9.068704, 9.253291, 9.43799, 9.622799, 
    9.807714, 9.992736, 10.17786, 10.36308, 10.5484, 10.73382, 10.91933, 
    11.10494, 11.29063, 11.47641, 11.66227, 11.84822, 12.03424, 12.22034, 
    12.40652, 12.59277, 12.77909, 12.96548, 13.15193, 13.33844, 13.52502, 
    13.71166, 13.89835, 14.08509, 14.27189, 14.45874, 14.64563, 14.83256, 
    15.01954, 15.20655, 15.39361, 15.58069, 15.76781, 15.95496, 16.14213, 
    16.32933, 16.51655, 16.70379, 16.89105, 17.07832, 17.26561, 17.4529, 
    17.6402, 17.82751, 18.01481, 18.20212, 18.38943, 18.57673, 18.76402, 
    18.9513, 19.13857, 19.32583, 19.51306, 19.70028, 19.88748, 20.07465, 
    20.26179, 20.4489, 20.63598, 20.82303, 21.01004, 21.19701, 21.38394, 
    21.57082, 21.75766, 21.94445, 22.13119, 22.31787, 22.5045, 22.69106, 
    22.87757, 23.06401, 23.25039, 23.4367, 23.62294, 23.8091, 23.99519, 
    24.1812, 24.36714, 24.55299, 24.73875, 24.92443, 25.11002, 25.29551, 
    25.48092, 25.66622, 25.85143, 26.03654, 26.22154, 26.40644, 26.59123, 
    26.77592, 26.96049, 27.14494, 27.32928, 27.5135, 27.6976, 27.88158, 
    28.06543, 28.24916, 28.43275, 28.61621, 28.79954, 28.98274, 29.1658, 
    29.34871, 29.53149, 29.71412, 29.8966, 30.07894, 30.26113, 30.44316, 
    30.62505, 30.80677, 30.98834, 31.16975, 31.35099, 31.53207, 31.71299, 
    31.89374, 32.07432, 32.25473, 32.43496, 32.61502, 32.7949, 32.97461, 
    33.15413, 33.33347, 33.51263, 33.6916, 33.87039, 34.04899, 34.22739, 
    34.40561, 34.58363, 34.76145, 34.93907, 35.1165, 35.29372, 35.47075, 
    35.64757, 35.82418, 36.00059, 36.17679, 36.35278, 36.52855, 36.70412, 
    36.87947, 37.0546, 37.22952, 37.40422, 37.57869, 37.75295, 37.92698, 
    38.10079, 38.27438, 38.44773, 38.62086, 38.79376, 38.96643, 39.13887, 
    39.31107, 39.48304, 39.65477, 39.82627, 39.99752, 40.16854, 40.33932, 
    40.50986, 40.68015, 40.8502, 41.02001, 41.18957, 41.35888, 41.52795, 
    41.69676, 41.86533, 42.03365, 42.20171, 42.36952, 42.53708, 42.70438, 
    42.87143, 43.03822, 43.20475, 43.37103, 43.53704, 43.7028, 43.8683, 
    44.03353, 44.19851, 44.36322, 44.52766, 44.69184, 44.85576, 45.01941, 
    45.1828, 45.34591, 45.50876, 45.67134, 45.83366, 45.9957, 46.15747, 
    46.31897, 46.48021, 46.64116, 46.80185, 46.96226, 47.1224, 47.28226, 
    47.44186, 47.60117, 47.76021, 47.91898, 48.07747, 48.23568,
  -25.78721, -25.65475, -25.52201, -25.38901, -25.25573, -25.12219, 
    -24.98838, -24.85429, -24.71994, -24.58531, -24.45041, -24.31524, 
    -24.1798, -24.04408, -23.90809, -23.77182, -23.63528, -23.49847, 
    -23.36138, -23.22401, -23.08637, -22.94845, -22.81025, -22.67178, 
    -22.53303, -22.394, -22.2547, -22.11511, -21.97525, -21.8351, -21.69468, 
    -21.55398, -21.413, -21.27174, -21.1302, -20.98837, -20.84627, -20.70388, 
    -20.56121, -20.41827, -20.27503, -20.13152, -19.98773, -19.84365, 
    -19.69929, -19.55464, -19.40972, -19.26451, -19.11901, -18.97323, 
    -18.82717, -18.68083, -18.5342, -18.38729, -18.24009, -18.09261, 
    -17.94484, -17.79679, -17.64846, -17.49984, -17.35094, -17.20175, 
    -17.05228, -16.90252, -16.75248, -16.60215, -16.45154, -16.30065, 
    -16.14947, -15.998, -15.84626, -15.69422, -15.54191, -15.38931, 
    -15.23643, -15.08326, -14.92981, -14.77607, -14.62206, -14.46776, 
    -14.31317, -14.15831, -14.00316, -13.84773, -13.69201, -13.53602, 
    -13.37975, -13.22319, -13.06635, -12.90923, -12.75184, -12.59416, 
    -12.4362, -12.27797, -12.11945, -11.96066, -11.80159, -11.64224, 
    -11.48261, -11.32271, -11.16253, -11.00208, -10.84135, -10.68034, 
    -10.51906, -10.35751, -10.19569, -10.03359, -9.87122, -9.708579, 
    -9.545668, -9.382485, -9.219034, -9.055314, -8.891326, -8.72707, 
    -8.562548, -8.397758, -8.232704, -8.067386, -7.901803, -7.735958, 
    -7.56985, -7.403481, -7.236851, -7.069962, -6.902813, -6.735406, 
    -6.567742, -6.399822, -6.231647, -6.063217, -5.894534, -5.725597, 
    -5.55641, -5.386972, -5.217285, -5.047349, -4.877165, -4.706736, 
    -4.536061, -4.365141, -4.193979, -4.022575, -3.85093, -3.679045, 
    -3.506922, -3.334562, -3.161966, -2.989135, -2.81607, -2.642773, 
    -2.469245, -2.295487, -2.121501, -1.947288, -1.772849, -1.598186, 
    -1.423299, -1.248191, -1.072863, -0.8973165, -0.7215523, -0.5455723, 
    -0.3693779, -0.1929706, -0.01635195, 0.1604766, 0.3375134, 0.514757, 
    0.6922058, 0.8698581, 1.047713, 1.225767, 1.404021, 1.582471, 1.761117, 
    1.939957, 2.118989, 2.298211, 2.477622, 2.657219, 2.837002, 3.016968, 
    3.197115, 3.377442, 3.557947, 3.738628, 3.919483, 4.100511, 4.281709, 
    4.463076, 4.644609, 4.826308, 5.008169, 5.19019, 5.372371, 5.554709, 
    5.737202, 5.919847, 6.102643, 6.285589, 6.468681, 6.651918, 6.835298, 
    7.018819, 7.202477, 7.386273, 7.570203, 7.754265, 7.938457, 8.122777, 
    8.307223, 8.491793, 8.676483, 8.861293, 9.04622, 9.231262, 9.416416, 
    9.601681, 9.787053, 9.972532, 10.15811, 10.3438, 10.52958, 10.71546, 
    10.90143, 11.0875, 11.27365, 11.4599, 11.64622, 11.83263, 12.01912, 
    12.20569, 12.39234, 12.57905, 12.76584, 12.9527, 13.13962, 13.32661, 
    13.51366, 13.70076, 13.88793, 14.07514, 14.26241, 14.44973, 14.6371, 
    14.82451, 15.01196, 15.19945, 15.38697, 15.57454, 15.76213, 15.94975, 
    16.1374, 16.32508, 16.51278, 16.70049, 16.88823, 17.07598, 17.26374, 
    17.45151, 17.63928, 17.82707, 18.01485, 18.20264, 18.39042, 18.5782, 
    18.76596, 18.95372, 19.14147, 19.3292, 19.51692, 19.70461, 19.89228, 
    20.07993, 20.26755, 20.45514, 20.64269, 20.83021, 21.0177, 21.20514, 
    21.39254, 21.5799, 21.76721, 21.95447, 22.14168, 22.32884, 22.51593, 
    22.70297, 22.88995, 23.07686, 23.26371, 23.45049, 23.63719, 23.82383, 
    24.01038, 24.19686, 24.38326, 24.56957, 24.7558, 24.94194, 25.12799, 
    25.31395, 25.49981, 25.68558, 25.87125, 26.05681, 26.24228, 26.42763, 
    26.61288, 26.79802, 26.98304, 27.16795, 27.35274, 27.53741, 27.72196, 
    27.90639, 28.09069, 28.27486, 28.4589, 28.64281, 28.82658, 29.01022, 
    29.19372, 29.37708, 29.56029, 29.74336, 29.92628, 30.10905, 30.29168, 
    30.47414, 30.65646, 30.83861, 31.02061, 31.20244, 31.38412, 31.56562, 
    31.74697, 31.92814, 32.10913, 32.28996, 32.47062, 32.6511, 32.83139, 
    33.01151, 33.19145, 33.3712, 33.55077, 33.73015, 33.90934, 34.08834, 
    34.26715, 34.44577, 34.62419, 34.80241, 34.98043, 35.15826, 35.33588, 
    35.51329, 35.69051, 35.86751, 36.0443, 36.22089, 36.39726, 36.57343, 
    36.74937, 36.9251, 37.10061, 37.27591, 37.45098, 37.62583, 37.80046, 
    37.97486, 38.14904, 38.32299, 38.49671, 38.6702, 38.84346, 39.01649, 
    39.18928, 39.36184, 39.53416, 39.70625, 39.8781, 40.04971, 40.22107, 
    40.39219, 40.56308, 40.73371, 40.9041, 41.07425, 41.24414, 41.41379, 
    41.58319, 41.75234, 41.92123, 42.08988, 42.25827, 42.4264, 42.59428, 
    42.76191, 42.92927, 43.09638, 43.26323, 43.42982, 43.59614, 43.76221, 
    43.92801, 44.09356, 44.25883, 44.42384, 44.58859, 44.75307, 44.91728, 
    45.08123, 45.24491, 45.40832, 45.57146, 45.73433, 45.89692, 46.05925, 
    46.2213, 46.38309, 46.54459, 46.70583, 46.86679, 47.02748, 47.18789, 
    47.34802, 47.50788, 47.66746, 47.82677, 47.98579, 48.14454, 48.30301,
  -25.87171, -25.73913, -25.60628, -25.47316, -25.33977, -25.2061, -25.07217, 
    -24.93796, -24.80348, -24.66873, -24.5337, -24.39841, -24.26283, 
    -24.12698, -23.99086, -23.85446, -23.71779, -23.58084, -23.44361, 
    -23.3061, -23.16832, -23.03026, -22.89192, -22.75331, -22.61441, 
    -22.47523, -22.33578, -22.19605, -22.05603, -21.91574, -21.77516, 
    -21.6343, -21.49317, -21.35175, -21.21004, -21.06806, -20.92579, 
    -20.78324, -20.64041, -20.49729, -20.35389, -20.21021, -20.06624, 
    -19.92199, -19.77745, -19.63263, -19.48753, -19.34214, -19.19646, 
    -19.0505, -18.90426, -18.75773, -18.61091, -18.46381, -18.31642, 
    -18.16875, -18.02079, -17.87254, -17.72401, -17.57519, -17.42609, 
    -17.2767, -17.12702, -16.97706, -16.82681, -16.67628, -16.52546, 
    -16.37435, -16.22296, -16.07128, -15.91931, -15.76706, -15.61453, 
    -15.4617, -15.3086, -15.1552, -15.00153, -14.84756, -14.69331, -14.53878, 
    -14.38396, -14.22886, -14.07347, -13.9178, -13.76185, -13.60561, 
    -13.44909, -13.29229, -13.1352, -12.97784, -12.82019, -12.66225, 
    -12.50404, -12.34555, -12.18677, -12.02772, -11.86838, -11.70877, 
    -11.54888, -11.38871, -11.22826, -11.06753, -10.90653, -10.74525, 
    -10.58369, -10.42186, -10.25976, -10.09737, -9.93472, -9.771792, 
    -9.608592, -9.44512, -9.281376, -9.117362, -8.953078, -8.788525, 
    -8.623702, -8.458612, -8.293255, -8.127631, -7.961741, -7.795588, 
    -7.629169, -7.462487, -7.295543, -7.128337, -6.960871, -6.793144, 
    -6.625159, -6.456915, -6.288414, -6.119658, -5.950645, -5.781378, 
    -5.611858, -5.442086, -5.272062, -5.101788, -4.931265, -4.760494, 
    -4.589475, -4.418211, -4.246701, -4.074948, -3.902953, -3.730716, 
    -3.558239, -3.385522, -3.212568, -3.039378, -2.865952, -2.692292, 
    -2.518399, -2.344275, -2.169921, -1.995338, -1.820527, -1.645491, 
    -1.470229, -1.294745, -1.119038, -0.9431112, -0.7669653, -0.5906019, 
    -0.4140224, -0.2372283, -0.06022129, 0.1169972, 0.2944257, 0.4720626, 
    0.6499062, 0.827955, 1.006207, 1.184662, 1.363316, 1.54217, 1.72122, 
    1.900465, 2.079905, 2.259536, 2.439357, 2.619366, 2.799562, 2.979943, 
    3.160506, 3.341251, 3.522175, 3.703277, 3.884554, 4.066005, 4.247628, 
    4.429421, 4.611382, 4.793509, 4.9758, 5.158253, 5.340867, 5.523638, 
    5.706566, 5.889648, 6.072883, 6.256267, 6.439799, 6.623478, 6.8073, 
    6.991264, 7.175368, 7.35961, 7.543987, 7.728497, 7.913138, 8.097909, 
    8.282806, 8.467828, 8.652972, 8.838237, 9.023619, 9.209117, 9.394729, 
    9.580452, 9.766283, 9.952222, 10.13826, 10.32441, 10.51065, 10.697, 
    10.88343, 11.06997, 11.25659, 11.44329, 11.63009, 11.81697, 12.00393, 
    12.19097, 12.37808, 12.56527, 12.75253, 12.93986, 13.12725, 13.31471, 
    13.50223, 13.68981, 13.87745, 14.06514, 14.25289, 14.44068, 14.62852, 
    14.81641, 15.00434, 15.1923, 15.38031, 15.56835, 15.75642, 15.94452, 
    16.13265, 16.3208, 16.50898, 16.69717, 16.88539, 17.07362, 17.26186, 
    17.45011, 17.63836, 17.82663, 18.01489, 18.20316, 18.39142, 18.57967, 
    18.76792, 18.95616, 19.14439, 19.3326, 19.52079, 19.70896, 19.89711, 
    20.08524, 20.27333, 20.4614, 20.64944, 20.83743, 21.02539, 21.21332, 
    21.4012, 21.58903, 21.77682, 21.96455, 22.15224, 22.33986, 22.52744, 
    22.71495, 22.9024, 23.08978, 23.2771, 23.46435, 23.65152, 23.83863, 
    24.02565, 24.2126, 24.39946, 24.58624, 24.77294, 24.95955, 25.14606, 
    25.33249, 25.51881, 25.70504, 25.89117, 26.0772, 26.26312, 26.44893, 
    26.63464, 26.82023, 27.00571, 27.19108, 27.37632, 27.56145, 27.74645, 
    27.93133, 28.11608, 28.3007, 28.48519, 28.66954, 28.85376, 29.03785, 
    29.22179, 29.40559, 29.58924, 29.77275, 29.95611, 30.13932, 30.32238, 
    30.50528, 30.68803, 30.87062, 31.05305, 31.23531, 31.41741, 31.59935, 
    31.78111, 31.96271, 32.14413, 32.32538, 32.50645, 32.68735, 32.86807, 
    33.0486, 33.22895, 33.40912, 33.5891, 33.76889, 33.94849, 34.1279, 
    34.30712, 34.48613, 34.66496, 34.84358, 35.022, 35.20022, 35.37824, 
    35.55605, 35.73365, 35.91105, 36.08823, 36.26521, 36.44197, 36.61852, 
    36.79484, 36.97095, 37.14685, 37.32252, 37.49797, 37.67319, 37.84819, 
    38.02297, 38.19752, 38.37183, 38.54592, 38.71978, 38.8934, 39.06679, 
    39.23994, 39.41286, 39.58554, 39.75798, 39.93018, 40.10213, 40.27385, 
    40.44532, 40.61654, 40.78753, 40.95826, 41.12874, 41.29897, 41.46896, 
    41.63869, 41.80817, 41.9774, 42.14637, 42.31509, 42.48355, 42.65175, 
    42.81969, 42.98738, 43.1548, 43.32197, 43.48887, 43.65551, 43.82189, 
    43.988, 44.15385, 44.31943, 44.48475, 44.64979, 44.81457, 44.97908, 
    45.14333, 45.3073, 45.471, 45.63443, 45.79758, 45.96047, 46.12308, 
    46.28542, 46.44748, 46.60927, 46.77078, 46.93201, 47.09298, 47.25366, 
    47.41406, 47.57419, 47.73404, 47.89361, 48.0529, 48.21191, 48.37064,
  -25.95649, -25.8238, -25.69083, -25.55759, -25.42408, -25.2903, -25.15624, 
    -25.02191, -24.88731, -24.75243, -24.61728, -24.48185, -24.34615, 
    -24.21017, -24.07392, -23.93739, -23.80058, -23.66349, -23.52613, 
    -23.38848, -23.25056, -23.11236, -22.97388, -22.83512, -22.69608, 
    -22.55676, -22.41716, -22.27727, -22.13711, -21.99666, -21.85593, 
    -21.71492, -21.57362, -21.43204, -21.29018, -21.14804, -21.00561, 
    -20.86289, -20.7199, -20.57661, -20.43304, -20.28919, -20.14505, 
    -20.00063, -19.85592, -19.71092, -19.56564, -19.42007, -19.27421, 
    -19.12807, -18.98164, -18.83492, -18.68792, -18.54063, -18.39305, 
    -18.24518, -18.09703, -17.94859, -17.79986, -17.65084, -17.50154, 
    -17.35195, -17.20207, -17.0519, -16.90145, -16.7507, -16.59967, 
    -16.44835, -16.29674, -16.14485, -15.99267, -15.8402, -15.68744, 
    -15.5344, -15.38106, -15.22744, -15.07354, -14.91935, -14.76487, 
    -14.6101, -14.45505, -14.29971, -14.14408, -13.98817, -13.83198, 
    -13.6755, -13.51873, -13.36168, -13.20435, -13.04673, -12.88883, 
    -12.73064, -12.57217, -12.41342, -12.25438, -12.09507, -11.93547, 
    -11.77559, -11.61543, -11.45499, -11.29427, -11.13327, -10.972, 
    -10.81044, -10.64861, -10.48649, -10.32411, -10.16144, -9.998502, 
    -9.835287, -9.671798, -9.508034, -9.343998, -9.179688, -9.015108, 
    -8.850256, -8.685133, -8.519741, -8.354079, -8.18815, -8.021953, 
    -7.855489, -7.688759, -7.521764, -7.354505, -7.186982, -7.019197, 
    -6.851149, -6.682841, -6.514273, -6.345446, -6.176361, -6.007019, 
    -5.83742, -5.667566, -5.497458, -5.327097, -5.156485, -4.98562, 
    -4.814506, -4.643143, -4.471532, -4.299675, -4.127572, -3.955224, 
    -3.782634, -3.609801, -3.436728, -3.263415, -3.089863, -2.916075, 
    -2.742051, -2.567792, -2.3933, -2.218576, -2.043622, -1.868438, 
    -1.693027, -1.517389, -1.341526, -1.16544, -0.9891313, -0.8126021, 
    -0.6358537, -0.4588876, -0.2817052, -0.1043082, 0.07330192, 0.2511236, 
    0.4291554, 0.6073955, 0.7858425, 0.9644946, 1.14335, 1.322408, 1.501666, 
    1.681122, 1.860775, 2.040623, 2.220665, 2.400898, 2.581321, 2.761932, 
    2.942729, 3.123711, 3.304876, 3.486221, 3.667745, 3.849446, 4.031322, 
    4.213372, 4.395593, 4.577983, 4.760541, 4.943264, 5.126151, 5.309199, 
    5.492407, 5.675772, 5.859293, 6.042967, 6.226793, 6.410768, 6.59489, 
    6.779157, 6.963567, 7.148118, 7.332807, 7.517633, 7.702594, 7.887687, 
    8.07291, 8.258261, 8.443738, 8.629337, 8.815059, 9.000899, 9.186855, 
    9.372927, 9.559111, 9.745404, 9.931805, 10.11831, 10.30492, 10.49163, 
    10.67844, 10.86534, 11.05234, 11.23943, 11.42661, 11.61387, 11.80122, 
    11.98865, 12.17616, 12.36375, 12.55141, 12.73914, 12.92694, 13.11481, 
    13.30275, 13.49075, 13.6788, 13.86692, 14.05509, 14.24331, 14.43158, 
    14.6199, 14.80826, 14.99667, 15.18512, 15.3736, 15.56212, 15.75068, 
    15.93926, 16.12787, 16.3165, 16.50516, 16.69384, 16.88253, 17.07124, 
    17.25997, 17.4487, 17.63744, 17.82618, 18.01493, 18.20367, 18.39242, 
    18.58116, 18.76989, 18.95861, 19.14732, 19.33601, 19.52468, 19.71334, 
    19.90197, 20.09057, 20.27915, 20.4677, 20.65621, 20.84469, 21.03313, 
    21.22153, 21.40989, 21.5982, 21.78647, 21.97468, 22.16284, 22.35095, 
    22.539, 22.72698, 22.91491, 23.10277, 23.29056, 23.47828, 23.66593, 
    23.85351, 24.041, 24.22842, 24.41576, 24.60301, 24.79017, 24.97725, 
    25.16423, 25.35112, 25.53791, 25.72461, 25.9112, 26.09769, 26.28407, 
    26.47035, 26.65651, 26.84257, 27.02851, 27.21433, 27.40003, 27.58561, 
    27.77107, 27.9564, 28.1416, 28.32667, 28.51161, 28.69642, 28.88108, 
    29.06561, 29.25, 29.43425, 29.61834, 29.8023, 29.9861, 30.16975, 
    30.35324, 30.53658, 30.71977, 30.90279, 31.08565, 31.26835, 31.45088, 
    31.63324, 31.81544, 31.99746, 32.17931, 32.36098, 32.54248, 32.72379, 
    32.90493, 33.08588, 33.26665, 33.44723, 33.62762, 33.80783, 33.98784, 
    34.16766, 34.34728, 34.5267, 34.70593, 34.88496, 35.06378, 35.2424, 
    35.42081, 35.59902, 35.77702, 35.95481, 36.13239, 36.30975, 36.4869, 
    36.66383, 36.84054, 37.01704, 37.19331, 37.36936, 37.54519, 37.72079, 
    37.89616, 38.07131, 38.24623, 38.42092, 38.59537, 38.76959, 38.94358, 
    39.11733, 39.29085, 39.46412, 39.63716, 39.80995, 39.9825, 40.15481, 
    40.32688, 40.4987, 40.67027, 40.84159, 41.01266, 41.18349, 41.35406, 
    41.52438, 41.69445, 41.86427, 42.03382, 42.20312, 42.37217, 42.54095, 
    42.70948, 42.87775, 43.04575, 43.2135, 43.38098, 43.5482, 43.71515, 
    43.88184, 44.04826, 44.21442, 44.3803, 44.54592, 44.71127, 44.87635, 
    45.04116, 45.2057, 45.36996, 45.53396, 45.69768, 45.86112, 46.0243, 
    46.18719, 46.34981, 46.51216, 46.67422, 46.83601, 46.99752, 47.15876, 
    47.31971, 47.48039, 47.64079, 47.8009, 47.96074, 48.12029, 48.27956, 
    48.43855,
  -26.04155, -25.90874, -25.77566, -25.64231, -25.50868, -25.37477, -25.2406, 
    -25.10615, -24.97142, -24.83642, -24.70115, -24.56559, -24.42976, 
    -24.29365, -24.15727, -24.0206, -23.88366, -23.74644, -23.60894, 
    -23.47116, -23.3331, -23.19476, -23.05613, -22.91723, -22.77804, 
    -22.63858, -22.49883, -22.35879, -22.21848, -22.07788, -21.93699, 
    -21.79583, -21.65438, -21.51264, -21.37062, -21.22831, -21.08572, 
    -20.94284, -20.79968, -20.65623, -20.51249, -20.36847, -20.22416, 
    -20.07956, -19.93468, -19.7895, -19.64404, -19.49829, -19.35226, 
    -19.20593, -19.05932, -18.91242, -18.76522, -18.61774, -18.46998, 
    -18.32192, -18.17357, -18.02493, -17.87601, -17.72679, -17.57729, 
    -17.42749, -17.27741, -17.12704, -16.97638, -16.82542, -16.67418, 
    -16.52265, -16.37083, -16.21872, -16.06632, -15.91363, -15.76065, 
    -15.60738, -15.45383, -15.29998, -15.14585, -14.99143, -14.83671, 
    -14.68172, -14.52643, -14.37085, -14.21499, -14.05884, -13.9024, 
    -13.74568, -13.58867, -13.43137, -13.27378, -13.11591, -12.95776, 
    -12.79932, -12.64059, -12.48158, -12.32229, -12.16271, -12.00285, 
    -11.8427, -11.68228, -11.52157, -11.36058, -11.1993, -11.03775, 
    -10.87592, -10.71381, -10.55141, -10.38874, -10.22579, -10.06257, 
    -9.899065, -9.735286, -9.571231, -9.4069, -9.242296, -9.077417, 
    -8.912267, -8.746843, -8.581148, -8.415181, -8.248945, -8.082439, 
    -7.915665, -7.748623, -7.581314, -7.413738, -7.245897, -7.077792, 
    -6.909423, -6.740792, -6.571898, -6.402744, -6.23333, -6.063656, 
    -5.893725, -5.723536, -5.553092, -5.382393, -5.21144, -5.040233, 
    -4.868775, -4.697066, -4.525108, -4.352901, -4.180447, -4.007747, 
    -3.834801, -3.661612, -3.48818, -3.314507, -3.140593, -2.966441, 
    -2.792051, -2.617425, -2.442564, -2.267469, -2.092142, -1.916584, 
    -1.740796, -1.564781, -1.388538, -1.21207, -1.035379, -0.8584647, 
    -0.6813298, -0.5039755, -0.3264032, -0.1486147, 0.02938871, 0.2076053, 
    0.3860336, 0.5646719, 0.7435187, 0.9225722, 1.101831, 1.281293, 1.460957, 
    1.640821, 1.820884, 2.001143, 2.181597, 2.362244, 2.543082, 2.724111, 
    2.905327, 3.086728, 3.268314, 3.450083, 3.632031, 3.814158, 3.996462, 
    4.17894, 4.361591, 4.544413, 4.727403, 4.910561, 5.093883, 5.277368, 
    5.461014, 5.644818, 5.82878, 6.012896, 6.197165, 6.381584, 6.566152, 
    6.750866, 6.935724, 7.120724, 7.305864, 7.491142, 7.676556, 7.862102, 
    8.04778, 8.233587, 8.41952, 8.605578, 8.791759, 8.978059, 9.164476, 
    9.35101, 9.537657, 9.724414, 9.91128, 10.09825, 10.28533, 10.4725, 
    10.65978, 10.84715, 11.03462, 11.22218, 11.40983, 11.59757, 11.78539, 
    11.97329, 12.16128, 12.34934, 12.53747, 12.72568, 12.91396, 13.10231, 
    13.29072, 13.4792, 13.66773, 13.85633, 14.04498, 14.23368, 14.42243, 
    14.61123, 14.80008, 14.98897, 15.1779, 15.36687, 15.55587, 15.7449, 
    15.93397, 16.12306, 16.31218, 16.50132, 16.69049, 16.87966, 17.06886, 
    17.25806, 17.44728, 17.63651, 17.82574, 18.01497, 18.2042, 18.39343, 
    18.58265, 18.77187, 18.96107, 19.15026, 19.33944, 19.5286, 19.71774, 
    19.90685, 20.09594, 20.285, 20.47403, 20.66303, 20.85199, 21.04091, 
    21.2298, 21.41863, 21.60743, 21.79617, 21.98487, 22.17351, 22.36209, 
    22.55062, 22.73908, 22.92749, 23.11582, 23.30409, 23.49229, 23.68042, 
    23.86847, 24.05644, 24.24433, 24.43214, 24.61986, 24.80749, 24.99504, 
    25.18249, 25.36985, 25.55711, 25.74427, 25.93133, 26.11829, 26.30514, 
    26.49187, 26.6785, 26.86502, 27.05142, 27.2377, 27.42386, 27.6099, 
    27.79581, 27.9816, 28.16726, 28.35278, 28.53818, 28.72343, 28.90855, 
    29.09353, 29.27836, 29.46305, 29.6476, 29.83199, 30.01624, 30.20033, 
    30.38427, 30.56805, 30.75167, 30.93513, 31.11842, 31.30155, 31.48452, 
    31.66731, 31.84994, 32.03239, 32.21466, 32.39676, 32.57868, 32.76042, 
    32.94198, 33.12335, 33.30454, 33.48553, 33.66634, 33.84696, 34.02739, 
    34.20761, 34.38764, 34.56747, 34.74711, 34.92654, 35.10577, 35.28479, 
    35.4636, 35.6422, 35.8206, 35.99878, 36.17675, 36.35451, 36.53204, 
    36.70937, 36.88646, 37.06334, 37.24, 37.41643, 37.59264, 37.76862, 
    37.94437, 38.11989, 38.29518, 38.47024, 38.64507, 38.81965, 38.994, 
    39.16812, 39.342, 39.51563, 39.68902, 39.86217, 40.03508, 40.20774, 
    40.38016, 40.55233, 40.72424, 40.89591, 41.06733, 41.2385, 41.40941, 
    41.58007, 41.75047, 41.92062, 42.09051, 42.26015, 42.42952, 42.59863, 
    42.76748, 42.93607, 43.1044, 43.27246, 43.44026, 43.6078, 43.77506, 
    43.94206, 44.1088, 44.27526, 44.44145, 44.60738, 44.77303, 44.93841, 
    45.10352, 45.26835, 45.43291, 45.5972, 45.76121, 45.92495, 46.08841, 
    46.25159, 46.41449, 46.57712, 46.73947, 46.90154, 47.06332, 47.22483, 
    47.38606, 47.54701, 47.70767, 47.86805, 48.02815, 48.18797, 48.3475, 
    48.50675,
  -26.1269, -25.99397, -25.86078, -25.72731, -25.59356, -25.45954, -25.32524, 
    -25.19067, -25.05582, -24.9207, -24.7853, -24.64962, -24.51366, 
    -24.37742, -24.2409, -24.10411, -23.96703, -23.82968, -23.69204, 
    -23.55412, -23.41592, -23.27744, -23.13868, -22.99963, -22.8603, 
    -22.72069, -22.58079, -22.44061, -22.30014, -22.15939, -22.01835, 
    -21.87703, -21.73543, -21.59353, -21.45135, -21.30889, -21.16613, 
    -21.02309, -20.87976, -20.73614, -20.59224, -20.44805, -20.30356, 
    -20.15879, -20.01373, -19.86839, -19.72275, -19.57682, -19.4306, 
    -19.28409, -19.1373, -18.99021, -18.84283, -18.69516, -18.5472, 
    -18.39895, -18.25041, -18.10158, -17.95246, -17.80304, -17.65334, 
    -17.50334, -17.35305, -17.20247, -17.05161, -16.90044, -16.74899, 
    -16.59725, -16.44521, -16.29289, -16.14027, -15.98736, -15.83416, 
    -15.68067, -15.52689, -15.37282, -15.21846, -15.06381, -14.90886, 
    -14.75363, -14.59811, -14.4423, -14.28619, -14.1298, -13.97312, 
    -13.81615, -13.6589, -13.50135, -13.34352, -13.1854, -13.02699, 
    -12.86829, -12.70931, -12.55004, -12.39048, -12.23064, -12.07052, 
    -11.91011, -11.74941, -11.58843, -11.42717, -11.26562, -11.1038, 
    -10.94169, -10.77929, -10.61662, -10.45367, -10.29043, -10.12692, 
    -9.963129, -9.799059, -9.634711, -9.470087, -9.305186, -9.14001, 
    -8.974559, -8.808833, -8.642835, -8.476562, -8.310019, -8.143204, 
    -7.976118, -7.808763, -7.641138, -7.473246, -7.305086, -7.13666, 
    -6.967969, -6.799013, -6.629793, -6.46031, -6.290566, -6.120561, 
    -5.950295, -5.779771, -5.608989, -5.437951, -5.266656, -5.095106, 
    -4.923303, -4.751247, -4.57894, -4.406383, -4.233576, -4.060522, 
    -3.88722, -3.713673, -3.539881, -3.365846, -3.19157, -3.017052, 
    -2.842295, -2.6673, -2.492069, -2.316602, -2.1409, -1.964966, -1.788801, 
    -1.612406, -1.435782, -1.258932, -1.081855, -0.9045551, -0.7270321, 
    -0.549288, -0.3713243, -0.1931425, -0.01474429, 0.1638689, 0.3426953, 
    0.5217335, 0.7009817, 0.8804384, 1.060102, 1.23997, 1.420042, 1.600316, 
    1.78079, 1.961462, 2.14233, 2.323393, 2.504649, 2.686096, 2.867732, 
    3.049556, 3.231565, 3.413758, 3.596133, 3.778688, 3.961421, 4.14433, 
    4.327413, 4.510668, 4.694093, 4.877687, 5.061447, 5.245371, 5.429457, 
    5.613703, 5.798108, 5.982668, 6.167382, 6.352248, 6.537263, 6.722426, 
    6.907735, 7.093187, 7.27878, 7.464511, 7.65038, 7.836382, 8.022517, 
    8.208782, 8.395175, 8.581694, 8.768335, 8.955097, 9.141979, 9.328977, 
    9.516088, 9.703312, 9.890645, 10.07808, 10.26563, 10.45328, 10.64102, 
    10.82887, 11.01681, 11.20484, 11.39296, 11.58117, 11.76947, 11.95785, 
    12.14631, 12.33485, 12.52347, 12.71215, 12.90091, 13.08974, 13.27863, 
    13.46759, 13.65661, 13.84568, 14.03481, 14.224, 14.41323, 14.60252, 
    14.79185, 14.98122, 15.17064, 15.36009, 15.54958, 15.7391, 15.92865, 
    16.11823, 16.30783, 16.49746, 16.68711, 16.87678, 17.06646, 17.25615, 
    17.44586, 17.63557, 17.82529, 18.01501, 18.20472, 18.39444, 18.58415, 
    18.77385, 18.96354, 19.15322, 19.34289, 19.53253, 19.72216, 19.91176, 
    20.10134, 20.29088, 20.4804, 20.66988, 20.85933, 21.04874, 21.2381, 
    21.42743, 21.6167, 21.80593, 21.99511, 22.18423, 22.3733, 22.56231, 
    22.75125, 22.94013, 23.12895, 23.3177, 23.50637, 23.69498, 23.8835, 
    24.07195, 24.26032, 24.4486, 24.6368, 24.82491, 25.01293, 25.20085, 
    25.38868, 25.57641, 25.76404, 25.95157, 26.139, 26.32631, 26.51352, 
    26.70061, 26.88759, 27.07445, 27.2612, 27.44782, 27.63432, 27.82069, 
    28.00694, 28.19305, 28.37903, 28.56488, 28.75059, 28.93616, 29.12159, 
    29.30687, 29.49201, 29.67701, 29.86185, 30.04654, 30.23107, 30.41545, 
    30.59967, 30.78373, 30.96763, 31.15137, 31.33493, 31.51833, 31.70156, 
    31.88461, 32.0675, 32.2502, 32.43273, 32.61507, 32.79724, 32.97922, 
    33.16101, 33.34262, 33.52404, 33.70526, 33.8863, 34.06713, 34.24777, 
    34.42822, 34.60846, 34.78849, 34.96833, 35.14796, 35.32738, 35.5066, 
    35.68561, 35.8644, 36.04298, 36.22134, 36.39949, 36.57742, 36.75513, 
    36.93262, 37.10988, 37.28692, 37.46374, 37.64032, 37.81668, 37.99281, 
    38.16871, 38.34437, 38.5198, 38.695, 38.86995, 39.04467, 39.21915, 
    39.39339, 39.56739, 39.74114, 39.91465, 40.08791, 40.26093, 40.4337, 
    40.60621, 40.77848, 40.9505, 41.12226, 41.29377, 41.46502, 41.63602, 
    41.80676, 41.97725, 42.14747, 42.31743, 42.48714, 42.65658, 42.82576, 
    42.99467, 43.16332, 43.3317, 43.49982, 43.66767, 43.83525, 44.00257, 
    44.16961, 44.33638, 44.50288, 44.66911, 44.83507, 45.00075, 45.16616, 
    45.33129, 45.49615, 45.66073, 45.82503, 45.98906, 46.15281, 46.31627, 
    46.47946, 46.64237, 46.805, 46.96735, 47.12941, 47.29119, 47.4527, 
    47.61391, 47.77485, 47.9355, 48.09587, 48.25595, 48.41574, 48.57525,
  -26.21253, -26.07949, -25.94618, -25.8126, -25.67873, -25.54459, -25.41018, 
    -25.27548, -25.14051, -25.00527, -24.86974, -24.73393, -24.59785, 
    -24.46148, -24.32483, -24.18791, -24.0507, -23.91321, -23.77544, 
    -23.63738, -23.49904, -23.36042, -23.22152, -23.08233, -22.94285, 
    -22.80309, -22.66305, -22.52272, -22.3821, -22.2412, -22.10001, 
    -21.95854, -21.81677, -21.67472, -21.53238, -21.38976, -21.24684, 
    -21.10364, -20.96014, -20.81636, -20.67229, -20.52792, -20.38327, 
    -20.23833, -20.09309, -19.94757, -19.80175, -19.65565, -19.50925, 
    -19.36256, -19.21558, -19.0683, -18.92074, -18.77288, -18.62473, 
    -18.47629, -18.32755, -18.17853, -18.02921, -17.87959, -17.72969, 
    -17.57949, -17.429, -17.27822, -17.12714, -16.97577, -16.8241, -16.67215, 
    -16.5199, -16.36736, -16.21452, -16.0614, -15.90797, -15.75426, 
    -15.60026, -15.44596, -15.29137, -15.13649, -14.98131, -14.82585, 
    -14.67009, -14.51404, -14.3577, -14.20107, -14.04414, -13.88693, 
    -13.72943, -13.57163, -13.41355, -13.25517, -13.09651, -12.93756, 
    -12.77832, -12.61879, -12.45898, -12.29887, -12.13848, -11.97781, 
    -11.81684, -11.65559, -11.49406, -11.33224, -11.17013, -11.00774, 
    -10.84507, -10.68212, -10.51888, -10.35536, -10.19156, -10.02748, 
    -9.863119, -9.698479, -9.533559, -9.368361, -9.202887, -9.037135, 
    -8.871107, -8.704803, -8.538225, -8.371373, -8.204247, -8.03685, 
    -7.86918, -7.70124, -7.53303, -7.364551, -7.195803, -7.026788, -6.857506, 
    -6.687959, -6.518147, -6.348072, -6.177733, -6.007133, -5.836272, 
    -5.665152, -5.493772, -5.322135, -5.150241, -4.978092, -4.805688, 
    -4.633031, -4.460122, -4.286962, -4.113551, -3.939893, -3.765986, 
    -3.591833, -3.417436, -3.242794, -3.06791, -2.892785, -2.71742, 
    -2.541816, -2.365976, -2.189899, -2.013587, -1.837043, -1.660267, 
    -1.483261, -1.306026, -1.128563, -0.9508752, -0.7729625, -0.5948271, 
    -0.4164703, -0.2378937, -0.05909901, 0.1199123, 0.2991386, 0.4785783, 
    0.6582298, 0.8380913, 1.018161, 1.198438, 1.37892, 1.559605, 1.740491, 
    1.921578, 2.102862, 2.284343, 2.466018, 2.647886, 2.829945, 3.012192, 
    3.194627, 3.377247, 3.56005, 3.743034, 3.926198, 4.10954, 4.293057, 
    4.476748, 4.66061, 4.844642, 5.028841, 5.213207, 5.397735, 5.582425, 
    5.767274, 5.952281, 6.137443, 6.322758, 6.508223, 6.693838, 6.879599, 
    7.065504, 7.251552, 7.437739, 7.624065, 7.810526, 7.99712, 8.183846, 
    8.370701, 8.557681, 8.744787, 8.932014, 9.119361, 9.306826, 9.494405, 
    9.682097, 9.8699, 10.05781, 10.24583, 10.43395, 10.62217, 10.81048, 
    10.9989, 11.18741, 11.37601, 11.56469, 11.75347, 11.94233, 12.13127, 
    12.32029, 12.50938, 12.69855, 12.88779, 13.0771, 13.26648, 13.45592, 
    13.64542, 13.83498, 14.0246, 14.21427, 14.40399, 14.59376, 14.78358, 
    14.97344, 15.16334, 15.35328, 15.54325, 15.73326, 15.9233, 16.11337, 
    16.30347, 16.49358, 16.68372, 16.87388, 17.06405, 17.25423, 17.44443, 
    17.63463, 17.82483, 18.01504, 18.20525, 18.39546, 18.58566, 18.77585, 
    18.96603, 19.1562, 19.34636, 19.53649, 19.7266, 19.9167, 20.10676, 
    20.29679, 20.4868, 20.67677, 20.8667, 21.0566, 21.24645, 21.43626, 
    21.62603, 21.81574, 22.0054, 22.19501, 22.38456, 22.57405, 22.76348, 
    22.95285, 23.14215, 23.33138, 23.52053, 23.70962, 23.89862, 24.08755, 
    24.2764, 24.46516, 24.65383, 24.84242, 25.03091, 25.21931, 25.40761, 
    25.59582, 25.78392, 25.97192, 26.15981, 26.3476, 26.53527, 26.72284, 
    26.91028, 27.09761, 27.28482, 27.4719, 27.65886, 27.8457, 28.0324, 
    28.21898, 28.40542, 28.59172, 28.77789, 28.96391, 29.1498, 29.33553, 
    29.52112, 29.70657, 29.89186, 30.07699, 30.26198, 30.4468, 30.63147, 
    30.81597, 31.00031, 31.18448, 31.36848, 31.55232, 31.73598, 31.91947, 
    32.10279, 32.28592, 32.46888, 32.65165, 32.83424, 33.01665, 33.19887, 
    33.38089, 33.56273, 33.74438, 33.92583, 34.10708, 34.28814, 34.46899, 
    34.64964, 34.83009, 35.01034, 35.19037, 35.3702, 35.54982, 35.72923, 
    35.90842, 36.08739, 36.26616, 36.4447, 36.62302, 36.80112, 36.979, 
    37.15665, 37.33408, 37.51128, 37.68824, 37.86499, 38.04149, 38.21777, 
    38.39381, 38.56961, 38.74517, 38.9205, 39.09559, 39.27044, 39.44504, 
    39.6194, 39.79351, 39.96738, 40.141, 40.31437, 40.48749, 40.66036, 
    40.83298, 41.00534, 41.17745, 41.3493, 41.5209, 41.69224, 41.86332, 
    42.03414, 42.2047, 42.37499, 42.54502, 42.7148, 42.8843, 43.05354, 
    43.22252, 43.39122, 43.55965, 43.72783, 43.89572, 44.06335, 44.2307, 
    44.39779, 44.56459, 44.73113, 44.89739, 45.06337, 45.22908, 45.39451, 
    45.55967, 45.72454, 45.88914, 46.05346, 46.21749, 46.38124, 46.54472, 
    46.70791, 46.87082, 47.03345, 47.19579, 47.35785, 47.51963, 47.68112, 
    47.84232, 48.00324, 48.16387, 48.32422, 48.48428, 48.64405,
  -26.29845, -26.1653, -26.03187, -25.89817, -25.76419, -25.62994, -25.4954, 
    -25.36059, -25.2255, -25.09012, -24.95447, -24.81854, -24.68233, 
    -24.54583, -24.40906, -24.272, -24.13466, -23.99703, -23.85913, 
    -23.72093, -23.58246, -23.4437, -23.30465, -23.16532, -23.0257, -22.8858, 
    -22.74561, -22.60513, -22.46437, -22.32331, -22.18197, -22.04034, 
    -21.89842, -21.75621, -21.61371, -21.47093, -21.32785, -21.18448, 
    -21.04082, -20.89688, -20.75263, -20.6081, -20.46328, -20.31816, 
    -20.17275, -20.02706, -19.88106, -19.73478, -19.5882, -19.44133, 
    -19.29416, -19.1467, -18.99895, -18.8509, -18.70256, -18.55393, -18.405, 
    -18.25578, -18.10626, -17.95645, -17.80634, -17.65594, -17.50525, 
    -17.35426, -17.20297, -17.0514, -16.89952, -16.74735, -16.59489, 
    -16.44213, -16.28908, -16.13573, -15.98209, -15.82816, -15.67393, 
    -15.5194, -15.36458, -15.20947, -15.05406, -14.89836, -14.74237, 
    -14.58608, -14.4295, -14.27263, -14.11546, -13.95801, -13.80026, 
    -13.64221, -13.48388, -13.32525, -13.16634, -13.00713, -12.84763, 
    -12.68785, -12.52777, -12.3674, -12.20675, -12.0458, -11.88457, 
    -11.72305, -11.56124, -11.39915, -11.23676, -11.0741, -10.91115, 
    -10.74791, -10.58439, -10.42058, -10.25649, -10.09212, -9.927469, 
    -9.762535, -9.59732, -9.431825, -9.26605, -9.099997, -8.933665, 
    -8.767056, -8.600171, -8.43301, -8.265574, -8.097862, -7.929878, 
    -7.761621, -7.593092, -7.424292, -7.255222, -7.085883, -6.916275, 
    -6.746399, -6.576257, -6.405849, -6.235177, -6.064241, -5.893042, 
    -5.721581, -5.54986, -5.37788, -5.205641, -5.033144, -4.860391, 
    -4.687383, -4.514121, -4.340605, -4.166838, -3.992821, -3.818554, 
    -3.644039, -3.469277, -3.29427, -3.119018, -2.943523, -2.767786, 
    -2.591809, -2.415593, -2.23914, -2.062449, -1.885525, -1.708366, 
    -1.530976, -1.353355, -1.175505, -0.9974269, -0.8191231, -0.6405947, 
    -0.4618432, -0.2828702, -0.1036774, 0.07573377, 0.2553616, 0.4352046, 
    0.6152609, 0.7955291, 0.9760072, 1.156694, 1.337587, 1.518685, 1.699987, 
    1.881489, 2.063192, 2.245092, 2.427188, 2.609479, 2.791962, 2.974635, 
    3.157497, 3.340546, 3.523779, 3.707196, 3.890793, 4.074569, 4.258523, 
    4.442651, 4.626952, 4.811425, 4.996066, 5.180874, 5.365847, 5.550983, 
    5.736279, 5.921734, 6.107346, 6.293111, 6.47903, 6.665097, 6.851313, 
    7.037674, 7.224179, 7.410825, 7.59761, 7.784532, 7.971589, 8.158777, 
    8.346095, 8.533542, 8.721113, 8.908808, 9.096622, 9.284556, 9.472606, 
    9.660769, 9.849043, 10.03743, 10.22592, 10.41451, 10.60321, 10.792, 
    10.98089, 11.16988, 11.35896, 11.54813, 11.73738, 11.92672, 12.11614, 
    12.30564, 12.49522, 12.68487, 12.8746, 13.06439, 13.25425, 13.44418, 
    13.63417, 13.82422, 14.01432, 14.20448, 14.39469, 14.58495, 14.77526, 
    14.96561, 15.156, 15.34643, 15.53689, 15.7274, 15.91793, 16.10849, 
    16.29907, 16.48968, 16.68031, 16.87096, 17.06162, 17.2523, 17.44299, 
    17.63368, 17.82438, 18.01508, 18.20578, 18.39648, 18.58718, 18.77786, 
    18.96854, 19.1592, 19.34984, 19.54047, 19.73108, 19.92166, 20.11222, 
    20.30274, 20.49324, 20.6837, 20.87412, 21.06451, 21.25485, 21.44515, 
    21.6354, 21.8256, 22.01575, 22.20585, 22.39589, 22.58587, 22.77578, 
    22.96563, 23.15542, 23.34513, 23.53477, 23.72434, 23.91383, 24.10324, 
    24.29256, 24.4818, 24.67096, 24.86002, 25.04899, 25.23787, 25.42665, 
    25.61533, 25.80391, 25.99238, 26.18075, 26.369, 26.55715, 26.74518, 
    26.93309, 27.12089, 27.30857, 27.49612, 27.68354, 27.87084, 28.05801, 
    28.24504, 28.43195, 28.61871, 28.80533, 28.99181, 29.17815, 29.36435, 
    29.55039, 29.73628, 29.92203, 30.10761, 30.29304, 30.47831, 30.66342, 
    30.84837, 31.03315, 31.21777, 31.40221, 31.58649, 31.77059, 31.95451, 
    32.13826, 32.32183, 32.50522, 32.68842, 32.87144, 33.05427, 33.23692, 
    33.41937, 33.60163, 33.7837, 33.96556, 34.14724, 34.3287, 34.50998, 
    34.69104, 34.8719, 35.05256, 35.233, 35.41323, 35.59326, 35.77307, 
    35.95266, 36.13204, 36.3112, 36.49014, 36.66885, 36.84734, 37.02561, 
    37.20365, 37.38147, 37.55905, 37.7364, 37.91353, 38.09042, 38.26707, 
    38.44349, 38.61966, 38.7956, 38.9713, 39.14676, 39.32197, 39.49694, 
    39.67166, 39.84614, 40.02036, 40.19434, 40.36807, 40.54155, 40.71477, 
    40.88773, 41.06045, 41.2329, 41.4051, 41.57704, 41.74872, 41.92014, 
    42.0913, 42.26219, 42.43282, 42.60319, 42.77329, 42.94312, 43.11269, 
    43.28198, 43.45101, 43.61977, 43.78825, 43.95647, 44.12441, 44.29208, 
    44.45947, 44.62659, 44.79343, 44.96, 45.12628, 45.29229, 45.45802, 
    45.62347, 45.78864, 45.95353, 46.11814, 46.28247, 46.44651, 46.61027, 
    46.77375, 46.93694, 47.09985, 47.26247, 47.4248, 47.58685, 47.74862, 
    47.91009, 48.07128, 48.23218, 48.39279, 48.55311, 48.71314,
  -26.38466, -26.25139, -26.11786, -25.98404, -25.84994, -25.71557, 
    -25.58092, -25.44598, -25.31077, -25.17528, -25.0395, -24.90344, 
    -24.7671, -24.63048, -24.49358, -24.35639, -24.21891, -24.08116, 
    -23.94311, -23.80479, -23.66617, -23.52727, -23.38809, -23.24861, 
    -23.10885, -22.9688, -22.82846, -22.68784, -22.54692, -22.40572, 
    -22.26423, -22.12244, -21.98037, -21.83801, -21.69535, -21.5524, 
    -21.40916, -21.26563, -21.12181, -20.9777, -20.83329, -20.68859, 
    -20.54359, -20.3983, -20.25272, -20.10685, -19.96068, -19.81421, 
    -19.66745, -19.5204, -19.37305, -19.22541, -19.07747, -18.92923, 
    -18.7807, -18.63188, -18.48276, -18.33334, -18.18362, -18.03361, 
    -17.88331, -17.7327, -17.58181, -17.43061, -17.27912, -17.12733, 
    -16.97525, -16.82286, -16.67019, -16.51721, -16.36394, -16.21038, 
    -16.05651, -15.90236, -15.7479, -15.59315, -15.4381, -15.28276, 
    -15.12712, -14.97119, -14.81496, -14.65843, -14.50161, -14.3445, 
    -14.18709, -14.02939, -13.87139, -13.7131, -13.55451, -13.39564, 
    -13.23647, -13.077, -12.91725, -12.7572, -12.59686, -12.43623, -12.27531, 
    -12.11409, -11.95259, -11.7908, -11.62872, -11.46635, -11.30369, 
    -11.14075, -10.97751, -10.81399, -10.65019, -10.48609, -10.32172, 
    -10.15706, -9.992111, -9.826882, -9.661371, -9.495577, -9.329502, 
    -9.163147, -8.996511, -8.829597, -8.662403, -8.494932, -8.327184, 
    -8.159159, -7.990859, -7.822284, -7.653436, -7.484314, -7.31492, 
    -7.145256, -6.97532, -6.805115, -6.634642, -6.463901, -6.292893, 
    -6.121621, -5.950083, -5.778282, -5.606217, -5.433892, -5.261306, 
    -5.088461, -4.915358, -4.741997, -4.568381, -4.39451, -4.220385, 
    -4.046007, -3.871379, -3.6965, -3.521373, -3.345998, -3.170377, 
    -2.994511, -2.818401, -2.64205, -2.465457, -2.288625, -2.111554, 
    -1.934247, -1.756705, -1.578929, -1.400921, -1.222681, -1.044212, 
    -0.8655158, -0.6865929, -0.5074451, -0.3280741, -0.1484814, 0.03133126, 
    0.2113624, 0.3916102, 0.5720732, 0.7527497, 0.9336379, 1.114736, 
    1.296043, 1.477556, 1.659274, 1.841195, 2.023317, 2.205639, 2.388158, 
    2.570873, 2.753782, 2.936883, 3.120175, 3.303654, 3.48732, 3.67117, 
    3.855203, 4.039416, 4.223807, 4.408375, 4.593118, 4.778032, 4.963118, 
    5.148371, 5.333791, 5.519374, 5.70512, 5.891026, 6.077089, 6.263309, 
    6.449681, 6.636205, 6.822877, 7.009697, 7.196661, 7.383768, 7.571015, 
    7.758399, 7.94592, 8.133574, 8.321359, 8.509272, 8.697312, 8.885476, 
    9.073762, 9.262167, 9.450688, 9.639325, 9.828074, 10.01693, 10.2059, 
    10.39497, 10.58414, 10.77342, 10.96279, 11.15226, 11.34182, 11.53147, 
    11.7212, 11.91103, 12.10093, 12.29092, 12.48098, 12.67112, 12.86133, 
    13.05162, 13.24197, 13.43238, 13.62286, 13.8134, 14.00399, 14.19464, 
    14.38534, 14.57609, 14.76689, 14.95773, 15.14862, 15.33954, 15.5305, 
    15.7215, 15.91252, 16.10357, 16.29466, 16.48576, 16.67689, 16.86803, 
    17.05919, 17.25036, 17.44154, 17.63273, 17.82393, 18.01512, 18.20632, 
    18.39751, 18.5887, 18.77988, 18.97105, 19.16221, 19.35335, 19.54447, 
    19.73557, 19.92665, 20.1177, 20.30872, 20.49971, 20.69066, 20.88158, 
    21.07246, 21.26329, 21.45408, 21.64483, 21.83552, 22.02616, 22.21675, 
    22.40728, 22.59774, 22.78815, 22.97849, 23.16876, 23.35896, 23.54909, 
    23.73914, 23.92911, 24.11901, 24.30882, 24.49854, 24.68818, 24.87772, 
    25.06717, 25.25653, 25.44579, 25.63494, 25.824, 26.01295, 26.20179, 
    26.39052, 26.57914, 26.76764, 26.95603, 27.1443, 27.33244, 27.52046, 
    27.70835, 27.89612, 28.08375, 28.27125, 28.45861, 28.64584, 28.83292, 
    29.01987, 29.20666, 29.39331, 29.57981, 29.76616, 29.95235, 30.13839, 
    30.32427, 30.50999, 30.69555, 30.88094, 31.06617, 31.25123, 31.43612, 
    31.62083, 31.80537, 31.98974, 32.17392, 32.35793, 32.54174, 32.72538, 
    32.90883, 33.09209, 33.27517, 33.45804, 33.64073, 33.82322, 34.0055, 
    34.1876, 34.36948, 34.55117, 34.73265, 34.91393, 35.09499, 35.27584, 
    35.45649, 35.63692, 35.81713, 35.99713, 36.17691, 36.35646, 36.5358, 
    36.71491, 36.8938, 37.07246, 37.25089, 37.42909, 37.60707, 37.78481, 
    37.96231, 38.13958, 38.31661, 38.49341, 38.66996, 38.84628, 39.02235, 
    39.19817, 39.37376, 39.54909, 39.72418, 39.89902, 40.07361, 40.24794, 
    40.42203, 40.59586, 40.76944, 40.94276, 41.11582, 41.28862, 41.46117, 
    41.63345, 41.80547, 41.97723, 42.14873, 42.31996, 42.49093, 42.66162, 
    42.83206, 43.00222, 43.17211, 43.34173, 43.51109, 43.68016, 43.84897, 
    44.0175, 44.18576, 44.35374, 44.52144, 44.68887, 44.85602, 45.02289, 
    45.18948, 45.35579, 45.52182, 45.68757, 45.85304, 46.01822, 46.18312, 
    46.34774, 46.51207, 46.67612, 46.83988, 47.00335, 47.16654, 47.32944, 
    47.49205, 47.65438, 47.81641, 47.97816, 48.13961, 48.30078, 48.46166, 
    48.62224, 48.78254,
  -26.47115, -26.33778, -26.20413, -26.0702, -25.93599, -25.8015, -25.66673, 
    -25.53167, -25.39634, -25.26072, -25.12482, -24.98864, -24.85217, 
    -24.71543, -24.57839, -24.44107, -24.30347, -24.16558, -24.0274, 
    -23.88894, -23.75019, -23.61115, -23.47182, -23.3322, -23.1923, 
    -23.05211, -22.91162, -22.77085, -22.62979, -22.48843, -22.34679, 
    -22.20485, -22.06262, -21.9201, -21.77729, -21.63418, -21.49078, 
    -21.34709, -21.2031, -21.05882, -20.91425, -20.76938, -20.62421, 
    -20.47875, -20.333, -20.18694, -20.0406, -19.89396, -19.74702, -19.59978, 
    -19.45225, -19.30442, -19.15629, -19.00787, -18.85915, -18.71013, 
    -18.56082, -18.41121, -18.26129, -18.11109, -17.96058, -17.80977, 
    -17.65867, -17.50727, -17.35557, -17.20358, -17.05128, -16.89869, 
    -16.74579, -16.5926, -16.43912, -16.28533, -16.13125, -15.97686, 
    -15.82218, -15.6672, -15.51193, -15.35636, -15.20049, -15.04432, 
    -14.88785, -14.73109, -14.57403, -14.41667, -14.25902, -14.10107, 
    -13.94283, -13.78429, -13.62545, -13.46632, -13.3069, -13.14718, 
    -12.98716, -12.82685, -12.66625, -12.50536, -12.34417, -12.18269, 
    -12.02092, -11.85885, -11.6965, -11.53385, -11.37092, -11.20769, 
    -11.04418, -10.88037, -10.71628, -10.5519, -10.38724, -10.22229, 
    -10.05705, -9.891523, -9.725715, -9.559622, -9.393246, -9.226587, 
    -9.059648, -8.892426, -8.724923, -8.557141, -8.38908, -8.220741, 
    -8.052124, -7.883231, -7.714062, -7.544618, -7.3749, -7.204908, 
    -7.034645, -6.86411, -6.693304, -6.522229, -6.350885, -6.179275, 
    -6.007397, -5.835253, -5.662846, -5.490174, -5.317241, -5.144046, 
    -4.970591, -4.796877, -4.622905, -4.448677, -4.274192, -4.099454, 
    -3.924462, -3.749219, -3.573725, -3.397981, -3.221989, -3.045751, 
    -2.869267, -2.692539, -2.515568, -2.338356, -2.160904, -1.983214, 
    -1.805286, -1.627123, -1.448725, -1.270095, -1.091234, -0.9121428, 
    -0.7328237, -0.5532779, -0.3735072, -0.1935131, -0.01329719, 0.1671388, 
    0.3477934, 0.5286648, 0.7097513, 0.8910513, 1.072563, 1.254285, 1.436215, 
    1.618351, 1.800692, 1.983236, 2.165981, 2.348926, 2.532067, 2.715404, 
    2.898935, 3.082658, 3.26657, 3.45067, 3.634956, 3.819426, 4.004078, 
    4.18891, 4.373919, 4.559105, 4.744464, 4.929996, 5.115696, 5.301565, 
    5.487599, 5.673796, 5.860155, 6.046672, 6.233347, 6.420176, 6.607158, 
    6.79429, 6.98157, 7.168996, 7.356566, 7.544277, 7.732127, 7.920114, 
    8.108235, 8.296489, 8.484872, 8.673383, 8.862019, 9.050777, 9.239656, 
    9.428654, 9.617766, 9.806993, 9.996329, 10.18577, 10.37533, 10.56498, 
    10.75473, 10.94459, 11.13454, 11.32458, 11.51472, 11.70494, 11.89525, 
    12.08564, 12.27612, 12.46667, 12.6573, 12.848, 13.03877, 13.22961, 
    13.42052, 13.61149, 13.80252, 13.9936, 14.18475, 14.37594, 14.56719, 
    14.75848, 14.94982, 15.1412, 15.33262, 15.52407, 15.71556, 15.90709, 
    16.09864, 16.29021, 16.48182, 16.67344, 16.86508, 17.05674, 17.24841, 
    17.44008, 17.63177, 17.82347, 18.01516, 18.20686, 18.39855, 18.59024, 
    18.78191, 18.97358, 19.16524, 19.35687, 19.54849, 19.74009, 19.93167, 
    20.12321, 20.31473, 20.50621, 20.69767, 20.88908, 21.08045, 21.27178, 
    21.46307, 21.65431, 21.84549, 22.03663, 22.22771, 22.41873, 22.60969, 
    22.80058, 22.99141, 23.18217, 23.37286, 23.56348, 23.75402, 23.94448, 
    24.13486, 24.32516, 24.51537, 24.70548, 24.89551, 25.08545, 25.27529, 
    25.46503, 25.65466, 25.8442, 26.03363, 26.22295, 26.41216, 26.60125, 
    26.79023, 26.97909, 27.16783, 27.35645, 27.54494, 27.7333, 27.92153, 
    28.10963, 28.2976, 28.48543, 28.67311, 28.86066, 29.04807, 29.23532, 
    29.42243, 29.60939, 29.79619, 29.98284, 30.16933, 30.35567, 30.54184, 
    30.72785, 30.91369, 31.09936, 31.28487, 31.4702, 31.65536, 31.84034, 
    32.02514, 32.20977, 32.39421, 32.57846, 32.76254, 32.94642, 33.13011, 
    33.31361, 33.49692, 33.68003, 33.86294, 34.04565, 34.22816, 34.41047, 
    34.59258, 34.77448, 34.95616, 35.13764, 35.31891, 35.49996, 35.6808, 
    35.86142, 36.04182, 36.222, 36.40196, 36.5817, 36.7612, 36.94049, 
    37.11954, 37.29837, 37.47696, 37.65532, 37.83345, 38.01134, 38.18899, 
    38.36641, 38.54358, 38.72051, 38.8972, 39.07365, 39.24984, 39.4258, 
    39.6015, 39.77695, 39.95216, 40.12711, 40.30181, 40.47625, 40.65044, 
    40.82437, 40.99805, 41.17146, 41.34461, 41.51751, 41.69014, 41.8625, 
    42.0346, 42.20644, 42.37801, 42.54931, 42.72034, 42.8911, 43.0616, 
    43.23182, 43.40176, 43.57144, 43.74084, 43.90997, 44.07882, 44.24739, 
    44.41568, 44.5837, 44.75144, 44.9189, 45.08607, 45.25297, 45.41958, 
    45.58591, 45.75196, 45.91772, 46.0832, 46.2484, 46.4133, 46.57793, 
    46.74226, 46.9063, 47.07006, 47.23353, 47.39671, 47.5596, 47.7222, 
    47.88451, 48.04653, 48.20825, 48.36969, 48.53083, 48.69168, 48.85223,
  -26.55794, -26.42446, -26.2907, -26.15665, -26.02233, -25.88772, -25.75283, 
    -25.61766, -25.4822, -25.34646, -25.21044, -25.07414, -24.93755, 
    -24.80067, -24.66351, -24.52606, -24.38832, -24.2503, -24.11199, 
    -23.97339, -23.8345, -23.69532, -23.55586, -23.4161, -23.27605, 
    -23.13572, -22.99509, -22.85417, -22.71296, -22.57145, -22.42966, 
    -22.28757, -22.14518, -22.00251, -21.85953, -21.71627, -21.57271, 
    -21.42885, -21.2847, -21.14025, -20.99551, -20.85048, -20.70514, 
    -20.55951, -20.41358, -20.26735, -20.12083, -19.97401, -19.82689, 
    -19.67947, -19.53176, -19.38374, -19.23543, -19.08682, -18.93791, 
    -18.7887, -18.63919, -18.48938, -18.33928, -18.18887, -18.03816, 
    -17.88716, -17.73585, -17.58424, -17.43234, -17.28013, -17.12762, 
    -16.97482, -16.82171, -16.66831, -16.5146, -16.36059, -16.20629, 
    -16.05168, -15.89678, -15.74157, -15.58607, -15.43026, -15.27416, 
    -15.11776, -14.96106, -14.80406, -14.64676, -14.48916, -14.33126, 
    -14.17307, -14.01458, -13.85579, -13.6967, -13.53732, -13.37764, 
    -13.21766, -13.05739, -12.89682, -12.73595, -12.57479, -12.41334, 
    -12.25159, -12.08955, -11.92721, -11.76458, -11.60166, -11.43845, 
    -11.27494, -11.11114, -10.94706, -10.78268, -10.61801, -10.45306, 
    -10.28781, -10.12228, -9.956459, -9.790353, -9.62396, -9.457283, 
    -9.290321, -9.123075, -8.955546, -8.787734, -8.61964, -8.451266, 
    -8.282611, -8.113677, -7.944464, -7.774974, -7.605206, -7.435163, 
    -7.264844, -7.094251, -6.923385, -6.752246, -6.580836, -6.409155, 
    -6.237205, -6.064986, -5.8925, -5.719747, -5.546729, -5.373446, 
    -5.199901, -5.026093, -4.852024, -4.677696, -4.503109, -4.328264, 
    -4.153163, -3.977807, -3.802197, -3.626335, -3.450221, -3.273858, 
    -3.097245, -2.920386, -2.74328, -2.56593, -2.388337, -2.210501, 
    -2.032426, -1.854111, -1.675559, -1.496771, -1.317749, -1.138493, 
    -0.9590061, -0.7792891, -0.5993438, -0.4191717, -0.2387744, -0.05815361, 
    0.1226891, 0.303752, 0.4850335, 0.6665319, 0.8482455, 1.030172, 1.212311, 
    1.39466, 1.577217, 1.75998, 1.942947, 2.126117, 2.309489, 2.493059, 
    2.676826, 2.860788, 3.044944, 3.229291, 3.413828, 3.598552, 3.783461, 
    3.968554, 4.153828, 4.339281, 4.524912, 4.710718, 4.896698, 5.082848, 
    5.269167, 5.455654, 5.642305, 5.829119, 6.016093, 6.203225, 6.390513, 
    6.577956, 6.765549, 6.953292, 7.141182, 7.329217, 7.517395, 7.705713, 
    7.894169, 8.08276, 8.271484, 8.46034, 8.649324, 8.838434, 9.027669, 
    9.217025, 9.406499, 9.59609, 9.785795, 9.975613, 10.16554, 10.35557, 
    10.54571, 10.73595, 10.92629, 11.11672, 11.30725, 11.49788, 11.68859, 
    11.87939, 12.07027, 12.26123, 12.45228, 12.64339, 12.83459, 13.02585, 
    13.21719, 13.40859, 13.60005, 13.79158, 13.98316, 14.1748, 14.36649, 
    14.55823, 14.75002, 14.94186, 15.13374, 15.32565, 15.51761, 15.7096, 
    15.90162, 16.09367, 16.28575, 16.47785, 16.66997, 16.86211, 17.05427, 
    17.24644, 17.43862, 17.63081, 17.82301, 18.0152, 18.2074, 18.39959, 
    18.59178, 18.78396, 18.97613, 19.16828, 19.36042, 19.55254, 19.74464, 
    19.93671, 20.12876, 20.32077, 20.51276, 20.70471, 20.89662, 21.08849, 
    21.28032, 21.4721, 21.66384, 21.85552, 22.04715, 22.23872, 22.43024, 
    22.62169, 22.81308, 23.00441, 23.19566, 23.38684, 23.57795, 23.76898, 
    23.95993, 24.1508, 24.34159, 24.53228, 24.72289, 24.91341, 25.10383, 
    25.29415, 25.48437, 25.67449, 25.86451, 26.05442, 26.24422, 26.43391, 
    26.62348, 26.81294, 27.00227, 27.19149, 27.38058, 27.56954, 27.75838, 
    27.94708, 28.13565, 28.32409, 28.51238, 28.70054, 28.88855, 29.07642, 
    29.26414, 29.4517, 29.63912, 29.82639, 30.01349, 30.20044, 30.38723, 
    30.57386, 30.76032, 30.94661, 31.13273, 31.31869, 31.50446, 31.69007, 
    31.87549, 32.06074, 32.2458, 32.43068, 32.61538, 32.79988, 32.9842, 
    33.16832, 33.35226, 33.53599, 33.71953, 33.90287, 34.08601, 34.26894, 
    34.45168, 34.6342, 34.81651, 34.99862, 35.18051, 35.36219, 35.54366, 
    35.7249, 35.90593, 36.08674, 36.26733, 36.44769, 36.62782, 36.80773, 
    36.98741, 37.16686, 37.34608, 37.52507, 37.70382, 37.88233, 38.06061, 
    38.23865, 38.41645, 38.594, 38.77131, 38.94838, 39.1252, 39.30177, 
    39.4781, 39.65417, 39.82999, 40.00556, 40.18088, 40.35594, 40.53074, 
    40.70529, 40.87958, 41.0536, 41.22737, 41.40088, 41.57412, 41.74709, 
    41.9198, 42.09225, 42.26442, 42.43633, 42.60797, 42.77934, 42.95043, 
    43.12125, 43.29181, 43.46208, 43.63208, 43.8018, 43.97125, 44.14042, 
    44.30931, 44.47792, 44.64625, 44.8143, 44.98206, 45.14955, 45.31675, 
    45.48367, 45.6503, 45.81665, 45.98271, 46.14848, 46.31397, 46.47917, 
    46.64408, 46.8087, 46.97303, 47.13707, 47.30082, 47.46428, 47.62745, 
    47.79033, 47.95291, 48.1152, 48.27719, 48.4389, 48.6003, 48.76142, 
    48.92224,
  -26.64503, -26.51143, -26.37756, -26.2434, -26.10896, -25.97424, -25.83923, 
    -25.70394, -25.56837, -25.43251, -25.29636, -25.15993, -25.02322, 
    -24.88621, -24.74892, -24.61134, -24.47348, -24.33532, -24.19688, 
    -24.05814, -23.91912, -23.77981, -23.6402, -23.5003, -23.36011, 
    -23.21963, -23.07886, -22.93779, -22.79643, -22.65478, -22.51283, 
    -22.37059, -22.22805, -22.08522, -21.94209, -21.79866, -21.65494, 
    -21.51093, -21.36661, -21.222, -21.07709, -20.93188, -20.78638, 
    -20.64058, -20.49447, -20.34807, -20.20137, -20.05437, -19.90708, 
    -19.75948, -19.61158, -19.46338, -19.31488, -19.16608, -19.01698, 
    -18.86758, -18.71788, -18.56787, -18.41757, -18.26696, -18.11606, 
    -17.96485, -17.81334, -17.66153, -17.50941, -17.357, -17.20428, 
    -17.05126, -16.89794, -16.74432, -16.5904, -16.43617, -16.28164, 
    -16.12681, -15.97168, -15.81625, -15.66052, -15.50448, -15.34815, 
    -15.19151, -15.03457, -14.87733, -14.71979, -14.56195, -14.40381, 
    -14.24537, -14.08663, -13.9276, -13.76826, -13.60862, -13.44868, 
    -13.28845, -13.12792, -12.96709, -12.80596, -12.64453, -12.48281, 
    -12.3208, -12.15848, -11.99587, -11.83297, -11.66977, -11.50628, 
    -11.34249, -11.17841, -11.01404, -10.84938, -10.68442, -10.51917, 
    -10.35364, -10.18781, -10.02169, -9.855289, -9.688597, -9.521617, 
    -9.35435, -9.186798, -9.01896, -8.850838, -8.682432, -8.513743, 
    -8.344772, -8.175519, -8.005986, -7.836174, -7.666082, -7.495712, 
    -7.325065, -7.154141, -6.982943, -6.81147, -6.639723, -6.467704, 
    -6.295414, -6.122853, -5.950023, -5.776924, -5.603558, -5.429925, 
    -5.256028, -5.081866, -4.907441, -4.732755, -4.557807, -4.382601, 
    -4.207137, -4.031415, -3.855438, -3.679206, -3.502721, -3.325984, 
    -3.148996, -2.97176, -2.794275, -2.616544, -2.438568, -2.260348, 
    -2.081886, -1.903183, -1.72424, -1.54506, -1.365644, -1.185992, 
    -1.006108, -0.8259912, -0.6456447, -0.4650695, -0.2842674, -0.10324, 
    0.07801108, 0.2594842, 0.4411776, 0.6230896, 0.8052185, 0.9875626, 
    1.17012, 1.352889, 1.535868, 1.719055, 1.902448, 2.086046, 2.269846, 
    2.453846, 2.638046, 2.822442, 3.007033, 3.191816, 3.376791, 3.561955, 
    3.747306, 3.932842, 4.11856, 4.30446, 4.490538, 4.676793, 4.863223, 
    5.049825, 5.236598, 5.423539, 5.610646, 5.797917, 5.98535, 6.172942, 
    6.360692, 6.548596, 6.736654, 6.924862, 7.113219, 7.301722, 7.490368, 
    7.679156, 7.868083, 8.057147, 8.246346, 8.435676, 8.625135, 8.814722, 
    9.004435, 9.194269, 9.384224, 9.574296, 9.764483, 9.954783, 10.14519, 
    10.33571, 10.52634, 10.71706, 10.90789, 11.09881, 11.28983, 11.48094, 
    11.67214, 11.86343, 12.05481, 12.24627, 12.4378, 12.62942, 12.82111, 
    13.01287, 13.2047, 13.39659, 13.58855, 13.78058, 13.97266, 14.16479, 
    14.35699, 14.54923, 14.74152, 14.93385, 15.12623, 15.31865, 15.51111, 
    15.7036, 15.89612, 16.08868, 16.28126, 16.47386, 16.66649, 16.85913, 
    17.05179, 17.24447, 17.43715, 17.62984, 17.82254, 18.01524, 18.20794, 
    18.40064, 18.59333, 18.78601, 18.97868, 19.17134, 19.36398, 19.55661, 
    19.74921, 19.94178, 20.13433, 20.32685, 20.51934, 20.71179, 20.9042, 
    21.09657, 21.2889, 21.48118, 21.67342, 21.8656, 22.05773, 22.2498, 
    22.44182, 22.63377, 22.82565, 23.01747, 23.20922, 23.4009, 23.5925, 
    23.78403, 23.97547, 24.16683, 24.35811, 24.54929, 24.74039, 24.9314, 
    25.1223, 25.31312, 25.50382, 25.69443, 25.88493, 26.07533, 26.26561, 
    26.45578, 26.64583, 26.83577, 27.02558, 27.21527, 27.40484, 27.59428, 
    27.78359, 27.97277, 28.16181, 28.35072, 28.53948, 28.72811, 28.91659, 
    29.10492, 29.2931, 29.48114, 29.66902, 29.85674, 30.04431, 30.23172, 
    30.41896, 30.60604, 30.79296, 30.9797, 31.16628, 31.35268, 31.53891, 
    31.72496, 31.91083, 32.09652, 32.28202, 32.46735, 32.65248, 32.83743, 
    33.02218, 33.20674, 33.39111, 33.57527, 33.75924, 33.94301, 34.12658, 
    34.30994, 34.49309, 34.67604, 34.85877, 35.04129, 35.22361, 35.4057, 
    35.58758, 35.76924, 35.95068, 36.13189, 36.31288, 36.49365, 36.67419, 
    36.8545, 37.03458, 37.21442, 37.39404, 37.57342, 37.75256, 37.93147, 
    38.11013, 38.28856, 38.46674, 38.64468, 38.82236, 38.99981, 39.17701, 
    39.35396, 39.53065, 39.7071, 39.88329, 40.05923, 40.23491, 40.41033, 
    40.5855, 40.76041, 40.93505, 41.10943, 41.28355, 41.45741, 41.631, 
    41.80432, 41.97738, 42.15017, 42.32269, 42.49493, 42.66691, 42.83861, 
    43.01004, 43.1812, 43.35208, 43.52268, 43.693, 43.86305, 44.03282, 
    44.20231, 44.37152, 44.54045, 44.70909, 44.87745, 45.04553, 45.21332, 
    45.38083, 45.54805, 45.71498, 45.88163, 46.04799, 46.21406, 46.37984, 
    46.54533, 46.71053, 46.87544, 47.04006, 47.20439, 47.36842, 47.53216, 
    47.69561, 47.85876, 48.02161, 48.18418, 48.34644, 48.50842, 48.67009, 
    48.83147, 48.99255,
  -26.73241, -26.5987, -26.46471, -26.33044, -26.19589, -26.06105, -25.92593, 
    -25.79052, -25.65483, -25.51885, -25.38258, -25.24603, -25.10919, 
    -24.97206, -24.83464, -24.69693, -24.55894, -24.42065, -24.28207, 
    -24.1432, -24.00404, -23.86459, -23.72485, -23.58481, -23.44448, 
    -23.30386, -23.16294, -23.02172, -22.88021, -22.73841, -22.59631, 
    -22.45392, -22.31123, -22.16824, -22.02495, -21.88137, -21.73749, 
    -21.59331, -21.44883, -21.30406, -21.15898, -21.01361, -20.86793, 
    -20.72196, -20.57568, -20.42911, -20.28223, -20.13505, -19.98757, 
    -19.83979, -19.69171, -19.54333, -19.39464, -19.24566, -19.09637, 
    -18.94677, -18.79688, -18.64668, -18.49618, -18.34538, -18.19427, 
    -18.04286, -17.89115, -17.73913, -17.58681, -17.43418, -17.28126, 
    -17.12802, -16.97449, -16.82065, -16.66651, -16.51206, -16.35731, 
    -16.20226, -16.0469, -15.89124, -15.73528, -15.57902, -15.42245, 
    -15.26557, -15.1084, -14.95092, -14.79314, -14.63506, -14.47668, 
    -14.31799, -14.159, -13.99971, -13.84012, -13.68023, -13.52004, 
    -13.35955, -13.19876, -13.03767, -12.87628, -12.71459, -12.5526, 
    -12.39031, -12.22773, -12.06484, -11.90166, -11.73819, -11.57442, 
    -11.41035, -11.24599, -11.08133, -10.91638, -10.75113, -10.58559, 
    -10.41976, -10.25364, -10.08723, -9.920526, -9.753531, -9.586248, 
    -9.418676, -9.250817, -9.08267, -8.914237, -8.745518, -8.576513, 
    -8.407226, -8.237654, -8.0678, -7.897663, -7.727246, -7.556549, 
    -7.385573, -7.214318, -7.042787, -6.870978, -6.698895, -6.526536, 
    -6.353905, -6.181, -6.007824, -5.834379, -5.660663, -5.48668, -5.312428, 
    -5.137912, -4.96313, -4.788085, -4.612776, -4.437207, -4.261377, 
    -4.085289, -3.908942, -3.73234, -3.555482, -3.37837, -3.201006, 
    -3.023391, -2.845526, -2.667412, -2.489052, -2.310446, -2.131595, 
    -1.952502, -1.773168, -1.593595, -1.413782, -1.233734, -1.05345, 
    -0.8729322, -0.6921827, -0.5112029, -0.3299942, -0.1485585, 0.03310277, 
    0.2149878, 0.3970949, 0.5794224, 0.7619684, 0.9447315, 1.12771, 1.310901, 
    1.494304, 1.677917, 1.861737, 2.045764, 2.229995, 2.414428, 2.599061, 
    2.783893, 2.968921, 3.154144, 3.339559, 3.525165, 3.710959, 3.89694, 
    4.083105, 4.269453, 4.455981, 4.642687, 4.829569, 5.016625, 5.203854, 
    5.391252, 5.578817, 5.766547, 5.954441, 6.142496, 6.330709, 6.519079, 
    6.707603, 6.896279, 7.085104, 7.274077, 7.463195, 7.652455, 7.841856, 
    8.031395, 8.221068, 8.410876, 8.600815, 8.790881, 8.981073, 9.17139, 
    9.361827, 9.552382, 9.743054, 9.93384, 10.12474, 10.31574, 10.50685, 
    10.69807, 10.88939, 11.0808, 11.27231, 11.46392, 11.65561, 11.84739, 
    12.03926, 12.23122, 12.42325, 12.61536, 12.80755, 12.99981, 13.19213, 
    13.38453, 13.57699, 13.76952, 13.9621, 14.15474, 14.34743, 14.54017, 
    14.73297, 14.92581, 15.11869, 15.31161, 15.50457, 15.69757, 15.8906, 
    16.08366, 16.27674, 16.46985, 16.66298, 16.85613, 17.0493, 17.24248, 
    17.43567, 17.62887, 17.82207, 18.01528, 18.20849, 18.40169, 18.59489, 
    18.78808, 18.98126, 19.17442, 19.36757, 19.5607, 19.7538, 19.94688, 
    20.13994, 20.33296, 20.52595, 20.71891, 20.91183, 21.1047, 21.29753, 
    21.49032, 21.68305, 21.87574, 22.06837, 22.26094, 22.45346, 22.64591, 
    22.83829, 23.03061, 23.22286, 23.41503, 23.60713, 23.79915, 23.99109, 
    24.18295, 24.37472, 24.5664, 24.75799, 24.94948, 25.14088, 25.33218, 
    25.52338, 25.71448, 25.90547, 26.09635, 26.28712, 26.47777, 26.6683, 
    26.85872, 27.04902, 27.23919, 27.42924, 27.61916, 27.80894, 27.9986, 
    28.18811, 28.37749, 28.56673, 28.75583, 28.94477, 29.13358, 29.32223, 
    29.51073, 29.69907, 29.88726, 30.07529, 30.26316, 30.45086, 30.6384, 
    30.82577, 31.01298, 31.2, 31.38686, 31.57354, 31.76004, 31.94636, 
    32.13249, 32.31844, 32.50421, 32.68979, 32.87517, 33.06036, 33.24536, 
    33.43016, 33.61476, 33.79916, 33.98336, 34.16735, 34.35114, 34.53472, 
    34.71809, 34.90125, 35.08419, 35.26692, 35.44943, 35.63173, 35.8138, 
    35.99565, 36.17727, 36.35867, 36.53984, 36.72079, 36.9015, 37.08198, 
    37.26223, 37.44224, 37.62202, 37.80155, 37.98085, 38.1599, 38.33871, 
    38.51728, 38.6956, 38.87368, 39.0515, 39.22908, 39.4064, 39.58347, 
    39.76029, 39.93686, 40.11316, 40.28921, 40.465, 40.64053, 40.81579, 
    40.9908, 41.16553, 41.34001, 41.51422, 41.68816, 41.86183, 42.03524, 
    42.20837, 42.38123, 42.55382, 42.72614, 42.89817, 43.06994, 43.24143, 
    43.41264, 43.58357, 43.75422, 43.92459, 44.09468, 44.2645, 44.43402, 
    44.60327, 44.77222, 44.9409, 45.10929, 45.27739, 45.4452, 45.61273, 
    45.77997, 45.94691, 46.11357, 46.27994, 46.44601, 46.6118, 46.77729, 
    46.94249, 47.1074, 47.272, 47.43632, 47.60034, 47.76406, 47.92749, 
    48.09063, 48.25346, 48.416, 48.57824, 48.74018, 48.90182, 49.06317,
  -26.82009, -26.68627, -26.55217, -26.41779, -26.28312, -26.14817, 
    -26.01293, -25.87741, -25.74159, -25.60549, -25.4691, -25.33243, 
    -25.19546, -25.05821, -24.92066, -24.78283, -24.6447, -24.50628, 
    -24.36757, -24.22857, -24.08928, -23.94969, -23.8098, -23.66963, 
    -23.52915, -23.38839, -23.24732, -23.10596, -22.96431, -22.82236, 
    -22.68011, -22.53756, -22.39472, -22.25157, -22.10813, -21.96439, 
    -21.82035, -21.67601, -21.53137, -21.38643, -21.24118, -21.09564, 
    -20.9498, -20.80365, -20.6572, -20.51045, -20.3634, -20.21605, -20.06839, 
    -19.92043, -19.77216, -19.6236, -19.47473, -19.32555, -19.17607, 
    -19.02629, -18.8762, -18.72581, -18.57511, -18.4241, -18.2728, -18.12119, 
    -17.96927, -17.81705, -17.66452, -17.51168, -17.35855, -17.2051, 
    -17.05135, -16.8973, -16.74294, -16.58827, -16.4333, -16.27802, 
    -16.12244, -15.96656, -15.81036, -15.65387, -15.49706, -15.33996, 
    -15.18255, -15.02483, -14.86681, -14.70848, -14.54986, -14.39092, 
    -14.23169, -14.07215, -13.91231, -13.75216, -13.59171, -13.43096, 
    -13.26991, -13.10856, -12.9469, -12.78495, -12.62269, -12.46013, 
    -12.29728, -12.13412, -11.97067, -11.80691, -11.64286, -11.47851, 
    -11.31387, -11.14892, -10.98368, -10.81815, -10.65232, -10.4862, 
    -10.31978, -10.15307, -9.986063, -9.818768, -9.65118, -9.483303, 
    -9.315135, -9.146679, -8.977933, -8.8089, -8.63958, -8.469974, -8.300082, 
    -8.129906, -7.959445, -7.788702, -7.617677, -7.446371, -7.274784, 
    -7.102918, -6.930773, -6.758351, -6.585652, -6.412678, -6.23943, 
    -6.065908, -5.892114, -5.718048, -5.543712, -5.369106, -5.194233, 
    -5.019093, -4.843687, -4.668016, -4.492083, -4.315887, -4.13943, 
    -3.962713, -3.785739, -3.608507, -3.431019, -3.253277, -3.075282, 
    -2.897035, -2.718537, -2.539791, -2.360797, -2.181557, -2.002073, 
    -1.822345, -1.642376, -1.462167, -1.281719, -1.101034, -0.9201141, 
    -0.73896, -0.5575737, -0.3759568, -0.194111, -0.0120379, 0.1702608, 
    0.3527834, 0.5355281, 0.7184932, 0.901677, 1.085078, 1.268693, 1.452522, 
    1.636563, 1.820813, 2.00527, 2.189934, 2.374801, 2.55987, 2.74514, 
    2.930608, 3.116271, 3.302129, 3.488179, 3.674419, 3.860847, 4.047461, 
    4.234259, 4.421238, 4.608398, 4.795735, 4.983248, 5.170933, 5.35879, 
    5.546816, 5.735009, 5.923366, 6.111885, 6.300565, 6.489402, 6.678394, 
    6.86754, 7.056837, 7.246282, 7.435874, 7.625609, 7.815486, 8.005502, 
    8.195655, 8.385942, 8.576361, 8.766909, 8.957584, 9.148384, 9.339307, 
    9.530349, 9.721508, 9.912782, 10.10417, 10.29566, 10.48727, 10.67897, 
    10.87078, 11.06269, 11.2547, 11.4468, 11.63899, 11.83127, 12.02363, 
    12.21608, 12.40862, 12.60123, 12.79391, 12.98667, 13.1795, 13.3724, 
    13.56537, 13.75839, 13.95148, 14.14462, 14.33782, 14.53107, 14.72437, 
    14.91771, 15.1111, 15.30453, 15.498, 15.6915, 15.88504, 16.07861, 
    16.2722, 16.46582, 16.65946, 16.85312, 17.04679, 17.24048, 17.43419, 
    17.62789, 17.82161, 18.01532, 18.20904, 18.40275, 18.59646, 18.79016, 
    18.98384, 19.17752, 19.37117, 19.56481, 19.75842, 19.95201, 20.14557, 
    20.33911, 20.5326, 20.72607, 20.91949, 21.11287, 21.30621, 21.4995, 
    21.69275, 21.88593, 22.07907, 22.27215, 22.46516, 22.65812, 22.851, 
    23.04382, 23.23657, 23.42924, 23.62184, 23.81436, 24.0068, 24.19915, 
    24.39142, 24.5836, 24.77568, 24.96767, 25.15957, 25.35136, 25.54305, 
    25.73464, 25.92612, 26.11748, 26.30874, 26.49988, 26.6909, 26.88181, 
    27.07259, 27.26324, 27.45377, 27.64417, 27.83443, 28.02456, 28.21456, 
    28.40441, 28.59413, 28.7837, 28.97312, 29.16239, 29.35151, 29.54048, 
    29.72929, 29.91795, 30.10644, 30.29477, 30.48294, 30.67094, 30.85877, 
    31.04642, 31.23391, 31.42122, 31.60835, 31.7953, 31.98207, 32.16866, 
    32.35505, 32.54126, 32.72728, 32.91311, 33.09874, 33.28418, 33.46942, 
    33.65446, 33.83929, 34.02392, 34.20835, 34.39256, 34.57657, 34.76036, 
    34.94395, 35.12732, 35.31046, 35.49339, 35.67611, 35.85859, 36.04086, 
    36.22289, 36.4047, 36.58628, 36.76763, 36.94875, 37.12963, 37.31028, 
    37.49069, 37.67086, 37.85079, 38.03048, 38.20993, 38.38913, 38.56808, 
    38.74679, 38.92525, 39.10345, 39.28141, 39.45911, 39.63656, 39.81375, 
    39.99068, 40.16736, 40.34378, 40.51993, 40.69582, 40.87145, 41.04681, 
    41.22191, 41.39674, 41.57131, 41.7456, 41.91962, 42.09338, 42.26685, 
    42.44006, 42.61299, 42.78564, 42.95802, 43.13012, 43.30194, 43.47349, 
    43.64475, 43.81573, 43.98643, 44.15685, 44.32698, 44.49682, 44.66638, 
    44.83566, 45.00465, 45.17334, 45.34175, 45.50988, 45.67771, 45.84525, 
    46.0125, 46.17946, 46.34612, 46.51249, 46.67857, 46.84435, 47.00984, 
    47.17503, 47.33993, 47.50453, 47.66883, 47.83284, 47.99654, 48.15995, 
    48.32306, 48.48587, 48.64838, 48.81059, 48.9725, 49.1341,
  -26.90806, -26.77414, -26.63993, -26.50543, -26.37065, -26.23559, 
    -26.10023, -25.96459, -25.82866, -25.69244, -25.55593, -25.41913, 
    -25.28205, -25.14466, -25.00699, -24.86903, -24.73077, -24.59223, 
    -24.45338, -24.31425, -24.17482, -24.03509, -23.89507, -23.75475, 
    -23.61414, -23.47323, -23.33202, -23.19052, -23.04872, -22.90661, 
    -22.76422, -22.62152, -22.47852, -22.33522, -22.19162, -22.04772, 
    -21.90352, -21.75902, -21.61422, -21.46911, -21.3237, -21.17799, 
    -21.03198, -20.88566, -20.73904, -20.59212, -20.44489, -20.29736, 
    -20.14952, -20.00138, -19.85293, -19.70418, -19.55512, -19.40576, 
    -19.25609, -19.10612, -18.95584, -18.80525, -18.65435, -18.50315, 
    -18.35165, -18.19983, -18.04771, -17.89528, -17.74255, -17.58951, 
    -17.43616, -17.2825, -17.12854, -16.97426, -16.81969, -16.6648, 
    -16.50961, -16.35411, -16.1983, -16.04218, -15.88576, -15.72904, -15.572, 
    -15.41466, -15.25701, -15.09906, -14.94079, -14.78223, -14.62335, 
    -14.46417, -14.30469, -14.1449, -13.98481, -13.82441, -13.6637, 
    -13.50269, -13.34138, -13.17976, -13.01785, -12.85562, -12.6931, 
    -12.53027, -12.36714, -12.20371, -12.03998, -11.87595, -11.71162, 
    -11.54699, -11.38206, -11.21683, -11.0513, -10.88547, -10.71935, 
    -10.55293, -10.38622, -10.21921, -10.05191, -9.884308, -9.716416, 
    -9.548232, -9.379756, -9.210988, -9.04193, -8.872582, -8.702945, 
    -8.53302, -8.362807, -8.192307, -8.021523, -7.850452, -7.679098, 
    -7.50746, -7.33554, -7.163339, -6.990857, -6.818096, -6.645056, 
    -6.471738, -6.298144, -6.124275, -5.950131, -5.775713, -5.601024, 
    -5.426063, -5.250833, -5.075333, -4.899565, -4.723531, -4.547232, 
    -4.370668, -4.193842, -4.016754, -3.839405, -3.661798, -3.483932, 
    -3.305811, -3.127434, -2.948804, -2.769921, -2.590788, -2.411405, 
    -2.231774, -2.051896, -1.871774, -1.691408, -1.5108, -1.329951, 
    -1.148864, -0.9675391, -0.7859787, -0.6041843, -0.4221574, -0.2398998, 
    -0.05741302, 0.1253011, 0.308241, 0.4914047, 0.6747907, 0.8583971, 
    1.042222, 1.226264, 1.410521, 1.594991, 1.779672, 1.964563, 2.149661, 
    2.334965, 2.520472, 2.706182, 2.892091, 3.078197, 3.264499, 3.450996, 
    3.637683, 3.824561, 4.011626, 4.198876, 4.38631, 4.573925, 4.761719, 
    4.94969, 5.137836, 5.326154, 5.514643, 5.7033, 5.892122, 6.081109, 
    6.270256, 6.459563, 6.649027, 6.838645, 7.028415, 7.218335, 7.408403, 
    7.598616, 7.788971, 7.979467, 8.1701, 8.360869, 8.551772, 8.742805, 
    8.933966, 9.125253, 9.316663, 9.508193, 9.699841, 9.891606, 10.08348, 
    10.27547, 10.46757, 10.65977, 10.85207, 11.04448, 11.23698, 11.42958, 
    11.62227, 11.81505, 12.00792, 12.20087, 12.3939, 12.58702, 12.7802, 
    12.97347, 13.1668, 13.36021, 13.55368, 13.74721, 13.9408, 14.13445, 
    14.32816, 14.52191, 14.71572, 14.90958, 15.10347, 15.29741, 15.49139, 
    15.68541, 15.87945, 16.07353, 16.26764, 16.46177, 16.65592, 16.85009, 
    17.04428, 17.23848, 17.43269, 17.62691, 17.82113, 18.01536, 18.20959, 
    18.40381, 18.59803, 18.79224, 18.98644, 19.18063, 19.3748, 19.56894, 
    19.76307, 19.95717, 20.15124, 20.34529, 20.5393, 20.73327, 20.9272, 
    21.12109, 21.31494, 21.50874, 21.70249, 21.89618, 22.08983, 22.28341, 
    22.47693, 22.67039, 22.86378, 23.05711, 23.25036, 23.44354, 23.63664, 
    23.82966, 24.0226, 24.21545, 24.40822, 24.60089, 24.79348, 24.98596, 
    25.17835, 25.37064, 25.56283, 25.7549, 25.94687, 26.13873, 26.33048, 
    26.52211, 26.71362, 26.90501, 27.09628, 27.28742, 27.47843, 27.66932, 
    27.86006, 28.05068, 28.24115, 28.43148, 28.62167, 28.81172, 29.00161, 
    29.19136, 29.38095, 29.57039, 29.75967, 29.9488, 30.13776, 30.32655, 
    30.51518, 30.70365, 30.89194, 31.08006, 31.268, 31.45576, 31.64335, 
    31.83076, 32.01798, 32.20501, 32.39186, 32.57852, 32.76498, 32.95126, 
    33.13733, 33.32321, 33.50888, 33.69436, 33.87963, 34.0647, 34.24955, 
    34.4342, 34.61864, 34.80286, 34.98687, 35.17066, 35.35423, 35.53758, 
    35.72071, 35.90362, 36.0863, 36.26875, 36.45097, 36.63296, 36.81471, 
    36.99624, 37.17752, 37.35857, 37.53939, 37.71996, 37.90028, 38.08037, 
    38.2602, 38.4398, 38.61914, 38.79823, 38.97708, 39.15567, 39.334, 
    39.51208, 39.68991, 39.86748, 40.04478, 40.22183, 40.39862, 40.57514, 
    40.7514, 40.92739, 41.10311, 41.27857, 41.45376, 41.62867, 41.80332, 
    41.9777, 42.1518, 42.32562, 42.49917, 42.67245, 42.84544, 43.01816, 
    43.1906, 43.36275, 43.53463, 43.70622, 43.87753, 44.04856, 44.2193, 
    44.38975, 44.55992, 44.7298, 44.89939, 45.06869, 45.23771, 45.40643, 
    45.57486, 45.74299, 45.91084, 46.07839, 46.24565, 46.41261, 46.57928, 
    46.74565, 46.91172, 47.0775, 47.24298, 47.40816, 47.57305, 47.73763, 
    47.90192, 48.0659, 48.22958, 48.39297, 48.55605, 48.71883, 48.88131, 
    49.04348, 49.20535,
  -26.99634, -26.86231, -26.72799, -26.59338, -26.45849, -26.32331, 
    -26.18784, -26.05208, -25.91603, -25.7797, -25.64307, -25.50615, 
    -25.36893, -25.23143, -25.09363, -24.95554, -24.81716, -24.67848, 
    -24.5395, -24.40023, -24.26067, -24.12081, -23.98065, -23.84019, 
    -23.69944, -23.55839, -23.41704, -23.27538, -23.13344, -22.99119, 
    -22.84864, -22.70579, -22.56264, -22.41918, -22.27543, -22.13137, 
    -21.98701, -21.84235, -21.69739, -21.55212, -21.40654, -21.26067, 
    -21.11448, -20.968, -20.8212, -20.6741, -20.5267, -20.37899, -20.23098, 
    -20.08265, -19.93402, -19.78509, -19.63585, -19.48629, -19.33644, 
    -19.18627, -19.0358, -18.88501, -18.73392, -18.58253, -18.43082, 
    -18.2788, -18.12648, -17.97384, -17.8209, -17.66765, -17.51409, 
    -17.36022, -17.20604, -17.05155, -16.89676, -16.74165, -16.58624, 
    -16.43051, -16.27448, -16.11814, -15.96149, -15.80453, -15.64726, 
    -15.48968, -15.3318, -15.1736, -15.0151, -14.85629, -14.69717, -14.53774, 
    -14.37801, -14.21797, -14.05762, -13.89697, -13.73601, -13.57474, 
    -13.41317, -13.25129, -13.08911, -12.92662, -12.76382, -12.60073, 
    -12.43732, -12.27362, -12.10961, -11.9453, -11.78069, -11.61577, 
    -11.45056, -11.28504, -11.11923, -10.95311, -10.78669, -10.61998, 
    -10.45297, -10.28566, -10.11806, -9.950154, -9.781957, -9.613465, 
    -9.44468, -9.2756, -9.106229, -8.936565, -8.766611, -8.596366, -8.425832, 
    -8.255008, -8.083897, -7.912498, -7.740814, -7.568844, -7.39659, 
    -7.224052, -7.051232, -6.878131, -6.704749, -6.531086, -6.357146, 
    -6.182928, -6.008433, -5.833663, -5.658619, -5.483302, -5.307712, 
    -5.131851, -4.955721, -4.779322, -4.602656, -4.425724, -4.248526, 
    -4.071065, -3.893342, -3.715357, -3.537113, -3.358611, -3.179851, 
    -3.000836, -2.821566, -2.642044, -2.46227, -2.282247, -2.101974, 
    -1.921456, -1.740691, -1.559682, -1.378432, -1.19694, -1.015209, 
    -0.833241, -0.6510367, -0.4685981, -0.2859269, -0.1030247, 0.08010672, 
    0.2634656, 0.4470503, 0.630859, 0.8148899, 0.9991412, 1.183611, 1.368298, 
    1.553199, 1.738314, 1.92364, 2.109175, 2.294917, 2.480865, 2.667016, 
    2.853368, 3.03992, 3.226669, 3.413613, 3.600751, 3.78808, 3.975598, 
    4.163303, 4.351193, 4.539266, 4.727519, 4.915951, 5.104558, 5.293341, 
    5.482294, 5.671418, 5.860708, 6.050164, 6.239782, 6.429562, 6.619499, 
    6.809591, 6.999838, 7.190236, 7.380782, 7.571474, 7.762311, 7.953289, 
    8.144406, 8.33566, 8.527048, 8.718568, 8.910217, 9.101993, 9.293893, 
    9.485915, 9.678056, 9.870314, 10.06269, 10.25517, 10.44776, 10.64046, 
    10.83326, 11.02617, 11.21917, 11.41227, 11.60546, 11.79874, 11.99211, 
    12.18557, 12.3791, 12.57272, 12.76642, 12.96019, 13.15403, 13.34794, 
    13.54192, 13.73596, 13.93006, 14.12422, 14.31844, 14.51271, 14.70703, 
    14.90139, 15.0958, 15.29025, 15.48475, 15.67927, 15.87383, 16.06842, 
    16.26304, 16.45769, 16.65235, 16.84704, 17.04174, 17.23646, 17.43118, 
    17.62592, 17.82066, 18.0154, 18.21015, 18.40488, 18.59962, 18.79434, 
    18.98906, 19.18376, 19.37844, 19.5731, 19.76774, 19.96236, 20.15694, 
    20.3515, 20.54602, 20.74051, 20.93495, 21.12936, 21.32372, 21.51803, 
    21.71229, 21.90649, 22.10065, 22.29474, 22.48877, 22.68274, 22.87664, 
    23.07047, 23.26423, 23.45791, 23.65152, 23.84504, 24.03848, 24.23184, 
    24.42511, 24.61828, 24.81137, 25.00435, 25.19724, 25.39003, 25.58271, 
    25.77529, 25.96775, 26.16011, 26.35234, 26.54447, 26.73647, 26.92835, 
    27.12011, 27.31174, 27.50323, 27.6946, 27.88583, 28.07693, 28.26789, 
    28.4587, 28.64937, 28.83989, 29.03027, 29.22049, 29.41056, 29.60047, 
    29.79022, 29.97982, 30.16924, 30.35851, 30.54761, 30.73653, 30.92529, 
    31.11387, 31.30227, 31.4905, 31.67854, 31.8664, 32.05408, 32.24157, 
    32.42886, 32.61597, 32.80289, 32.9896, 33.17612, 33.36245, 33.54856, 
    33.73448, 33.92019, 34.10569, 34.29098, 34.47606, 34.66093, 34.84558, 
    35.03002, 35.21424, 35.39823, 35.582, 35.76555, 35.94888, 36.13197, 
    36.31484, 36.49747, 36.67987, 36.86204, 37.04397, 37.22567, 37.40712, 
    37.58833, 37.7693, 37.95003, 38.13051, 38.31074, 38.49072, 38.67046, 
    38.84994, 39.02917, 39.20815, 39.38686, 39.56533, 39.74353, 39.92147, 
    40.09916, 40.27657, 40.45373, 40.63062, 40.80724, 40.9836, 41.15969, 
    41.33551, 41.51105, 41.68633, 41.86133, 42.03605, 42.21051, 42.38468, 
    42.55857, 42.73219, 42.90553, 43.07859, 43.25137, 43.42386, 43.59607, 
    43.76799, 43.93963, 44.11098, 44.28205, 44.45283, 44.62331, 44.79351, 
    44.96342, 45.13304, 45.30236, 45.4714, 45.64014, 45.80858, 45.97673, 
    46.14459, 46.31215, 46.47941, 46.64637, 46.81304, 46.97941, 47.14547, 
    47.31124, 47.47671, 47.64188, 47.80675, 47.97131, 48.13557, 48.29953, 
    48.46319, 48.62654, 48.7896, 48.95234, 49.11478, 49.27692,
  -27.08492, -26.95078, -26.81635, -26.68163, -26.54663, -26.41134, 
    -26.27575, -26.13988, -26.00371, -25.86726, -25.73051, -25.59347, 
    -25.45613, -25.3185, -25.18058, -25.04236, -24.90385, -24.76504, 
    -24.62593, -24.48653, -24.34683, -24.20683, -24.06654, -23.92595, 
    -23.78505, -23.64386, -23.50236, -23.36057, -23.21847, -23.07608, 
    -22.93338, -22.79038, -22.64707, -22.50347, -22.35956, -22.21534, 
    -22.07083, -21.926, -21.78087, -21.63544, -21.4897, -21.34366, -21.19731, 
    -21.05065, -20.90368, -20.75641, -20.60884, -20.46095, -20.31275, 
    -20.16425, -20.01544, -19.86632, -19.71689, -19.56715, -19.4171, 
    -19.26675, -19.11608, -18.9651, -18.81382, -18.66222, -18.51031, 
    -18.3581, -18.20557, -18.05273, -17.89958, -17.74612, -17.59235, 
    -17.43826, -17.28387, -17.12917, -16.97415, -16.81883, -16.66319, 
    -16.50724, -16.35098, -16.19441, -16.03753, -15.88034, -15.72284, 
    -15.56503, -15.4069, -15.24847, -15.08973, -14.93067, -14.77131, 
    -14.61164, -14.45166, -14.29136, -14.13076, -13.96985, -13.80864, 
    -13.64711, -13.48528, -13.32313, -13.16068, -12.99793, -12.83487, 
    -12.6715, -12.50782, -12.34384, -12.17956, -12.01497, -11.85007, 
    -11.68488, -11.51937, -11.35357, -11.18746, -11.02106, -10.85435, 
    -10.68734, -10.52003, -10.35242, -10.18451, -10.01631, -9.847806, 
    -9.679007, -9.509911, -9.340519, -9.170834, -9.000854, -8.83058, 
    -8.660014, -8.489157, -8.318009, -8.146571, -7.974844, -7.802828, 
    -7.630526, -7.457936, -7.285061, -7.111902, -6.938459, -6.764733, 
    -6.590725, -6.416437, -6.241869, -6.067023, -5.8919, -5.716499, 
    -5.540824, -5.364874, -5.188652, -5.012157, -4.835392, -4.658358, 
    -4.481055, -4.303485, -4.12565, -3.94755, -3.769187, -3.590563, 
    -3.411678, -3.232534, -3.053133, -2.873475, -2.693562, -2.513396, 
    -2.332978, -2.15231, -1.971393, -1.790228, -1.608818, -1.427163, 
    -1.245266, -1.063127, -0.880749, -0.6981331, -0.515281, -0.3321944, 
    -0.1488751, 0.03467543, 0.2184553, 0.4024627, 0.586696, 0.7711533, 
    0.9558328, 1.140733, 1.325851, 1.511186, 1.696736, 1.882499, 2.068473, 
    2.254655, 2.441045, 2.62764, 2.814438, 3.001437, 3.188635, 3.376029, 
    3.563619, 3.751402, 3.939375, 4.127537, 4.315886, 4.504418, 4.693133, 
    4.882028, 5.0711, 5.260348, 5.449769, 5.639362, 5.829123, 6.019051, 
    6.209142, 6.399395, 6.589808, 6.780379, 6.971104, 7.161981, 7.353008, 
    7.544183, 7.735503, 7.926966, 8.118569, 8.31031, 8.502188, 8.694197, 
    8.886336, 9.078604, 9.270997, 9.463513, 9.656149, 9.848903, 10.04177, 
    10.23475, 10.42784, 10.62104, 10.81435, 11.00775, 11.20126, 11.39486, 
    11.58855, 11.78234, 11.97622, 12.17018, 12.36422, 12.55835, 12.75255, 
    12.94683, 13.14119, 13.33561, 13.5301, 13.72465, 13.91926, 14.11394, 
    14.30867, 14.50345, 14.69828, 14.89316, 15.08809, 15.28306, 15.47806, 
    15.67311, 15.86818, 16.06329, 16.25843, 16.45359, 16.64877, 16.84397, 
    17.03919, 17.23443, 17.42967, 17.62492, 17.82018, 18.01544, 18.2107, 
    18.40596, 18.60121, 18.79646, 18.99169, 19.18691, 19.38211, 19.57729, 
    19.77244, 19.96758, 20.16268, 20.35775, 20.55279, 20.74779, 20.94275, 
    21.13767, 21.33254, 21.52737, 21.72214, 21.91686, 22.11152, 22.30613, 
    22.50067, 22.69515, 22.88956, 23.0839, 23.27817, 23.47236, 23.66648, 
    23.86051, 24.05446, 24.24832, 24.44209, 24.63577, 24.82936, 25.02285, 
    25.21624, 25.40952, 25.60271, 25.79578, 25.98874, 26.18159, 26.37433, 
    26.56695, 26.75945, 26.95182, 27.14407, 27.33619, 27.52817, 27.72003, 
    27.91175, 28.10333, 28.29477, 28.48607, 28.67722, 28.86822, 29.05908, 
    29.24978, 29.44032, 29.63071, 29.82094, 30.011, 30.2009, 30.39064, 
    30.58021, 30.7696, 30.95882, 31.14786, 31.33673, 31.52542, 31.71392, 
    31.90224, 32.09037, 32.27832, 32.46607, 32.65363, 32.84099, 33.02816, 
    33.21512, 33.40189, 33.58845, 33.77481, 33.96096, 34.1469, 34.33263, 
    34.51815, 34.70345, 34.88853, 35.07339, 35.25804, 35.44246, 35.62666, 
    35.81063, 35.99437, 36.17789, 36.36117, 36.54422, 36.72704, 36.90961, 
    37.09195, 37.27406, 37.45591, 37.63753, 37.8189, 38.00003, 38.1809, 
    38.36153, 38.54191, 38.72204, 38.90191, 39.08153, 39.26089, 39.43999, 
    39.61884, 39.79742, 39.97574, 40.1538, 40.33159, 40.50912, 40.68638, 
    40.86337, 41.04009, 41.21655, 41.39272, 41.56863, 41.74426, 41.91962, 
    42.0947, 42.2695, 42.44403, 42.61827, 42.79223, 42.96591, 43.13931, 
    43.31243, 43.48526, 43.6578, 43.83006, 44.00203, 44.17371, 44.3451, 
    44.5162, 44.68702, 44.85753, 45.02776, 45.19769, 45.36733, 45.53668, 
    45.70573, 45.87448, 46.04294, 46.21109, 46.37896, 46.54652, 46.71378, 
    46.88074, 47.0474, 47.21376, 47.37982, 47.54557, 47.71103, 47.87618, 
    48.04102, 48.20557, 48.3698, 48.53373, 48.69736, 48.86068, 49.02369, 
    49.1864, 49.3488,
  -27.1738, -27.03956, -26.90502, -26.7702, -26.63508, -26.49967, -26.36397, 
    -26.22799, -26.0917, -25.95513, -25.81826, -25.6811, -25.54364, 
    -25.40589, -25.26784, -25.1295, -24.99085, -24.85192, -24.71268, 
    -24.57314, -24.43331, -24.29318, -24.15275, -24.01201, -23.87098, 
    -23.72965, -23.58801, -23.44607, -23.30383, -23.16129, -23.01844, 
    -22.87529, -22.73183, -22.58807, -22.44401, -22.29963, -22.15496, 
    -22.00997, -21.86469, -21.71909, -21.57318, -21.42697, -21.28045, 
    -21.13363, -20.98649, -20.83904, -20.69129, -20.54323, -20.39485, 
    -20.24617, -20.09718, -19.94787, -19.79826, -19.64833, -19.4981, 
    -19.34755, -19.19669, -19.04552, -18.89404, -18.74224, -18.59013, 
    -18.43772, -18.28498, -18.13194, -17.97858, -17.82491, -17.67093, 
    -17.51664, -17.36203, -17.20711, -17.05188, -16.89633, -16.74047, 
    -16.5843, -16.42781, -16.27102, -16.11391, -15.95648, -15.79875, 
    -15.6407, -15.48234, -15.32367, -15.16468, -15.00538, -14.84577, 
    -14.68585, -14.52562, -14.36508, -14.20423, -14.04306, -13.88159, 
    -13.7198, -13.5577, -13.3953, -13.23258, -13.06956, -12.90623, -12.74259, 
    -12.57864, -12.41438, -12.24982, -12.08495, -11.91978, -11.7543, 
    -11.58851, -11.42242, -11.25602, -11.08932, -10.92232, -10.75501, 
    -10.58741, -10.4195, -10.25129, -10.08278, -9.913966, -9.744857, 
    -9.57545, -9.405746, -9.235744, -9.065448, -8.894855, -8.723968, 
    -8.552787, -8.381313, -8.209547, -8.037491, -7.865143, -7.692506, 
    -7.519581, -7.346367, -7.172868, -6.999082, -6.825012, -6.650658, 
    -6.476021, -6.301102, -6.125903, -5.950424, -5.774667, -5.598632, 
    -5.422321, -5.245735, -5.068876, -4.891743, -4.714339, -4.536665, 
    -4.358722, -4.180511, -4.002033, -3.823291, -3.644285, -3.465016, 
    -3.285486, -3.105697, -2.925649, -2.745345, -2.564785, -2.383971, 
    -2.202905, -2.021588, -1.840022, -1.658208, -1.476148, -1.293843, 
    -1.111294, -0.9285049, -0.7454757, -0.5622084, -0.3787047, -0.1949663, 
    -0.0109949, 0.1732077, 0.3576398, 0.5422994, 0.7271851, 0.9122947, 
    1.097626, 1.283179, 1.468949, 1.654936, 1.841138, 2.027553, 2.214178, 
    2.401012, 2.588053, 2.775298, 2.962747, 3.150395, 3.338243, 3.526287, 
    3.714526, 3.902956, 4.091578, 4.280387, 4.469382, 4.65856, 4.84792, 
    5.03746, 5.227176, 5.417067, 5.607131, 5.797364, 5.987766, 6.178333, 
    6.369063, 6.559955, 6.751005, 6.942211, 7.13357, 7.325081, 7.516741, 
    7.708548, 7.900498, 8.092589, 8.284821, 8.477188, 8.66969, 8.862323, 
    9.055085, 9.247973, 9.440986, 9.63412, 9.827372, 10.02074, 10.21422, 
    10.40782, 10.60152, 10.79532, 10.98923, 11.18324, 11.37735, 11.57155, 
    11.76585, 11.96023, 12.15471, 12.34926, 12.5439, 12.73861, 12.9334, 
    13.12827, 13.3232, 13.51821, 13.71327, 13.9084, 14.10359, 14.29884, 
    14.49414, 14.68949, 14.88489, 15.08033, 15.27582, 15.47134, 15.6669, 
    15.8625, 16.05813, 16.25378, 16.44946, 16.64517, 16.84089, 17.03663, 
    17.23238, 17.42815, 17.62392, 17.8197, 18.01548, 18.21127, 18.40705, 
    18.60282, 18.79858, 18.99433, 19.19007, 19.38579, 19.58149, 19.77717, 
    19.97282, 20.16844, 20.36403, 20.55959, 20.75511, 20.95059, 21.14603, 
    21.34142, 21.53676, 21.73205, 21.92729, 22.12247, 22.31759, 22.51264, 
    22.70764, 22.90256, 23.09741, 23.29219, 23.4869, 23.68152, 23.87606, 
    24.07052, 24.26489, 24.45917, 24.65336, 24.84745, 25.04145, 25.23534, 
    25.42913, 25.62281, 25.81639, 26.00986, 26.20321, 26.39644, 26.58955, 
    26.78255, 26.97542, 27.16816, 27.36077, 27.55325, 27.7456, 27.93781, 
    28.12988, 28.3218, 28.51359, 28.70522, 28.89671, 29.08805, 29.27923, 
    29.47025, 29.66112, 29.85182, 30.04236, 30.23274, 30.42295, 30.61298, 
    30.80285, 30.99253, 31.18204, 31.37138, 31.56053, 31.74949, 31.93827, 
    32.12686, 32.31526, 32.50347, 32.69149, 32.8793, 33.06692, 33.25433, 
    33.44155, 33.62856, 33.81536, 34.00195, 34.18833, 34.3745, 34.56045, 
    34.74619, 34.93171, 35.117, 35.30207, 35.48693, 35.67155, 35.85595, 
    36.04011, 36.22404, 36.40775, 36.59121, 36.77444, 36.95744, 37.14019, 
    37.3227, 37.50496, 37.68699, 37.86876, 38.05029, 38.23156, 38.41259, 
    38.59336, 38.77388, 38.95415, 39.13416, 39.3139, 39.49339, 39.67262, 
    39.85158, 40.03028, 40.20872, 40.38689, 40.56479, 40.74242, 40.91978, 
    41.09687, 41.27369, 41.45023, 41.6265, 41.80249, 41.9782, 42.15364, 
    42.32879, 42.50367, 42.67826, 42.85257, 43.02659, 43.20033, 43.37379, 
    43.54696, 43.71983, 43.89243, 44.06473, 44.23674, 44.40846, 44.57988, 
    44.75102, 44.92186, 45.09241, 45.26266, 45.43261, 45.60227, 45.77163, 
    45.94069, 46.10945, 46.27791, 46.44608, 46.61394, 46.7815, 46.94876, 
    47.11571, 47.28236, 47.44871, 47.61475, 47.78049, 47.94593, 48.11105, 
    48.27588, 48.44039, 48.6046, 48.76849, 48.93209, 49.09537, 49.25834, 
    49.42101,
  -27.26299, -27.12864, -26.994, -26.85906, -26.72383, -26.58832, -26.45251, 
    -26.3164, -26.18, -26.04331, -25.90632, -25.76904, -25.63146, -25.49359, 
    -25.35542, -25.21694, -25.07818, -24.93911, -24.79974, -24.66008, 
    -24.52011, -24.37984, -24.23927, -24.0984, -23.95723, -23.81575, 
    -23.67397, -23.53189, -23.38951, -23.24681, -23.10382, -22.96052, 
    -22.81691, -22.673, -22.52878, -22.38425, -22.23941, -22.09427, 
    -21.94882, -21.80306, -21.65699, -21.51061, -21.36393, -21.21693, 
    -21.06962, -20.922, -20.77407, -20.62583, -20.47728, -20.32842, 
    -20.17924, -20.02976, -19.87996, -19.72984, -19.57942, -19.42868, 
    -19.27763, -19.12626, -18.97458, -18.82259, -18.67028, -18.51766, 
    -18.36473, -18.21148, -18.05792, -17.90404, -17.74985, -17.59534, 
    -17.44052, -17.28538, -17.12993, -16.97416, -16.81808, -16.66168, 
    -16.50497, -16.34795, -16.19061, -16.03295, -15.87498, -15.7167, 
    -15.5581, -15.39919, -15.23996, -15.08042, -14.92057, -14.7604, 
    -14.59992, -14.43912, -14.27802, -14.11659, -13.95486, -13.79282, 
    -13.63046, -13.46779, -13.30481, -13.14152, -12.97792, -12.814, 
    -12.64978, -12.48525, -12.32041, -12.15526, -11.9898, -11.82403, 
    -11.65796, -11.49158, -11.32489, -11.1579, -10.9906, -10.823, -10.6551, 
    -10.48689, -10.31837, -10.14956, -9.980438, -9.81102, -9.641302, 
    -9.471284, -9.300966, -9.130351, -8.959438, -8.788229, -8.616724, 
    -8.444923, -8.272829, -8.100441, -7.927761, -7.754788, -7.581526, 
    -7.407973, -7.234132, -7.060003, -6.885587, -6.710885, -6.535899, 
    -6.360628, -6.185075, -6.00924, -5.833124, -5.656729, -5.480056, 
    -5.303105, -5.125879, -4.948378, -4.770603, -4.592556, -4.414238, 
    -4.23565, -4.056794, -3.87767, -3.69828, -3.518626, -3.33871, -3.158531, 
    -2.978092, -2.797394, -2.616439, -2.435228, -2.253762, -2.072044, 
    -1.890074, -1.707855, -1.525387, -1.342673, -1.159714, -0.9765111, 
    -0.7930667, -0.6093825, -0.4254598, -0.2413005, -0.05690642, 0.1277208, 
    0.3125793, 0.4976674, 0.6829832, 0.8685248, 1.054291, 1.240278, 1.426486, 
    1.612913, 1.799556, 1.986413, 2.173483, 2.360763, 2.548252, 2.735947, 
    2.923847, 3.111949, 3.300252, 3.488752, 3.677449, 3.86634, 4.055422, 
    4.244694, 4.434154, 4.623798, 4.813626, 5.003634, 5.193821, 5.384185, 
    5.574722, 5.765431, 5.956309, 6.147354, 6.338564, 6.529936, 6.721468, 
    6.913157, 7.105002, 7.296999, 7.489146, 7.681442, 7.873882, 8.066465, 
    8.259189, 8.452049, 8.645046, 8.838175, 9.031434, 9.224821, 9.418332, 
    9.611966, 9.80572, 9.999591, 10.19358, 10.38767, 10.58188, 10.77619, 
    10.97061, 11.16513, 11.35975, 11.55446, 11.74926, 11.94416, 12.13914, 
    12.33421, 12.52936, 12.72459, 12.9199, 13.11528, 13.31073, 13.50625, 
    13.70184, 13.89748, 14.09319, 14.28895, 14.48477, 14.68064, 14.87656, 
    15.07253, 15.26853, 15.46458, 15.66066, 15.85678, 16.05293, 16.24911, 
    16.44531, 16.64154, 16.83779, 17.03405, 17.23033, 17.42662, 17.62292, 
    17.81922, 18.01553, 18.21183, 18.40813, 18.60443, 18.80072, 18.99699, 
    19.19326, 19.3895, 19.58572, 19.78192, 19.9781, 20.17424, 20.37036, 
    20.56643, 20.76247, 20.95848, 21.15443, 21.35034, 21.54621, 21.74202, 
    21.93777, 22.13347, 22.32911, 22.52468, 22.72019, 22.91563, 23.111, 
    23.3063, 23.50151, 23.69665, 23.8917, 24.08668, 24.28156, 24.47635, 
    24.67105, 24.86565, 25.06015, 25.25455, 25.44885, 25.64304, 25.83712, 
    26.03108, 26.22494, 26.41867, 26.61229, 26.80578, 26.99915, 27.19238, 
    27.38549, 27.57847, 27.77131, 27.96401, 28.15657, 28.34899, 28.54126, 
    28.73338, 28.92535, 29.11717, 29.30884, 29.50035, 29.69169, 29.88288, 
    30.0739, 30.26475, 30.45543, 30.64594, 30.83628, 31.02643, 31.21641, 
    31.40621, 31.59583, 31.78526, 31.9745, 32.16355, 32.35241, 32.54108, 
    32.72955, 32.91782, 33.10589, 33.29376, 33.48142, 33.66888, 33.85612, 
    34.04316, 34.22998, 34.41659, 34.60298, 34.78916, 34.97511, 35.16084, 
    35.34634, 35.53162, 35.71668, 35.9015, 36.08609, 36.27045, 36.45457, 
    36.63845, 36.8221, 37.00551, 37.18867, 37.37159, 37.55427, 37.73669, 
    37.91888, 38.10081, 38.28249, 38.46391, 38.64508, 38.826, 39.00665, 
    39.18705, 39.36719, 39.54706, 39.72667, 39.90602, 40.0851, 40.26392, 
    40.44246, 40.62074, 40.79874, 40.97647, 41.15393, 41.33112, 41.50802, 
    41.68465, 41.861, 42.03707, 42.21286, 42.38837, 42.5636, 42.73854, 
    42.9132, 43.08757, 43.26165, 43.43545, 43.60895, 43.78217, 43.95509, 
    44.12773, 44.30007, 44.47212, 44.64387, 44.81533, 44.98649, 45.15736, 
    45.32793, 45.4982, 45.66817, 45.83784, 46.00721, 46.17628, 46.34505, 
    46.51351, 46.68167, 46.84953, 47.01709, 47.18434, 47.35128, 47.51792, 
    47.68425, 47.85028, 48.016, 48.1814, 48.3465, 48.5113, 48.67578, 
    48.83995, 49.00381, 49.16737, 49.33061, 49.49354,
  -27.35249, -27.21803, -27.08328, -26.94824, -26.8129, -26.67727, -26.54135, 
    -26.40513, -26.26862, -26.13181, -25.9947, -25.8573, -25.7196, -25.5816, 
    -25.44331, -25.30471, -25.16581, -25.02662, -24.88712, -24.74732, 
    -24.60723, -24.46682, -24.32612, -24.18511, -24.0438, -23.90218, 
    -23.76026, -23.61804, -23.47551, -23.33267, -23.18952, -23.04607, 
    -22.90231, -22.75825, -22.61387, -22.46919, -22.3242, -22.17889, 
    -22.03328, -21.88736, -21.74113, -21.59458, -21.44773, -21.30056, 
    -21.15308, -21.00529, -20.85719, -20.70877, -20.56004, -20.411, 
    -20.26164, -20.11197, -19.96198, -19.81169, -19.66107, -19.51014, 
    -19.3589, -19.20734, -19.05546, -18.90327, -18.75077, -18.59794, 
    -18.44481, -18.29135, -18.13758, -17.9835, -17.82909, -17.67437, 
    -17.51933, -17.36398, -17.20831, -17.05232, -16.89602, -16.7394, 
    -16.58246, -16.42521, -16.26764, -16.10975, -15.95155, -15.79303, 
    -15.63419, -15.47504, -15.31557, -15.15579, -14.99569, -14.83527, 
    -14.67454, -14.51349, -14.35213, -14.19046, -14.02847, -13.86616, 
    -13.70354, -13.54061, -13.37736, -13.2138, -13.04993, -12.88575, 
    -12.72125, -12.55644, -12.39132, -12.22589, -12.06015, -11.8941, 
    -11.72774, -11.56107, -11.39409, -11.2268, -11.05921, -10.89131, 
    -10.7231, -10.55459, -10.38577, -10.21665, -10.04723, -9.877499, 
    -9.707467, -9.537134, -9.3665, -9.195566, -9.024332, -8.852799, 
    -8.680969, -8.508842, -8.336417, -8.163697, -7.990684, -7.817376, 
    -7.643775, -7.469882, -7.295698, -7.121224, -6.946462, -6.771411, 
    -6.596074, -6.42045, -6.244542, -6.068349, -5.891874, -5.715117, 
    -5.538081, -5.360765, -5.18317, -5.005299, -4.827152, -4.648731, 
    -4.470036, -4.29107, -4.111833, -3.932327, -3.752553, -3.572512, 
    -3.392206, -3.211637, -3.030805, -2.849712, -2.66836, -2.48675, 
    -2.304884, -2.122762, -1.940388, -1.757761, -1.574885, -1.391759, 
    -1.208387, -1.02477, -0.8409085, -0.6568053, -0.4724619, -0.28788, 
    -0.1030613, 0.08199235, 0.2672793, 0.4527976, 0.6385455, 0.8245212, 
    1.010723, 1.197148, 1.383796, 1.570664, 1.75775, 1.945052, 2.132568, 
    2.320297, 2.508236, 2.696383, 2.884737, 3.073294, 3.262053, 3.451013, 
    3.64017, 3.829523, 4.019069, 4.208806, 4.398732, 4.588845, 4.779143, 
    4.969623, 5.160283, 5.351121, 5.542134, 5.733321, 5.924678, 6.116203, 
    6.307895, 6.499751, 6.691767, 6.883943, 7.076274, 7.268761, 7.461398, 
    7.654184, 7.847117, 8.040195, 8.233413, 8.42677, 8.620264, 8.813891, 
    9.00765, 9.201538, 9.395552, 9.589688, 9.783946, 9.978323, 10.17281, 
    10.36742, 10.56213, 10.75696, 10.95188, 11.14691, 11.34204, 11.53727, 
    11.73258, 11.92799, 12.12349, 12.31908, 12.51474, 12.71049, 12.90632, 
    13.10221, 13.29819, 13.49423, 13.69033, 13.8865, 14.08273, 14.27901, 
    14.47536, 14.67175, 14.86819, 15.06468, 15.26121, 15.45778, 15.65439, 
    15.85103, 16.04771, 16.24441, 16.44114, 16.6379, 16.83467, 17.03146, 
    17.22826, 17.42508, 17.6219, 17.81874, 18.01557, 18.2124, 18.40923, 
    18.60605, 18.80287, 18.99967, 19.19646, 19.39323, 19.58998, 19.7867, 
    19.9834, 20.18007, 20.37671, 20.57331, 20.76988, 20.96641, 21.16289, 
    21.35932, 21.55571, 21.75204, 21.94832, 22.14454, 22.34069, 22.53679, 
    22.73282, 22.92878, 23.12466, 23.32048, 23.51621, 23.71187, 23.90744, 
    24.10292, 24.29832, 24.49362, 24.68883, 24.88395, 25.07896, 25.27387, 
    25.46867, 25.66337, 25.85796, 26.05243, 26.24679, 26.44103, 26.63515, 
    26.82914, 27.02301, 27.21675, 27.41035, 27.60382, 27.79716, 27.99036, 
    28.18341, 28.37632, 28.56908, 28.7617, 28.95416, 29.14647, 29.33862, 
    29.53061, 29.72244, 29.9141, 30.1056, 30.29693, 30.48809, 30.67908, 
    30.86989, 31.06052, 31.25097, 31.44124, 31.63132, 31.82122, 32.01093, 
    32.20044, 32.38976, 32.57889, 32.76782, 32.95655, 33.14507, 33.33339, 
    33.52151, 33.70941, 33.89711, 34.08459, 34.27186, 34.45891, 34.64574, 
    34.83236, 35.01875, 35.20491, 35.39085, 35.57656, 35.76205, 35.9473, 
    36.13231, 36.31709, 36.50164, 36.68594, 36.87001, 37.05383, 37.23741, 
    37.42074, 37.60383, 37.78667, 37.96925, 38.15159, 38.33367, 38.5155, 
    38.69706, 38.87838, 39.05943, 39.24022, 39.42075, 39.60101, 39.78101, 
    39.96074, 40.1402, 40.3194, 40.49832, 40.67697, 40.85535, 41.03345, 
    41.21128, 41.38883, 41.5661, 41.7431, 41.91981, 42.09624, 42.27238, 
    42.44825, 42.62383, 42.79912, 42.97412, 43.14884, 43.32327, 43.49741, 
    43.67125, 43.84481, 44.01807, 44.19104, 44.36371, 44.53609, 44.70817, 
    44.87995, 45.05144, 45.22263, 45.39351, 45.5641, 45.73438, 45.90437, 
    46.07405, 46.24342, 46.4125, 46.58127, 46.74973, 46.91789, 47.08574, 
    47.25328, 47.42052, 47.58745, 47.75407, 47.92038, 48.08639, 48.25208, 
    48.41746, 48.58253, 48.74729, 48.91174, 49.07587, 49.2397, 49.40321, 
    49.5664,
  -27.4423, -27.30774, -27.17288, -27.03773, -26.90228, -26.76654, -26.6305, 
    -26.49417, -26.35754, -26.22062, -26.0834, -25.94587, -25.80805, 
    -25.66993, -25.53151, -25.39279, -25.25377, -25.11445, -24.97482, 
    -24.83489, -24.69466, -24.55413, -24.41329, -24.27214, -24.13069, 
    -23.98894, -23.84687, -23.70451, -23.56183, -23.41885, -23.27555, 
    -23.13195, -22.98804, -22.84382, -22.6993, -22.55445, -22.40931, 
    -22.26384, -22.11807, -21.97199, -21.82559, -21.67888, -21.53186, 
    -21.38452, -21.23687, -21.08891, -20.94063, -20.79204, -20.64313, 
    -20.49391, -20.34437, -20.19451, -20.04434, -19.89386, -19.74306, 
    -19.59194, -19.4405, -19.28875, -19.13668, -18.98429, -18.83158, 
    -18.67856, -18.52522, -18.37156, -18.21758, -18.06329, -17.90867, 
    -17.75374, -17.59849, -17.44292, -17.28703, -17.13082, -16.9743, 
    -16.81745, -16.66029, -16.50281, -16.34501, -16.18689, -16.02845, 
    -15.86969, -15.71062, -15.55123, -15.39152, -15.23149, -15.07114, 
    -14.91048, -14.7495, -14.5882, -14.42658, -14.26465, -14.1024, -13.93983, 
    -13.77695, -13.61376, -13.45024, -13.28641, -13.12227, -12.95781, 
    -12.79304, -12.62796, -12.46256, -12.29685, -12.13082, -11.96448, 
    -11.79784, -11.63088, -11.46361, -11.29603, -11.12814, -10.95994, 
    -10.79143, -10.62262, -10.4535, -10.28407, -10.11433, -9.944294, 
    -9.77395, -9.603301, -9.432349, -9.261095, -9.08954, -8.917684, 
    -8.745526, -8.573071, -8.400315, -8.227263, -8.053914, -7.88027, 
    -7.706329, -7.532095, -7.357568, -7.182749, -7.007638, -6.832238, 
    -6.656548, -6.48057, -6.304306, -6.127755, -5.950919, -5.773799, 
    -5.596398, -5.418715, -5.240751, -5.062508, -4.883988, -4.705191, 
    -4.526119, -4.346773, -4.167154, -3.987264, -3.807104, -3.626675, 
    -3.445979, -3.265017, -3.083791, -2.902302, -2.720551, -2.538541, 
    -2.356272, -2.173746, -1.990965, -1.807929, -1.624642, -1.441104, 
    -1.257317, -1.073283, -0.8890032, -0.7044794, -0.5197135, -0.334707, 
    -0.1494619, 0.03602016, 0.2217374, 0.4076879, 0.5938699, 0.7802815, 
    0.9669209, 1.153786, 1.340875, 1.528186, 1.715717, 1.903467, 2.091432, 
    2.279611, 2.468003, 2.656604, 2.845413, 3.034428, 3.223647, 3.413067, 
    3.602687, 3.792504, 3.982516, 4.17272, 4.363116, 4.5537, 4.74447, 
    4.935424, 5.126559, 5.317874, 5.509366, 5.701032, 5.892871, 6.084879, 
    6.277056, 6.469397, 6.661901, 6.854565, 7.047387, 7.240364, 7.433494, 
    7.626774, 7.820202, 8.013776, 8.207492, 8.401348, 8.595342, 8.789471, 
    8.983732, 9.178123, 9.372642, 9.567285, 9.76205, 9.956934, 10.15193, 
    10.34705, 10.54227, 10.73761, 10.93305, 11.12859, 11.32423, 11.51997, 
    11.71581, 11.91174, 12.10775, 12.30386, 12.50004, 12.69631, 12.89266, 
    13.08908, 13.28557, 13.48213, 13.67876, 13.87545, 14.07221, 14.26902, 
    14.46588, 14.6628, 14.85977, 15.05679, 15.25385, 15.45094, 15.64808, 
    15.84525, 16.04246, 16.23969, 16.43695, 16.63423, 16.83153, 17.02885, 
    17.22619, 17.42353, 17.62089, 17.81825, 18.01561, 18.21297, 18.41033, 
    18.60769, 18.80503, 19.00236, 19.19968, 19.39698, 19.59426, 19.79151, 
    19.98874, 20.18594, 20.3831, 20.58024, 20.77733, 20.97438, 21.17139, 
    21.36835, 21.56526, 21.76212, 21.95892, 22.15566, 22.35235, 22.54897, 
    22.74552, 22.942, 23.13841, 23.33474, 23.531, 23.72717, 23.92326, 
    24.11926, 24.31517, 24.51099, 24.70672, 24.90235, 25.09787, 25.2933, 
    25.48862, 25.68382, 25.87892, 26.0739, 26.26877, 26.46351, 26.65814, 
    26.85263, 27.047, 27.24125, 27.43535, 27.62933, 27.82316, 28.01685, 
    28.21041, 28.40381, 28.59707, 28.79017, 28.98313, 29.17592, 29.36856, 
    29.56104, 29.75336, 29.94551, 30.13749, 30.3293, 30.52094, 30.7124, 
    30.90369, 31.09479, 31.28572, 31.47646, 31.66702, 31.85738, 32.04755, 
    32.23753, 32.42732, 32.61691, 32.8063, 32.99548, 33.18447, 33.37325, 
    33.56181, 33.75017, 33.93832, 34.12625, 34.31396, 34.50146, 34.68874, 
    34.87579, 35.06262, 35.24922, 35.4356, 35.62174, 35.80766, 35.99334, 
    36.17878, 36.36399, 36.54896, 36.73368, 36.91817, 37.10241, 37.28641, 
    37.47015, 37.65365, 37.8369, 38.01989, 38.20264, 38.38512, 38.56735, 
    38.74932, 38.93103, 39.11248, 39.29366, 39.47458, 39.65524, 39.83562, 
    40.01574, 40.19558, 40.37516, 40.55446, 40.73349, 40.91225, 41.09072, 
    41.26892, 41.44684, 41.62448, 41.80183, 41.97891, 42.1557, 42.33221, 
    42.50843, 42.68436, 42.86, 43.03536, 43.21042, 43.3852, 43.55968, 
    43.73386, 43.90776, 44.08136, 44.25466, 44.42766, 44.60037, 44.77278, 
    44.94489, 45.1167, 45.2882, 45.45941, 45.63031, 45.80091, 45.97121, 
    46.1412, 46.31089, 46.48027, 46.64934, 46.81811, 46.98657, 47.15472, 
    47.32256, 47.49009, 47.65731, 47.82422, 47.99082, 48.1571, 48.32308, 
    48.48874, 48.65409, 48.81913, 48.98385, 49.14826, 49.31235, 49.47613, 
    49.63959,
  -27.53242, -27.39775, -27.26279, -27.12753, -26.99197, -26.85612, 
    -26.71998, -26.58353, -26.44679, -26.30975, -26.17241, -26.03477, 
    -25.89683, -25.75858, -25.62004, -25.4812, -25.34205, -25.2026, 
    -25.06285, -24.92279, -24.78242, -24.64175, -24.50078, -24.3595, 
    -24.21791, -24.07602, -23.93381, -23.7913, -23.64848, -23.50535, 
    -23.36191, -23.21816, -23.0741, -22.92973, -22.78505, -22.64005, 
    -22.49475, -22.34912, -22.20319, -22.05694, -21.91038, -21.76351, 
    -21.61632, -21.46881, -21.32099, -21.17286, -21.0244, -20.87564, 
    -20.72655, -20.57715, -20.42743, -20.27739, -20.12704, -19.97637, 
    -19.82537, -19.67407, -19.52244, -19.37049, -19.21822, -19.06564, 
    -18.91273, -18.75951, -18.60596, -18.4521, -18.29792, -18.14341, 
    -17.98859, -17.83344, -17.67798, -17.52219, -17.36608, -17.20966, 
    -17.05291, -16.89584, -16.73845, -16.58074, -16.42271, -16.26436, 
    -16.10569, -15.94669, -15.78738, -15.62775, -15.4678, -15.30752, 
    -15.14693, -14.98602, -14.82479, -14.66324, -14.50137, -14.33918, 
    -14.17667, -14.01384, -13.8507, -13.68723, -13.52346, -13.35936, 
    -13.19494, -13.03021, -12.86517, -12.6998, -12.53412, -12.36813, 
    -12.20182, -12.0352, -11.86826, -11.70101, -11.53345, -11.36558, 
    -11.19739, -11.02889, -10.86009, -10.69097, -10.52154, -10.3518, 
    -10.18176, -10.01141, -9.840751, -9.669786, -9.498516, -9.326941, 
    -9.155064, -8.982882, -8.810398, -8.637612, -8.464526, -8.291141, 
    -8.117455, -7.943473, -7.769193, -7.594616, -7.419745, -7.244579, 
    -7.069119, -6.893368, -6.717325, -6.540992, -6.364369, -6.187459, 
    -6.010261, -5.832778, -5.65501, -5.476958, -5.298624, -5.120009, 
    -4.941114, -4.76194, -4.582489, -4.402761, -4.22276, -4.042484, 
    -3.861936, -3.681118, -3.50003, -3.318675, -3.137053, -2.955165, 
    -2.773015, -2.590602, -2.407929, -2.224997, -2.041807, -1.858361, 
    -1.674662, -1.490709, -1.306506, -1.122053, -0.937353, -0.7524069, 
    -0.5672165, -0.3817838, -0.1961103, -0.010198, 0.1759514, 0.362336, 
    0.5489541, 0.7358036, 0.9228828, 1.11019, 1.297722, 1.485479, 1.673457, 
    1.861656, 2.050072, 2.238704, 2.42755, 2.616607, 2.805874, 2.995349, 
    3.185029, 3.374913, 3.564997, 3.755281, 3.945761, 4.136436, 4.327303, 
    4.51836, 4.709605, 4.901035, 5.092648, 5.284442, 5.476415, 5.668564, 
    5.860887, 6.053381, 6.246044, 6.438873, 6.631867, 6.825022, 7.018336, 
    7.211807, 7.405433, 7.599209, 7.793136, 7.987208, 8.181424, 8.375782, 
    8.570279, 8.764912, 8.959679, 9.154576, 9.349602, 9.544753, 9.740028, 
    9.935423, 10.13093, 10.32656, 10.5223, 10.71815, 10.91411, 11.11017, 
    11.30633, 11.50259, 11.69894, 11.89539, 12.09192, 12.28855, 12.48526, 
    12.68205, 12.87892, 13.07586, 13.27288, 13.46997, 13.66712, 13.86434, 
    14.06162, 14.25896, 14.45636, 14.65381, 14.8513, 15.04885, 15.24644, 
    15.44407, 15.64174, 15.83944, 16.03717, 16.23494, 16.43273, 16.63054, 
    16.82838, 17.02623, 17.2241, 17.42198, 17.61986, 17.81776, 18.01565, 
    18.21355, 18.41144, 18.60933, 18.8072, 19.00507, 19.20292, 19.40075, 
    19.59856, 19.79635, 19.99411, 20.19184, 20.38954, 20.5872, 20.78482, 
    20.9824, 21.17994, 21.37743, 21.57487, 21.77226, 21.96959, 22.16686, 
    22.36407, 22.56121, 22.75829, 22.9553, 23.15223, 23.34909, 23.54586, 
    23.74256, 23.93917, 24.13569, 24.33213, 24.52847, 24.72471, 24.92085, 
    25.1169, 25.31284, 25.50867, 25.70439, 25.9, 26.09549, 26.29087, 
    26.48612, 26.68126, 26.87626, 27.07114, 27.26588, 27.4605, 27.65497, 
    27.84931, 28.0435, 28.23755, 28.43145, 28.62521, 28.81881, 29.01225, 
    29.20554, 29.39867, 29.59164, 29.78444, 29.97708, 30.16955, 30.36184, 
    30.55396, 30.74591, 30.93767, 31.12926, 31.32066, 31.51188, 31.7029, 
    31.89374, 32.08438, 32.27483, 32.46508, 32.65514, 32.84499, 33.03464, 
    33.22408, 33.41331, 33.60234, 33.79115, 33.97975, 34.16813, 34.35629, 
    34.54424, 34.73196, 34.91945, 35.10672, 35.29377, 35.48058, 35.66716, 
    35.85351, 36.03962, 36.2255, 36.41113, 36.59653, 36.78168, 36.96659, 
    37.15125, 37.33566, 37.51982, 37.70374, 37.8874, 38.0708, 38.25395, 
    38.43684, 38.61947, 38.80185, 38.98396, 39.1658, 39.34738, 39.52869, 
    39.70974, 39.89051, 40.07102, 40.25125, 40.43121, 40.61089, 40.7903, 
    40.96943, 41.14828, 41.32685, 41.50514, 41.68315, 41.86087, 42.03831, 
    42.21546, 42.39233, 42.5689, 42.74519, 42.92119, 43.09689, 43.27231, 
    43.44743, 43.62225, 43.79678, 43.97101, 44.14495, 44.31859, 44.49192, 
    44.66496, 44.8377, 45.01014, 45.18227, 45.3541, 45.52563, 45.69685, 
    45.86777, 46.03838, 46.20868, 46.37867, 46.54836, 46.71774, 46.88681, 
    47.05557, 47.22402, 47.39215, 47.55998, 47.72749, 47.89469, 48.06158, 
    48.22815, 48.39441, 48.56035, 48.72598, 48.89129, 49.05629, 49.22097, 
    49.38534, 49.54939, 49.71311,
  -27.62286, -27.48808, -27.35301, -27.21765, -27.08198, -26.94602, 
    -26.80976, -26.67321, -26.53635, -26.39919, -26.26174, -26.12398, 
    -25.98592, -25.84756, -25.70889, -25.56992, -25.43065, -25.29107, 
    -25.15119, -25.011, -24.87051, -24.72971, -24.5886, -24.44718, -24.30545, 
    -24.16342, -24.02108, -23.87842, -23.73546, -23.59218, -23.4486, 
    -23.3047, -23.16049, -23.01597, -22.87113, -22.72598, -22.58052, 
    -22.43474, -22.28864, -22.14224, -21.99551, -21.84847, -21.70111, 
    -21.55344, -21.40545, -21.25714, -21.10852, -20.95957, -20.81031, 
    -20.66073, -20.51083, -20.36061, -20.21007, -20.05921, -19.90803, 
    -19.75653, -19.60471, -19.45257, -19.30011, -19.14733, -18.99422, 
    -18.8408, -18.68705, -18.53298, -18.37859, -18.22388, -18.06884, 
    -17.91348, -17.7578, -17.6018, -17.44547, -17.28883, -17.13186, 
    -16.97456, -16.81695, -16.65901, -16.50075, -16.34217, -16.18326, 
    -16.02403, -15.86448, -15.70461, -15.54441, -15.3839, -15.22306, 
    -15.0619, -14.90041, -14.73861, -14.57649, -14.41404, -14.25127, 
    -14.08819, -13.92478, -13.76105, -13.597, -13.43264, -13.26795, 
    -13.10295, -12.93762, -12.77198, -12.60602, -12.43975, -12.27315, 
    -12.10625, -11.93902, -11.77148, -11.60362, -11.43546, -11.26697, 
    -11.09818, -10.92907, -10.75964, -10.58991, -10.41987, -10.24951, 
    -10.07885, -9.907874, -9.736592, -9.565003, -9.393107, -9.220905, 
    -9.048398, -8.875587, -8.702471, -8.529053, -8.355332, -8.181311, 
    -8.006989, -7.832367, -7.657447, -7.48223, -7.306716, -7.130908, 
    -6.954803, -6.778406, -6.601717, -6.424736, -6.247464, -6.069903, 
    -5.892055, -5.713919, -5.535498, -5.356792, -5.177803, -4.998532, 
    -4.81898, -4.639148, -4.459039, -4.278652, -4.09799, -3.917053, 
    -3.735843, -3.554362, -3.372611, -3.190592, -3.008305, -2.825753, 
    -2.642936, -2.459857, -2.276517, -2.092917, -1.90906, -1.724946, 
    -1.540577, -1.355956, -1.171083, -0.9859605, -0.8005901, -0.6149735, 
    -0.4291126, -0.2430089, -0.0566644, 0.1299191, 0.3167398, 0.5037959, 
    0.6910853, 0.8786063, 1.066357, 1.254335, 1.442539, 1.630967, 1.819617, 
    2.008486, 2.197573, 2.386875, 2.576391, 2.766119, 2.956055, 3.146199, 
    3.336548, 3.5271, 3.717852, 3.908803, 4.09995, 4.291291, 4.482823, 
    4.674545, 4.866454, 5.058548, 5.250824, 5.44328, 5.635914, 5.828723, 
    6.021705, 6.214858, 6.408178, 6.601664, 6.795313, 6.989122, 7.18309, 
    7.377213, 7.571489, 7.765915, 7.96049, 8.15521, 8.350072, 8.545074, 
    8.740213, 8.935489, 9.130895, 9.326431, 9.522094, 9.717881, 9.913789, 
    10.10982, 10.30596, 10.50222, 10.69858, 10.89506, 11.09163, 11.28832, 
    11.4851, 11.68197, 11.87894, 12.076, 12.27315, 12.47039, 12.6677, 
    12.8651, 13.06257, 13.26012, 13.45773, 13.65542, 13.85317, 14.05098, 
    14.24885, 14.44678, 14.64476, 14.84279, 15.04086, 15.23899, 15.43715, 
    15.63535, 15.83359, 16.03186, 16.23016, 16.42848, 16.62683, 16.8252, 
    17.02359, 17.222, 17.42041, 17.61883, 17.81726, 18.01569, 18.21413, 
    18.41255, 18.61098, 18.80939, 19.00779, 19.20617, 19.40454, 19.60289, 
    19.80121, 19.99951, 20.19777, 20.396, 20.5942, 20.79236, 20.99047, 
    21.18854, 21.38656, 21.58454, 21.78245, 21.98031, 22.17812, 22.37586, 
    22.57353, 22.77114, 22.96867, 23.16613, 23.36351, 23.56082, 23.75804, 
    23.95517, 24.15222, 24.34918, 24.54604, 24.7428, 24.93947, 25.13603, 
    25.33249, 25.52884, 25.72507, 25.9212, 26.11721, 26.3131, 26.50887, 
    26.70451, 26.90002, 27.09541, 27.29066, 27.48578, 27.68076, 27.8756, 
    28.0703, 28.26485, 28.45925, 28.6535, 28.8476, 29.04155, 29.23533, 
    29.42895, 29.62241, 29.81571, 30.00883, 30.20179, 30.39457, 30.58718, 
    30.7796, 30.97185, 31.16392, 31.35579, 31.54749, 31.73899, 31.9303, 
    32.12141, 32.31234, 32.50306, 32.69358, 32.88389, 33.07401, 33.26391, 
    33.4536, 33.64309, 33.83235, 34.0214, 34.21024, 34.39885, 34.58725, 
    34.77541, 34.96336, 35.15107, 35.33855, 35.52581, 35.71283, 35.89961, 
    36.08616, 36.27246, 36.45853, 36.64435, 36.82993, 37.01526, 37.20034, 
    37.38518, 37.56976, 37.75409, 37.93816, 38.12198, 38.30553, 38.48883, 
    38.67187, 38.85465, 39.03716, 39.2194, 39.40138, 39.58309, 39.76453, 
    39.94569, 40.12659, 40.30721, 40.48755, 40.66761, 40.8474, 41.02691, 
    41.20613, 41.38508, 41.56374, 41.74212, 41.92021, 42.09801, 42.27552, 
    42.45275, 42.62968, 42.80633, 42.98268, 43.15874, 43.3345, 43.50997, 
    43.68514, 43.86001, 44.03458, 44.20886, 44.38283, 44.5565, 44.72987, 
    44.90294, 45.07571, 45.24817, 45.42032, 45.59217, 45.76371, 45.93494, 
    46.10587, 46.27648, 46.44678, 46.61678, 46.78646, 46.95584, 47.1249, 
    47.29364, 47.46208, 47.6302, 47.798, 47.96549, 48.13267, 48.29953, 
    48.46607, 48.63229, 48.7982, 48.96379, 49.12907, 49.29402, 49.45866, 
    49.62297, 49.78697,
  -27.71361, -27.57873, -27.44355, -27.30808, -27.17231, -27.03624, 
    -26.89987, -26.7632, -26.62623, -26.48896, -26.35139, -26.21351, 
    -26.07534, -25.93685, -25.79807, -25.65898, -25.51958, -25.37987, 
    -25.23986, -25.09954, -24.95892, -24.81799, -24.67674, -24.53519, 
    -24.39333, -24.25116, -24.10867, -23.96588, -23.82277, -23.67935, 
    -23.53562, -23.39157, -23.24721, -23.10254, -22.95755, -22.81224, 
    -22.66662, -22.52069, -22.37443, -22.22786, -22.08098, -21.93377, 
    -21.78625, -21.6384, -21.49025, -21.34176, -21.19297, -21.04385, 
    -20.89441, -20.74465, -20.59457, -20.44416, -20.29344, -20.1424, 
    -19.99103, -19.83934, -19.68733, -19.53499, -19.38234, -19.22936, 
    -19.07605, -18.92243, -18.76848, -18.6142, -18.4596, -18.30468, 
    -18.14944, -17.99387, -17.83797, -17.68175, -17.52521, -17.36834, 
    -17.21115, -17.05363, -16.89579, -16.73762, -16.57913, -16.42032, 
    -16.26118, -16.10171, -15.94192, -15.78181, -15.62137, -15.46061, 
    -15.29952, -15.13811, -14.97638, -14.81432, -14.65194, -14.48924, 
    -14.32621, -14.16287, -13.9992, -13.8352, -13.67089, -13.50625, 
    -13.34129, -13.17601, -13.01041, -12.84449, -12.67826, -12.5117, 
    -12.34482, -12.17762, -12.01011, -11.84228, -11.67413, -11.50566, 
    -11.33688, -11.16778, -10.99837, -10.82865, -10.65861, -10.48825, 
    -10.31759, -10.14661, -9.975322, -9.803722, -9.631813, -9.459596, 
    -9.287069, -9.114235, -8.941094, -8.767648, -8.593896, -8.41984, 
    -8.245481, -8.070819, -7.895855, -7.720592, -7.545028, -7.369165, 
    -7.193005, -7.016548, -6.839795, -6.662748, -6.485407, -6.307773, 
    -6.129848, -5.951633, -5.773129, -5.594337, -5.415258, -5.235894, 
    -5.056245, -4.876314, -4.6961, -4.515606, -4.334833, -4.153783, 
    -3.972456, -3.790854, -3.608978, -3.42683, -3.244411, -3.061723, 
    -2.878768, -2.695546, -2.512059, -2.32831, -2.144298, -1.960027, 
    -1.775497, -1.590711, -1.405669, -1.220374, -1.034828, -0.8490314, 
    -0.6629868, -0.4766957, -0.2901599, -0.1033813, 0.08363826, 0.270897, 
    0.458393, 0.6461244, 0.8340893, 1.022286, 1.210712, 1.399365, 1.588245, 
    1.777347, 1.966672, 2.156216, 2.345977, 2.535954, 2.726144, 2.916544, 
    3.107154, 3.297971, 3.488992, 3.680216, 3.871639, 4.063261, 4.255078, 
    4.447089, 4.63929, 4.83168, 5.024257, 5.217017, 5.409959, 5.603081, 
    5.796379, 5.989851, 6.183496, 6.37731, 6.57129, 6.765436, 6.959743, 
    7.15421, 7.348834, 7.543612, 7.738541, 7.93362, 8.128845, 8.324215, 
    8.519725, 8.715375, 8.91116, 9.107079, 9.303127, 9.499305, 9.695607, 
    9.892032, 10.08858, 10.28524, 10.48201, 10.6789, 10.8759, 11.073, 
    11.2702, 11.46751, 11.66491, 11.8624, 12.05999, 12.25767, 12.45543, 
    12.65328, 12.8512, 13.0492, 13.24728, 13.44543, 13.64365, 13.84193, 
    14.04027, 14.23868, 14.43714, 14.63566, 14.83422, 15.03283, 15.23149, 
    15.43019, 15.62893, 15.82771, 16.02651, 16.22535, 16.42422, 16.6231, 
    16.82201, 17.02094, 17.21988, 17.41883, 17.6178, 17.81677, 18.01574, 
    18.21471, 18.41368, 18.61264, 18.81159, 19.01053, 19.20945, 19.40836, 
    19.60724, 19.8061, 20.00494, 20.20374, 20.40251, 20.60124, 20.79993, 
    20.99859, 21.19719, 21.39575, 21.59426, 21.79271, 21.9911, 22.18944, 
    22.38771, 22.58592, 22.78406, 22.98212, 23.18011, 23.37803, 23.57586, 
    23.77361, 23.97127, 24.16884, 24.36633, 24.56371, 24.761, 24.95819, 
    25.15527, 25.35225, 25.54912, 25.74588, 25.94252, 26.13905, 26.33545, 
    26.53174, 26.72789, 26.92392, 27.11982, 27.31558, 27.51121, 27.7067, 
    27.90205, 28.09725, 28.2923, 28.48721, 28.68196, 28.87656, 29.071, 
    29.26529, 29.45941, 29.65336, 29.84715, 30.04076, 30.23421, 30.42748, 
    30.62057, 30.81349, 31.00622, 31.19876, 31.39112, 31.5833, 31.77528, 
    31.96706, 32.15865, 32.35004, 32.54124, 32.73223, 32.92301, 33.11359, 
    33.30396, 33.49411, 33.68406, 33.87378, 34.06329, 34.25258, 34.44165, 
    34.63049, 34.81911, 35.0075, 35.19566, 35.38359, 35.57128, 35.75874, 
    35.94596, 36.13294, 36.31968, 36.50618, 36.69243, 36.87844, 37.06419, 
    37.2497, 37.43496, 37.61996, 37.8047, 37.98919, 38.17342, 38.35739, 
    38.5411, 38.72454, 38.90773, 39.09064, 39.27328, 39.45566, 39.63776, 
    39.8196, 40.00116, 40.18244, 40.36345, 40.54417, 40.72462, 40.90479, 
    41.08468, 41.26429, 41.4436, 41.62264, 41.80138, 41.97984, 42.15801, 
    42.33589, 42.51348, 42.69077, 42.86777, 43.04448, 43.22089, 43.397, 
    43.57282, 43.74834, 43.92355, 44.09847, 44.27308, 44.44739, 44.6214, 
    44.7951, 44.9685, 45.14159, 45.31438, 45.48686, 45.65903, 45.83089, 
    46.00244, 46.17368, 46.3446, 46.51522, 46.68552, 46.85551, 47.02519, 
    47.19455, 47.3636, 47.53233, 47.70075, 47.86885, 48.03663, 48.20409, 
    48.37124, 48.53807, 48.70457, 48.87076, 49.03663, 49.20218, 49.36741, 
    49.53231, 49.6969, 49.86116,
  -27.80467, -27.66969, -27.53441, -27.39884, -27.26296, -27.12678, -26.9903, 
    -26.85352, -26.71644, -26.57906, -26.44137, -26.30338, -26.16508, 
    -26.02648, -25.88757, -25.74835, -25.60883, -25.469, -25.32886, 
    -25.18842, -25.04766, -24.9066, -24.76522, -24.62353, -24.48153, 
    -24.33922, -24.1966, -24.05366, -23.91041, -23.76685, -23.62297, 
    -23.47878, -23.33427, -23.18944, -23.0443, -22.89884, -22.75307, 
    -22.60697, -22.46056, -22.31383, -22.16678, -22.01941, -21.87172, 
    -21.72371, -21.57538, -21.42673, -21.27776, -21.12846, -20.97885, 
    -20.82891, -20.67864, -20.52806, -20.37715, -20.22592, -20.07437, 
    -19.92249, -19.77029, -19.61776, -19.46491, -19.31173, -19.15823, 
    -19.0044, -18.85025, -18.69577, -18.54096, -18.38583, -18.23038, 
    -18.07459, -17.91849, -17.76205, -17.60529, -17.4482, -17.29078, 
    -17.13304, -16.97497, -16.81658, -16.65786, -16.49881, -16.33944, 
    -16.17973, -16.01971, -15.85935, -15.69867, -15.53766, -15.37633, 
    -15.21467, -15.05269, -14.89038, -14.72774, -14.56478, -14.4015, 
    -14.23789, -14.07395, -13.90969, -13.74511, -13.5802, -13.41497, 
    -13.24942, -13.08354, -12.91735, -12.75083, -12.58398, -12.41682, 
    -12.24934, -12.08153, -11.91341, -11.74497, -11.57621, -11.40713, 
    -11.23773, -11.06801, -10.89798, -10.72763, -10.55697, -10.38599, 
    -10.2147, -10.0431, -9.871179, -9.698949, -9.526408, -9.353557, 
    -9.180395, -9.006925, -8.833146, -8.65906, -8.484668, -8.30997, 
    -8.134967, -7.95966, -7.784051, -7.60814, -7.431927, -7.255414, 
    -7.078603, -6.901494, -6.724088, -6.546386, -6.368389, -6.190099, 
    -6.011516, -5.832642, -5.653477, -5.474024, -5.294283, -5.114256, 
    -4.933943, -4.753346, -4.572467, -4.391307, -4.209867, -4.028147, 
    -3.846151, -3.663879, -3.481333, -3.298514, -3.115423, -2.932063, 
    -2.748434, -2.564538, -2.380377, -2.195952, -2.011265, -1.826318, 
    -1.641112, -1.455649, -1.26993, -1.083958, -0.8977332, -0.7112586, 
    -0.5245355, -0.3375657, -0.1503511, 0.03710651, 0.2248053, 0.4127433, 
    0.6009187, 0.7893294, 0.9779737, 1.166849, 1.355955, 1.545288, 1.734846, 
    1.924628, 2.114631, 2.304853, 2.495293, 2.685947, 2.876815, 3.067893, 
    3.25918, 3.450673, 3.64237, 3.834269, 4.026367, 4.218663, 4.411154, 
    4.603837, 4.796711, 4.989773, 5.18302, 5.376451, 5.570062, 5.763852, 
    5.957818, 6.151957, 6.346266, 6.540745, 6.735389, 6.930197, 7.125165, 
    7.320292, 7.515574, 7.71101, 7.906596, 8.10233, 8.298209, 8.494231, 
    8.690392, 8.886692, 9.083125, 9.27969, 9.476384, 9.673204, 9.870149, 
    10.06721, 10.2644, 10.46169, 10.6591, 10.85662, 11.05425, 11.25198, 
    11.44981, 11.64774, 11.84577, 12.04389, 12.24209, 12.44039, 12.63876, 
    12.83722, 13.03576, 13.23437, 13.43305, 13.63181, 13.83062, 14.02951, 
    14.22845, 14.42745, 14.6265, 14.8256, 15.02476, 15.22396, 15.42319, 
    15.62247, 15.82179, 16.02114, 16.22052, 16.41992, 16.61935, 16.8188, 
    17.01827, 17.21776, 17.41725, 17.61676, 17.81627, 18.01578, 18.21529, 
    18.4148, 18.61431, 18.8138, 19.01328, 19.21275, 19.4122, 19.61162, 
    19.81102, 20.0104, 20.20974, 20.40905, 20.60832, 20.80756, 21.00675, 
    21.20589, 21.40499, 21.60403, 21.80302, 22.00196, 22.20083, 22.39964, 
    22.59838, 22.79705, 22.99565, 23.19418, 23.39262, 23.59099, 23.78927, 
    23.98746, 24.18556, 24.38357, 24.58149, 24.7793, 24.97702, 25.17463, 
    25.37213, 25.56952, 25.7668, 25.96397, 26.16101, 26.35794, 26.55474, 
    26.75141, 26.94796, 27.14437, 27.34065, 27.53679, 27.73278, 27.92864, 
    28.12435, 28.31991, 28.51533, 28.71058, 28.90569, 29.10063, 29.29541, 
    29.49003, 29.68448, 29.87877, 30.07288, 30.26682, 30.46058, 30.65416, 
    30.84756, 31.04078, 31.23381, 31.42665, 31.61931, 31.81177, 32.00403, 
    32.1961, 32.38797, 32.57963, 32.77109, 32.96235, 33.15339, 33.34423, 
    33.53485, 33.72525, 33.91544, 34.10541, 34.29515, 34.48468, 34.67397, 
    34.86304, 35.05188, 35.24049, 35.42886, 35.617, 35.8049, 35.99256, 
    36.17998, 36.36716, 36.55409, 36.74077, 36.92721, 37.11339, 37.29932, 
    37.485, 37.67043, 37.85559, 38.0405, 38.22514, 38.40953, 38.59364, 
    38.7775, 38.96109, 39.1444, 39.32745, 39.51023, 39.69273, 39.87496, 
    40.05691, 40.23859, 40.41998, 40.6011, 40.78193, 40.96249, 41.14275, 
    41.32273, 41.50243, 41.68184, 41.86095, 42.03978, 42.21832, 42.39656, 
    42.57452, 42.75217, 42.92953, 43.10659, 43.28336, 43.45982, 43.63599, 
    43.81185, 43.98741, 44.16267, 44.33762, 44.51228, 44.68662, 44.86066, 
    45.03439, 45.20781, 45.38092, 45.55372, 45.72622, 45.8984, 46.07026, 
    46.24182, 46.41306, 46.58399, 46.7546, 46.9249, 47.09488, 47.26455, 
    47.43389, 47.60292, 47.77163, 47.94003, 48.1081, 48.27585, 48.44328, 
    48.6104, 48.77719, 48.94366, 49.10981, 49.27563, 49.44113, 49.60631, 
    49.77117, 49.9357,
  -27.89606, -27.76098, -27.6256, -27.48991, -27.35393, -27.21764, -27.08106, 
    -26.94416, -26.80697, -26.66947, -26.53167, -26.39356, -26.25515, 
    -26.11642, -25.97739, -25.83806, -25.69841, -25.55846, -25.41819, 
    -25.27762, -25.13673, -24.99554, -24.85403, -24.71221, -24.57007, 
    -24.42762, -24.28486, -24.14178, -23.99839, -23.85468, -23.71066, 
    -23.56632, -23.42166, -23.27669, -23.13139, -22.98578, -22.83985, 
    -22.6936, -22.54702, -22.40013, -22.25292, -22.10539, -21.95753, 
    -21.80935, -21.66085, -21.51203, -21.36289, -21.21342, -21.06363, 
    -20.91351, -20.76307, -20.6123, -20.46121, -20.30979, -20.15805, 
    -20.00598, -19.85359, -19.70087, -19.54782, -19.39445, -19.24075, 
    -19.08672, -18.93236, -18.77768, -18.62267, -18.46733, -18.31166, 
    -18.15567, -17.99934, -17.84269, -17.68571, -17.5284, -17.37077, 
    -17.2128, -17.0545, -16.89588, -16.73693, -16.57765, -16.41804, -16.2581, 
    -16.09784, -15.93724, -15.77632, -15.61507, -15.45349, -15.29158, 
    -15.12934, -14.96678, -14.80389, -14.64067, -14.47712, -14.31325, 
    -14.14905, -13.98453, -13.81968, -13.6545, -13.489, -13.32317, -13.15701, 
    -12.99054, -12.82374, -12.65661, -12.48916, -12.32139, -12.1533, 
    -11.98488, -11.81614, -11.64708, -11.4777, -11.30801, -11.13799, 
    -10.96765, -10.79699, -10.62602, -10.45473, -10.28312, -10.1112, 
    -9.938964, -9.766413, -9.593548, -9.42037, -9.246881, -9.073079, 
    -8.898968, -8.724547, -8.549817, -8.37478, -8.199435, -8.023784, 
    -7.847828, -7.671568, -7.495005, -7.318139, -7.140972, -6.963505, 
    -6.785739, -6.607675, -6.429314, -6.250657, -6.071705, -5.892459, 
    -5.712922, -5.533093, -5.352974, -5.172566, -4.991871, -4.81089, 
    -4.629624, -4.448075, -4.266243, -4.084131, -3.901739, -3.719069, 
    -3.536123, -3.352901, -3.169406, -2.985639, -2.801602, -2.617295, 
    -2.432721, -2.247881, -2.062778, -1.877411, -1.691783, -1.505897, 
    -1.319752, -1.133352, -0.9466979, -0.7597914, -0.5726344, -0.3852287, 
    -0.1975761, -0.009678453, 0.1784623, 0.3668443, 0.5554657, 0.7443244, 
    0.9334186, 1.122746, 1.312305, 1.502094, 1.69211, 1.882351, 2.072816, 
    2.263501, 2.454406, 2.645528, 2.836864, 3.028413, 3.220172, 3.412139, 
    3.604312, 3.796689, 3.989266, 4.182044, 4.375017, 4.568185, 4.761545, 
    4.955094, 5.148831, 5.342753, 5.536857, 5.731141, 5.925601, 6.120238, 
    6.315046, 6.510025, 6.705171, 6.900482, 7.095955, 7.291588, 7.487378, 
    7.683322, 7.879418, 8.075664, 8.272055, 8.468591, 8.665267, 8.862082, 
    9.059033, 9.256117, 9.453331, 9.650673, 9.848139, 10.04573, 10.24343, 
    10.44126, 10.63919, 10.83724, 11.0354, 11.23366, 11.43202, 11.63048, 
    11.82904, 12.02769, 12.22643, 12.42526, 12.62417, 12.82316, 13.02224, 
    13.22138, 13.42061, 13.6199, 13.81925, 14.01868, 14.21816, 14.4177, 
    14.61729, 14.81694, 15.01663, 15.21637, 15.41616, 15.61598, 15.81584, 
    16.01573, 16.21565, 16.4156, 16.61558, 16.81557, 17.01559, 17.21562, 
    17.41566, 17.61571, 17.81576, 18.01582, 18.21588, 18.41594, 18.61599, 
    18.81602, 19.01605, 19.21606, 19.41606, 19.61603, 19.81597, 20.01589, 
    20.21578, 20.41563, 20.61545, 20.81523, 21.01496, 21.21465, 21.41428, 
    21.61387, 21.8134, 22.01287, 22.21229, 22.41163, 22.61091, 22.81012, 
    23.00926, 23.20832, 23.4073, 23.6062, 23.80502, 24.00374, 24.20238, 
    24.40092, 24.59937, 24.79771, 24.99596, 25.19409, 25.39212, 25.59004, 
    25.78785, 25.98554, 26.18311, 26.38055, 26.57787, 26.77507, 26.97213, 
    27.16906, 27.36585, 27.56251, 27.75902, 27.95539, 28.15161, 28.34768, 
    28.5436, 28.73937, 28.93498, 29.13042, 29.32571, 29.52083, 29.71578, 
    29.91056, 30.10517, 30.2996, 30.49386, 30.68793, 30.88183, 31.07553, 
    31.26905, 31.46238, 31.65552, 31.84846, 32.04121, 32.23376, 32.4261, 
    32.61824, 32.81018, 33.0019, 33.19342, 33.38472, 33.57581, 33.76668, 
    33.95733, 34.14776, 34.33796, 34.52794, 34.71769, 34.90722, 35.09651, 
    35.28556, 35.47439, 35.66297, 35.85131, 36.03942, 36.22728, 36.41489, 
    36.60226, 36.78938, 36.97624, 37.16285, 37.34921, 37.53532, 37.72116, 
    37.90675, 38.09208, 38.27714, 38.46194, 38.64647, 38.83073, 39.01472, 
    39.19845, 39.3819, 39.56508, 39.74798, 39.93061, 40.11296, 40.29502, 
    40.47681, 40.65832, 40.83954, 41.02047, 41.20112, 41.38148, 41.56156, 
    41.74134, 41.92083, 42.10003, 42.27894, 42.45755, 42.63586, 42.81388, 
    42.9916, 43.16902, 43.34614, 43.52295, 43.69947, 43.87568, 44.05159, 
    44.22719, 44.40249, 44.57748, 44.75216, 44.92653, 45.10059, 45.27435, 
    45.44778, 45.62091, 45.79373, 45.96623, 46.13842, 46.31029, 46.48185, 
    46.65309, 46.82401, 46.99461, 47.1649, 47.33487, 47.50452, 47.67385, 
    47.84285, 48.01154, 48.17991, 48.34795, 48.51567, 48.68307, 48.85014, 
    49.01689, 49.18332, 49.34942, 49.5152, 49.68065, 49.84578, 50.01057,
  -27.98777, -27.85258, -27.7171, -27.58131, -27.44522, -27.30883, -27.17213, 
    -27.03513, -26.89783, -26.76022, -26.6223, -26.48407, -26.34554, 
    -26.2067, -26.06755, -25.92809, -25.78833, -25.64825, -25.50786, 
    -25.36716, -25.22614, -25.08481, -24.94317, -24.80122, -24.65895, 
    -24.51636, -24.37346, -24.23024, -24.08671, -23.94286, -23.79869, 
    -23.6542, -23.50939, -23.36427, -23.21882, -23.07306, -22.92697, 
    -22.78056, -22.63383, -22.48678, -22.33941, -22.19171, -22.04369, 
    -21.89534, -21.74668, -21.59768, -21.44836, -21.29872, -21.14875, 
    -20.99846, -20.84784, -20.69689, -20.54561, -20.39401, -20.24208, 
    -20.08982, -19.93724, -19.78433, -19.63108, -19.47751, -19.32361, 
    -19.16938, -19.01483, -18.85994, -18.70472, -18.54917, -18.3933, 
    -18.23709, -18.08055, -17.92368, -17.76649, -17.60896, -17.4511, 
    -17.29291, -17.13438, -16.97553, -16.81635, -16.65684, -16.49699, 
    -16.33682, -16.17631, -16.01548, -15.85431, -15.69281, -15.53099, 
    -15.36883, -15.20634, -15.04353, -14.88038, -14.7169, -14.5531, 
    -14.38896, -14.2245, -14.05971, -13.89459, -13.72914, -13.56336, 
    -13.39726, -13.23083, -13.06407, -12.89699, -12.72958, -12.56184, 
    -12.39378, -12.2254, -12.05669, -11.88766, -11.7183, -11.54862, 
    -11.37862, -11.2083, -11.03765, -10.86669, -10.6954, -10.5238, -10.35188, 
    -10.17964, -10.00708, -9.834208, -9.661018, -9.487514, -9.313695, 
    -9.139562, -8.965117, -8.790359, -8.615292, -8.439914, -8.264226, 
    -8.08823, -7.911927, -7.735317, -7.558401, -7.381181, -7.203658, 
    -7.025832, -6.847705, -6.669277, -6.49055, -6.311525, -6.132203, 
    -5.952585, -5.772673, -5.592467, -5.411969, -5.23118, -5.050101, 
    -4.868734, -4.68708, -4.50514, -4.322916, -4.140408, -3.957619, -3.77455, 
    -3.591202, -3.407577, -3.223676, -3.039501, -2.855053, -2.670334, 
    -2.485345, -2.300089, -2.114566, -1.928778, -1.742727, -1.556415, 
    -1.369843, -1.183014, -0.9959278, -0.8085876, -0.6209947, -0.4331511, 
    -0.2450586, -0.05671899, 0.1318658, 0.3206938, 0.5097632, 0.699072, 
    0.8886182, 1.0784, 1.268415, 1.458661, 1.649137, 1.83984, 2.030768, 
    2.22192, 2.413291, 2.604882, 2.79669, 2.988711, 3.180945, 3.373389, 
    3.56604, 3.758897, 3.951957, 4.145217, 4.338676, 4.532331, 4.72618, 
    4.920219, 5.114448, 5.308863, 5.503462, 5.698243, 5.893202, 6.088338, 
    6.283648, 6.47913, 6.67478, 6.870597, 7.066577, 7.262719, 7.459018, 
    7.655474, 7.852083, 8.048842, 8.245749, 8.442802, 8.639997, 8.837331, 
    9.034802, 9.232408, 9.430145, 9.62801, 9.826001, 10.02412, 10.22235, 
    10.4207, 10.61917, 10.81775, 11.01643, 11.21522, 11.41412, 11.61311, 
    11.81221, 12.01139, 12.21067, 12.41004, 12.60949, 12.80902, 13.00863, 
    13.20832, 13.40808, 13.60792, 13.80782, 14.00778, 14.20781, 14.40789, 
    14.60803, 14.80822, 15.00846, 15.20875, 15.40908, 15.60945, 15.80985, 
    16.01029, 16.21076, 16.41126, 16.61178, 16.81233, 17.01289, 17.21347, 
    17.41405, 17.61465, 17.81526, 18.01587, 18.21647, 18.41708, 18.61768, 
    18.81826, 19.01884, 19.2194, 19.41994, 19.62046, 19.82095, 20.02142, 
    20.22185, 20.42225, 20.62262, 20.82294, 21.02322, 21.22345, 21.42363, 
    21.62376, 21.82384, 22.02386, 22.22381, 22.4237, 22.62352, 22.82327, 
    23.02295, 23.22255, 23.42207, 23.62151, 23.82086, 24.02012, 24.21929, 
    24.41837, 24.61735, 24.81623, 25.01501, 25.21367, 25.41223, 25.61068, 
    25.80902, 26.00723, 26.20533, 26.4033, 26.60114, 26.79886, 26.99644, 
    27.19389, 27.3912, 27.58838, 27.78541, 27.98229, 28.17903, 28.37561, 
    28.57204, 28.76832, 28.96444, 29.16039, 29.35618, 29.5518, 29.74726, 
    29.94254, 30.13765, 30.33258, 30.52733, 30.7219, 30.91629, 31.11049, 
    31.3045, 31.49832, 31.69194, 31.88537, 32.07859, 32.27162, 32.46445, 
    32.65707, 32.84948, 33.04168, 33.23367, 33.42544, 33.617, 33.80833, 
    33.99945, 34.19034, 34.38101, 34.57145, 34.76166, 34.95164, 35.14138, 
    35.33089, 35.52016, 35.70919, 35.89798, 36.08653, 36.27483, 36.46288, 
    36.65068, 36.83824, 37.02554, 37.21259, 37.39937, 37.5859, 37.77217, 
    37.95818, 38.14393, 38.32941, 38.51463, 38.69957, 38.88425, 39.06865, 
    39.25278, 39.43664, 39.62022, 39.80353, 39.98655, 40.1693, 40.35176, 
    40.53394, 40.71583, 40.89744, 41.07877, 41.2598, 41.44054, 41.62099, 
    41.80115, 41.98102, 42.16059, 42.33986, 42.51884, 42.69752, 42.8759, 
    43.05398, 43.23176, 43.40923, 43.58641, 43.76328, 43.93983, 44.11609, 
    44.29204, 44.46767, 44.64301, 44.81802, 44.99273, 45.16713, 45.34121, 
    45.51498, 45.68843, 45.86158, 46.0344, 46.20691, 46.3791, 46.55097, 
    46.72252, 46.89375, 47.06467, 47.23526, 47.40553, 47.57548, 47.74511, 
    47.91442, 48.0834, 48.25206, 48.42039, 48.5884, 48.75608, 48.92344, 
    49.09047, 49.25718, 49.42356, 49.58961, 49.75533, 49.92073, 50.0858,
  -28.0798, -27.94452, -27.80893, -27.67304, -27.53684, -27.40034, -27.26354, 
    -27.12643, -26.98901, -26.85129, -26.71326, -26.57492, -26.43627, 
    -26.29731, -26.15804, -26.01846, -25.87857, -25.73837, -25.59785, 
    -25.45703, -25.31588, -25.17443, -25.03265, -24.89056, -24.74816, 
    -24.60544, -24.4624, -24.31904, -24.17537, -24.03137, -23.88706, 
    -23.74242, -23.59747, -23.45219, -23.3066, -23.16068, -23.01443, 
    -22.86787, -22.72098, -22.57377, -22.42624, -22.27838, -22.13019, 
    -21.98168, -21.83284, -21.68368, -21.53419, -21.38437, -21.23422, 
    -21.08375, -20.93295, -20.78182, -20.63037, -20.47858, -20.32646, 
    -20.17402, -20.02124, -19.86813, -19.7147, -19.56093, -19.40683, 
    -19.2524, -19.09764, -18.94255, -18.78712, -18.63137, -18.47528, 
    -18.31886, -18.16211, -18.00503, -17.84761, -17.68986, -17.53178, 
    -17.37336, -17.21461, -17.05553, -16.89612, -16.73638, -16.5763, 
    -16.41589, -16.25514, -16.09406, -15.93266, -15.77091, -15.60884, 
    -15.44643, -15.28369, -15.12062, -14.95722, -14.79349, -14.62942, 
    -14.46502, -14.30029, -14.13524, -13.96985, -13.80413, -13.63808, 
    -13.4717, -13.30499, -13.13795, -12.97059, -12.80289, -12.63487, 
    -12.46652, -12.29784, -12.12884, -11.95951, -11.78986, -11.61988, 
    -11.44957, -11.27895, -11.108, -10.93672, -10.76513, -10.59321, 
    -10.42097, -10.24841, -10.07553, -9.902336, -9.728822, -9.554989, 
    -9.38084, -9.206375, -9.031595, -8.856502, -8.681094, -8.505374, 
    -8.329343, -8.153, -7.976348, -7.799388, -7.622119, -7.444544, -7.266663, 
    -7.088477, -6.909987, -6.731195, -6.552101, -6.372707, -6.193014, 
    -6.013022, -5.832734, -5.652149, -5.471271, -5.290099, -5.108635, 
    -4.92688, -4.744836, -4.562504, -4.379886, -4.196982, -4.013794, 
    -3.830324, -3.646574, -3.462543, -3.278235, -3.09365, -2.90879, 
    -2.723657, -2.538252, -2.352576, -2.166633, -1.980422, -1.793946, 
    -1.607207, -1.420206, -1.232945, -1.045426, -0.8576496, -0.669619, 
    -0.4813355, -0.2928011, -0.1040175, 0.08501332, 0.2742895, 0.463809, 
    0.6535699, 0.8435702, 1.033808, 1.224281, 1.414988, 1.605925, 1.797092, 
    1.988486, 2.180105, 2.371947, 2.564009, 2.75629, 2.948787, 3.141498, 
    3.334421, 3.527553, 3.720892, 3.914436, 4.108183, 4.302129, 4.496274, 
    4.690613, 4.885146, 5.079869, 5.27478, 5.469877, 5.665157, 5.860618, 
    6.056256, 6.25207, 6.448057, 6.644215, 6.840539, 7.03703, 7.233683, 
    7.430496, 7.627466, 7.82459, 8.021867, 8.219292, 8.416863, 8.614579, 
    8.812436, 9.01043, 9.208561, 9.406823, 9.605216, 9.803735, 10.00238, 
    10.20114, 10.40003, 10.59902, 10.79814, 10.99736, 11.19668, 11.39612, 
    11.59565, 11.79528, 11.995, 12.19482, 12.39473, 12.59472, 12.79479, 
    12.99495, 13.19518, 13.39549, 13.59587, 13.79631, 13.99682, 14.19739, 
    14.39803, 14.59871, 14.79945, 15.00024, 15.20108, 15.40195, 15.60287, 
    15.80383, 16.00482, 16.20584, 16.40689, 16.60796, 16.80906, 17.01017, 
    17.2113, 17.41244, 17.61359, 17.81475, 18.01591, 18.21707, 18.41823, 
    18.61938, 18.82051, 19.02164, 19.22275, 19.42385, 19.62491, 19.82596, 
    20.02698, 20.22796, 20.42891, 20.62983, 20.8307, 21.03152, 21.23231, 
    21.43304, 21.63371, 21.83434, 22.0349, 22.2354, 22.43583, 22.6362, 
    22.8365, 23.03672, 23.23686, 23.43692, 23.6369, 23.83679, 24.0366, 
    24.23631, 24.43592, 24.63544, 24.83485, 25.03416, 25.23337, 25.43246, 
    25.63144, 25.83031, 26.02905, 26.22768, 26.42618, 26.62455, 26.82279, 
    27.0209, 27.21887, 27.41671, 27.6144, 27.81195, 28.00935, 28.2066, 
    28.4037, 28.60065, 28.79744, 28.99406, 29.19053, 29.38683, 29.58296, 
    29.77892, 29.9747, 30.17031, 30.36575, 30.561, 30.75606, 30.95094, 
    31.14564, 31.34014, 31.53445, 31.72856, 31.92248, 32.11619, 32.3097, 
    32.50301, 32.69611, 32.889, 33.08168, 33.27414, 33.46638, 33.65841, 
    33.85022, 34.04181, 34.23316, 34.42429, 34.6152, 34.80586, 34.9963, 
    35.1865, 35.37646, 35.56618, 35.75567, 35.9449, 36.1339, 36.32264, 
    36.51114, 36.69938, 36.88737, 37.0751, 37.26258, 37.4498, 37.63676, 
    37.82346, 38.0099, 38.19606, 38.38197, 38.5676, 38.75296, 38.93805, 
    39.12287, 39.30741, 39.49167, 39.67566, 39.85936, 40.04279, 40.22593, 
    40.40879, 40.59137, 40.77365, 40.95565, 41.13736, 41.31878, 41.4999, 
    41.68073, 41.86127, 42.04152, 42.22146, 42.4011, 42.58045, 42.7595, 
    42.93824, 43.11668, 43.29482, 43.47265, 43.65018, 43.8274, 44.00431, 
    44.18092, 44.35721, 44.53319, 44.70886, 44.88422, 45.05927, 45.23399, 
    45.40841, 45.58251, 45.75629, 45.92976, 46.1029, 46.27573, 46.44824, 
    46.62043, 46.79229, 46.96384, 47.13506, 47.30596, 47.47654, 47.64679, 
    47.81672, 47.98632, 48.1556, 48.32455, 48.49317, 48.66147, 48.82944, 
    48.99708, 49.16439, 49.33138, 49.49804, 49.66436, 49.83036, 49.99603, 
    50.16137,
  -28.17216, -28.03677, -27.90108, -27.76509, -27.62879, -27.49218, 
    -27.35527, -27.21805, -27.08053, -26.94269, -26.80455, -26.66609, 
    -26.52733, -26.38825, -26.24887, -26.10917, -25.96915, -25.82883, 
    -25.68819, -25.54723, -25.40596, -25.26437, -25.12247, -24.98025, 
    -24.83771, -24.69485, -24.55168, -24.40818, -24.26436, -24.12023, 
    -23.97577, -23.83099, -23.68589, -23.54046, -23.39471, -23.24864, 
    -23.10225, -22.95553, -22.80848, -22.66111, -22.51341, -22.36539, 
    -22.21704, -22.06836, -21.91936, -21.77002, -21.62036, -21.47037, 
    -21.32005, -21.1694, -21.01842, -20.86711, -20.71547, -20.5635, 
    -20.41119, -20.25856, -20.10559, -19.95229, -19.79866, -19.6447, 
    -19.4904, -19.33577, -19.18081, -19.02551, -18.86988, -18.71392, 
    -18.55762, -18.40099, -18.24402, -18.08672, -17.92909, -17.77112, 
    -17.61281, -17.45417, -17.2952, -17.13589, -16.97625, -16.81627, 
    -16.65595, -16.49531, -16.33432, -16.17301, -16.01135, -15.84937, 
    -15.68704, -15.52439, -15.3614, -15.19807, -15.03441, -14.87042, 
    -14.70609, -14.54143, -14.37644, -14.21111, -14.04545, -13.87946, 
    -13.71314, -13.54648, -13.3795, -13.21218, -13.04453, -12.87655, 
    -12.70824, -12.5396, -12.37064, -12.20134, -12.03171, -11.86176, 
    -11.69148, -11.52087, -11.34994, -11.17868, -11.0071, -10.83519, 
    -10.66296, -10.4904, -10.31752, -10.14432, -9.970802, -9.796961, 
    -9.622799, -9.448319, -9.273521, -9.098406, -8.922974, -8.747226, 
    -8.571164, -8.394788, -8.218098, -8.041097, -7.863784, -7.686162, 
    -7.50823, -7.32999, -7.151443, -6.972589, -6.793432, -6.61397, -6.434205, 
    -6.254139, -6.073772, -5.893106, -5.712142, -5.530882, -5.349326, 
    -5.167475, -4.985332, -4.802897, -4.620172, -4.437158, -4.253856, 
    -4.070268, -3.886395, -3.70224, -3.517802, -3.333085, -3.148088, 
    -2.962815, -2.777266, -2.591443, -2.405347, -2.218981, -2.032346, 
    -1.845443, -1.658275, -1.470843, -1.283148, -1.095193, -0.9069799, 
    -0.7185096, -0.5297843, -0.3408059, -0.1515764, 0.03790253, 0.2276288, 
    0.4176005, 0.6078156, 0.7982723, 0.9889683, 1.179902, 1.371071, 1.562472, 
    1.754106, 1.945968, 2.138057, 2.330371, 2.522907, 2.715663, 2.908638, 
    3.101828, 3.295232, 3.488848, 3.682672, 3.876703, 4.070938, 4.265375, 
    4.460011, 4.654844, 4.849872, 5.045093, 5.240502, 5.4361, 5.631882, 
    5.827846, 6.023989, 6.22031, 6.416805, 6.613472, 6.810309, 7.007312, 
    7.204479, 7.401807, 7.599295, 7.796937, 7.994734, 8.19268, 8.390775, 
    8.589014, 8.787395, 8.985917, 9.184574, 9.383366, 9.582288, 9.781339, 
    9.980514, 10.17981, 10.37923, 10.57876, 10.77841, 10.97817, 11.17803, 
    11.37801, 11.57808, 11.77825, 11.97852, 12.17888, 12.37933, 12.57986, 
    12.78048, 12.98119, 13.18196, 13.38282, 13.58374, 13.78474, 13.9858, 
    14.18692, 14.3881, 14.58934, 14.79063, 14.99197, 15.19336, 15.39479, 
    15.59626, 15.79777, 15.99932, 16.20089, 16.40249, 16.60412, 16.80577, 
    17.00744, 17.20913, 17.41082, 17.61253, 17.81424, 18.01595, 18.21767, 
    18.41938, 18.62108, 18.82278, 19.02446, 19.22613, 19.42777, 19.6294, 
    19.831, 20.03257, 20.23411, 20.43561, 20.63708, 20.8385, 21.03988, 
    21.24121, 21.4425, 21.64373, 21.8449, 22.04601, 22.24706, 22.44804, 
    22.64896, 22.8498, 23.05057, 23.25126, 23.45186, 23.65239, 23.85282, 
    24.05317, 24.25342, 24.45358, 24.65363, 24.85359, 25.05344, 25.25318, 
    25.45281, 25.65232, 25.85172, 26.051, 26.25016, 26.44919, 26.64809, 
    26.84686, 27.0455, 27.24399, 27.44235, 27.64057, 27.83864, 28.03656, 
    28.23434, 28.43196, 28.62942, 28.82672, 29.02386, 29.22084, 29.41765, 
    29.61429, 29.81076, 30.00705, 30.20317, 30.3991, 30.59485, 30.79042, 
    30.9858, 31.18099, 31.37599, 31.57079, 31.7654, 31.9598, 32.154, 32.348, 
    32.54179, 32.73537, 32.92875, 33.1219, 33.31484, 33.50756, 33.70007, 
    33.89235, 34.0844, 34.27622, 34.46782, 34.65918, 34.85032, 35.04121, 
    35.23187, 35.42229, 35.61246, 35.8024, 35.99209, 36.18153, 36.37072, 
    36.55965, 36.74834, 36.93677, 37.12494, 37.31285, 37.50051, 37.6879, 
    37.87503, 38.06189, 38.24848, 38.4348, 38.62085, 38.80663, 38.99214, 
    39.17737, 39.36232, 39.547, 39.73139, 39.9155, 40.09933, 40.28287, 
    40.46613, 40.64909, 40.83178, 41.01416, 41.19626, 41.37806, 41.55957, 
    41.74079, 41.9217, 42.10232, 42.28264, 42.46266, 42.64238, 42.82179, 
    43.0009, 43.17971, 43.3582, 43.5364, 43.71428, 43.89185, 44.06911, 
    44.24607, 44.42271, 44.59903, 44.77505, 44.95074, 45.12613, 45.30119, 
    45.47594, 45.65037, 45.82448, 45.99827, 46.17174, 46.34489, 46.51772, 
    46.69022, 46.8624, 47.03426, 47.20579, 47.377, 47.54788, 47.71844, 
    47.88866, 48.05857, 48.22814, 48.39738, 48.5663, 48.73489, 48.90314, 
    49.07107, 49.23867, 49.40593, 49.57287, 49.73947, 49.90574, 50.07168, 
    50.23729,
  -28.26484, -28.12935, -27.99356, -27.85747, -27.72106, -27.58435, 
    -27.44734, -27.31001, -27.17237, -27.03443, -26.89617, -26.7576, 
    -26.61872, -26.47953, -26.34003, -26.20021, -26.06007, -25.91962, 
    -25.77886, -25.63778, -25.49638, -25.35466, -25.21263, -25.07028, 
    -24.9276, -24.78461, -24.6413, -24.49766, -24.3537, -24.20943, -24.06483, 
    -23.9199, -23.77465, -23.62908, -23.48318, -23.33696, -23.19041, 
    -23.04353, -22.89633, -22.7488, -22.60094, -22.45275, -22.30424, 
    -22.1554, -22.00622, -21.85672, -21.70688, -21.55672, -21.40623, 
    -21.2554, -21.10424, -20.95275, -20.80092, -20.64877, -20.49628, 
    -20.34345, -20.1903, -20.03681, -19.88298, -19.72882, -19.57433, 
    -19.4195, -19.26433, -19.10883, -18.953, -18.79683, -18.64032, -18.48347, 
    -18.32629, -18.16878, -18.01092, -17.85273, -17.69421, -17.53534, 
    -17.37614, -17.2166, -17.05673, -16.89652, -16.73597, -16.57508, 
    -16.41386, -16.2523, -16.09041, -15.92817, -15.7656, -15.6027, -15.43945, 
    -15.27588, -15.11196, -14.94771, -14.78312, -14.6182, -14.45294, 
    -14.28735, -14.12142, -13.95515, -13.78856, -13.62162, -13.45436, 
    -13.28676, -13.11883, -12.95056, -12.78197, -12.61304, -12.44378, 
    -12.27418, -12.10426, -11.93401, -11.76343, -11.59252, -11.42128, 
    -11.24971, -11.07782, -10.90559, -10.73305, -10.56017, -10.38697, 
    -10.21345, -10.03961, -9.865438, -9.690948, -9.516135, -9.341003, 
    -9.165551, -8.98978, -8.813692, -8.637286, -8.460564, -8.283525, 
    -8.106174, -7.928509, -7.750531, -7.572241, -7.393641, -7.214732, 
    -7.035514, -6.855989, -6.676158, -6.496022, -6.315582, -6.134839, 
    -5.953794, -5.772449, -5.590806, -5.408864, -5.226625, -5.044092, 
    -4.861264, -4.678144, -4.494732, -4.311031, -4.127042, -3.942765, 
    -3.758203, -3.573357, -3.388229, -3.20282, -3.017131, -2.831164, 
    -2.644921, -2.458404, -2.271613, -2.084552, -1.89722, -1.709621, 
    -1.521756, -1.333626, -1.145234, -0.956581, -0.767669, -0.5785, 
    -0.3890757, -0.1993981, -0.009469034, 0.1807095, 0.3711354, 0.5618069, 
    0.7527219, 0.9438784, 1.135274, 1.326908, 1.518776, 1.710878, 1.90321, 
    2.095772, 2.28856, 2.481572, 2.674807, 2.868261, 3.061934, 3.255821, 
    3.449922, 3.644234, 3.838754, 4.03348, 4.22841, 4.423541, 4.61887, 
    4.814396, 5.010116, 5.206028, 5.402128, 5.598414, 5.794885, 5.991536, 
    6.188366, 6.385373, 6.582552, 6.779903, 6.977422, 7.175106, 7.372952, 
    7.57096, 7.769124, 7.967443, 8.165914, 8.364533, 8.563299, 8.762209, 
    8.961259, 9.160447, 9.35977, 9.559225, 9.75881, 9.958521, 10.15835, 
    10.35831, 10.55838, 10.75857, 10.95887, 11.15928, 11.35979, 11.5604, 
    11.76112, 11.96193, 12.16284, 12.36384, 12.56492, 12.76609, 12.96734, 
    13.16867, 13.37007, 13.57155, 13.7731, 13.97471, 14.17638, 14.37812, 
    14.57991, 14.78176, 14.98365, 15.18559, 15.38758, 15.58961, 15.79168, 
    15.99378, 16.19591, 16.39807, 16.60026, 16.80247, 17.00469, 17.20693, 
    17.40919, 17.61145, 17.81372, 18.016, 18.21827, 18.42054, 18.6228, 
    18.82506, 19.0273, 19.22952, 19.43173, 19.63391, 19.83607, 20.03819, 
    20.24029, 20.44235, 20.64437, 20.84635, 21.04829, 21.25018, 21.45201, 
    21.6538, 21.85552, 22.05719, 22.25879, 22.46033, 22.66179, 22.86318, 
    23.0645, 23.26574, 23.46689, 23.66796, 23.86895, 24.06984, 24.27064, 
    24.47134, 24.67194, 24.87243, 25.07282, 25.27311, 25.47327, 25.67333, 
    25.87326, 26.07308, 26.27277, 26.47233, 26.67177, 26.87107, 27.07024, 
    27.26926, 27.46815, 27.66689, 27.86549, 28.06394, 28.26223, 28.46037, 
    28.65835, 28.85618, 29.05383, 29.25133, 29.44865, 29.6458, 29.84278, 
    30.03958, 30.23621, 30.43265, 30.6289, 30.82498, 31.02086, 31.21655, 
    31.41204, 31.60734, 31.80244, 31.99734, 32.19203, 32.38652, 32.5808, 
    32.77486, 32.96872, 33.16235, 33.35577, 33.54897, 33.74195, 33.9347, 
    34.12723, 34.31953, 34.51159, 34.70342, 34.89502, 35.08638, 35.27749, 
    35.46837, 35.659, 35.84939, 36.03953, 36.22942, 36.41906, 36.60844, 
    36.79757, 36.98644, 37.17505, 37.3634, 37.55149, 37.73932, 37.92687, 
    38.11416, 38.30118, 38.48793, 38.6744, 38.8606, 39.04652, 39.23217, 
    39.41753, 39.60262, 39.78742, 39.97194, 40.15617, 40.34011, 40.52377, 
    40.70713, 40.89021, 41.07299, 41.25547, 41.43766, 41.61956, 41.80116, 
    41.98245, 42.16345, 42.34414, 42.52454, 42.70462, 42.88441, 43.06388, 
    43.24305, 43.42191, 43.60046, 43.77871, 43.95663, 44.13425, 44.31155, 
    44.48854, 44.66521, 44.84157, 45.0176, 45.19333, 45.36873, 45.54381, 
    45.71857, 45.89301, 46.06713, 46.24092, 46.41439, 46.58754, 46.76036, 
    46.93286, 47.10503, 47.27687, 47.44839, 47.61958, 47.79043, 47.96096, 
    48.13116, 48.30103, 48.47057, 48.63978, 48.80866, 48.9772, 49.14541, 
    49.31329, 49.48084, 49.64805, 49.81493, 49.98148, 50.14769, 50.31356,
  -28.35785, -28.22227, -28.08638, -27.95018, -27.81367, -27.67686, 
    -27.53973, -27.4023, -27.26455, -27.1265, -26.98813, -26.84945, 
    -26.71046, -26.57115, -26.43153, -26.29159, -26.15133, -26.01076, 
    -25.86987, -25.72867, -25.58714, -25.4453, -25.30313, -25.16065, 
    -25.01784, -24.87471, -24.73126, -24.58749, -24.44339, -24.29897, 
    -24.15423, -24.00916, -23.86376, -23.71804, -23.57199, -23.42562, 
    -23.27892, -23.13189, -22.98453, -22.83684, -22.68882, -22.54047, 
    -22.39179, -22.24278, -22.09344, -21.94377, -21.79376, -21.64342, 
    -21.49276, -21.34175, -21.19041, -21.03874, -20.88674, -20.7344, 
    -20.58172, -20.42871, -20.27536, -20.12168, -19.96766, -19.8133, 
    -19.65861, -19.50358, -19.34822, -19.19251, -19.03647, -18.88009, 
    -18.72337, -18.56631, -18.40892, -18.25119, -18.09312, -17.93471, 
    -17.77596, -17.61687, -17.45744, -17.29768, -17.13757, -16.97713, 
    -16.81634, -16.65522, -16.49376, -16.33196, -16.16982, -16.00734, 
    -15.84452, -15.68137, -15.51787, -15.35404, -15.18986, -15.02535, 
    -14.86051, -14.69532, -14.5298, -14.36393, -14.19773, -14.0312, 
    -13.86433, -13.69712, -13.52957, -13.36169, -13.19348, -13.02493, 
    -12.85604, -12.68682, -12.51727, -12.34738, -12.17716, -12.00661, 
    -11.83572, -11.66451, -11.49296, -11.32109, -11.14888, -10.97635, 
    -10.80348, -10.63029, -10.45677, -10.28292, -10.10875, -9.934257, 
    -9.759436, -9.584291, -9.408824, -9.233035, -9.056924, -8.880493, 
    -8.703743, -8.526673, -8.349287, -8.171583, -7.993564, -7.815229, 
    -7.636581, -7.457621, -7.278347, -7.098764, -6.918871, -6.738669, 
    -6.55816, -6.377345, -6.196224, -6.0148, -5.833072, -5.651044, -5.468715, 
    -5.286088, -5.103162, -4.91994, -4.736424, -4.552614, -4.368512, 
    -4.184119, -3.999437, -3.814467, -3.629211, -3.44367, -3.257846, 
    -3.07174, -2.885354, -2.69869, -2.511748, -2.324532, -2.137042, -1.94928, 
    -1.761248, -1.572948, -1.384381, -1.19555, -1.006455, -0.8170998, 
    -0.627485, -0.4376127, -0.247485, -0.05710382, 0.133529, 0.3244114, 
    0.5155413, 0.7069169, 0.898536, 1.090397, 1.282496, 1.474834, 1.667406, 
    1.860211, 2.053247, 2.246512, 2.440003, 2.633718, 2.827655, 3.021812, 
    3.216186, 3.410775, 3.605576, 3.800588, 3.995808, 4.191233, 4.386861, 
    4.582689, 4.778716, 4.974938, 5.171353, 5.367959, 5.564754, 5.761733, 
    5.958895, 6.156237, 6.353757, 6.551453, 6.74932, 6.947357, 7.145561, 
    7.343929, 7.542459, 7.741147, 7.939992, 8.138989, 8.338138, 8.537434, 
    8.736874, 8.936457, 9.136178, 9.336036, 9.536027, 9.736148, 9.936398, 
    10.13677, 10.33727, 10.53788, 10.73861, 10.93945, 11.1404, 11.34146, 
    11.54263, 11.74389, 11.94525, 12.14671, 12.34825, 12.54989, 12.75161, 
    12.95341, 13.15529, 13.35725, 13.55928, 13.76138, 13.96355, 14.16578, 
    14.36808, 14.57043, 14.77283, 14.97528, 15.17778, 15.38033, 15.58292, 
    15.78555, 15.98821, 16.1909, 16.39362, 16.59637, 16.79914, 17.00193, 
    17.20473, 17.40755, 17.61037, 17.81321, 18.01604, 18.21888, 18.42171, 
    18.62453, 18.82735, 19.03015, 19.23294, 19.4357, 19.63845, 19.84116, 
    20.04385, 20.24651, 20.44913, 20.65171, 20.85425, 21.05675, 21.25919, 
    21.46159, 21.66393, 21.86621, 22.06843, 22.27059, 22.47268, 22.6747, 
    22.87665, 23.07852, 23.28031, 23.48201, 23.68364, 23.88517, 24.08661, 
    24.28795, 24.4892, 24.69035, 24.89139, 25.09233, 25.29315, 25.49386, 
    25.69446, 25.89493, 26.09529, 26.29552, 26.49562, 26.69559, 26.89542, 
    27.09512, 27.29468, 27.4941, 27.69337, 27.8925, 28.09147, 28.29029, 
    28.48896, 28.68746, 28.8858, 29.08398, 29.28199, 29.47983, 29.6775, 
    29.87499, 30.07231, 30.26944, 30.46639, 30.66315, 30.85973, 31.05611, 
    31.25231, 31.4483, 31.6441, 31.83969, 32.03509, 32.23027, 32.42525, 
    32.62002, 32.81458, 33.00891, 33.20304, 33.39694, 33.59062, 33.78407, 
    33.9773, 34.1703, 34.36307, 34.55561, 34.74791, 34.93997, 35.13179, 
    35.32337, 35.51471, 35.7058, 35.89664, 36.08723, 36.27758, 36.46766, 
    36.6575, 36.84707, 37.03638, 37.22544, 37.41423, 37.60275, 37.79101, 
    37.979, 38.16672, 38.35416, 38.54134, 38.72824, 38.91486, 39.1012, 
    39.28726, 39.47304, 39.65854, 39.84375, 40.02867, 40.21331, 40.39765, 
    40.58171, 40.76547, 40.94894, 41.13212, 41.31499, 41.49758, 41.67986, 
    41.86184, 42.04352, 42.2249, 42.40597, 42.58673, 42.76719, 42.94735, 
    43.12719, 43.30673, 43.48595, 43.66486, 43.84346, 44.02174, 44.19971, 
    44.37737, 44.5547, 44.73172, 44.90842, 45.0848, 45.26086, 45.4366, 
    45.61202, 45.78711, 45.96188, 46.13633, 46.31045, 46.48424, 46.65771, 
    46.83085, 47.00366, 47.17614, 47.3483, 47.52012, 47.69162, 47.86278, 
    48.03361, 48.20411, 48.37428, 48.54411, 48.71361, 48.88278, 49.05161, 
    49.22011, 49.38827, 49.5561, 49.72359, 49.89075, 50.05756, 50.22405, 
    50.39019,
  -28.45119, -28.31551, -28.17952, -28.04322, -27.90661, -27.7697, -27.63247, 
    -27.49493, -27.35707, -27.21891, -27.08043, -26.94164, -26.80253, 
    -26.66311, -26.52337, -26.38331, -26.24293, -26.10224, -25.96123, 
    -25.8199, -25.67825, -25.53627, -25.39398, -25.25136, -25.10842, 
    -24.96516, -24.82158, -24.67767, -24.53343, -24.38887, -24.24398, 
    -24.09877, -23.95323, -23.80736, -23.66116, -23.51463, -23.36778, 
    -23.22059, -23.07308, -22.92523, -22.77705, -22.62854, -22.4797, 
    -22.33052, -22.18102, -22.03117, -21.881, -21.73049, -21.57964, 
    -21.42846, -21.27695, -21.1251, -20.97291, -20.82038, -20.66752, 
    -20.51432, -20.36078, -20.20691, -20.0527, -19.89815, -19.74326, 
    -19.58803, -19.43246, -19.27655, -19.1203, -18.96371, -18.80679, 
    -18.64952, -18.49191, -18.33396, -18.17567, -18.01704, -17.85807, 
    -17.69876, -17.5391, -17.37911, -17.21877, -17.0581, -16.89708, 
    -16.73572, -16.57402, -16.41198, -16.24959, -16.08687, -15.9238, 
    -15.7604, -15.59665, -15.43256, -15.26813, -15.10336, -14.93825, 
    -14.7728, -14.60701, -14.44088, -14.27441, -14.1076, -13.94046, 
    -13.77297, -13.60515, -13.43698, -13.26848, -13.09965, -12.93047, 
    -12.76096, -12.59111, -12.42093, -12.25041, -12.07956, -11.90837, 
    -11.73685, -11.565, -11.39281, -11.22029, -11.04745, -10.87426, 
    -10.70075, -10.52691, -10.35274, -10.17825, -10.00342, -9.828268, 
    -9.65279, -9.476987, -9.300859, -9.124408, -8.947634, -8.770537, 
    -8.593121, -8.415383, -8.237328, -8.058953, -7.880261, -7.701253, 
    -7.52193, -7.342293, -7.162342, -6.98208, -6.801506, -6.620623, 
    -6.439431, -6.257931, -6.076126, -5.894015, -5.7116, -5.528883, 
    -5.345864, -5.162546, -4.978929, -4.795015, -4.610805, -4.4263, 
    -4.241502, -4.056413, -3.871034, -3.685366, -3.499411, -3.31317, 
    -3.126646, -2.939839, -2.752751, -2.565384, -2.37774, -2.18982, 
    -2.001626, -1.813159, -1.624422, -1.435416, -1.246144, -1.056606, 
    -0.8668045, -0.6767418, -0.4864196, -0.2958398, -0.1050043, 0.08608489, 
    0.2774258, 0.4690164, 0.6608547, 0.8529387, 1.045266, 1.237835, 1.430643, 
    1.623688, 1.816969, 2.010482, 2.204226, 2.398198, 2.592396, 2.786818, 
    2.981461, 3.176324, 3.371403, 3.566697, 3.762203, 3.957919, 4.153841, 
    4.349969, 4.546299, 4.742829, 4.939557, 5.136478, 5.333593, 5.530897, 
    5.728388, 5.926064, 6.123921, 6.321958, 6.520171, 6.718558, 6.917116, 
    7.115843, 7.314735, 7.513791, 7.713006, 7.912379, 8.111907, 8.311586, 
    8.511415, 8.71139, 8.911507, 9.111765, 9.31216, 9.512691, 9.713352, 
    9.914143, 10.11506, 10.3161, 10.51726, 10.71853, 10.91992, 11.12142, 
    11.32303, 11.52474, 11.72655, 11.92847, 12.13048, 12.33258, 12.53477, 
    12.73704, 12.9394, 13.14184, 13.34435, 13.54694, 13.7496, 13.95233, 
    14.15512, 14.35797, 14.56088, 14.76385, 14.96686, 15.16993, 15.37304, 
    15.57619, 15.77938, 15.9826, 16.18586, 16.38915, 16.59246, 16.79579, 
    16.99915, 17.20251, 17.4059, 17.60929, 17.81269, 18.01609, 18.21949, 
    18.42288, 18.62627, 18.82965, 19.03302, 19.23637, 19.4397, 19.64301, 
    19.84629, 20.04955, 20.25277, 20.45595, 20.65909, 20.8622, 21.06525, 
    21.26826, 21.47122, 21.67412, 21.87696, 22.07974, 22.28246, 22.48511, 
    22.68769, 22.89019, 23.09262, 23.29496, 23.49722, 23.6994, 23.90149, 
    24.10348, 24.30538, 24.50717, 24.70887, 24.91046, 25.11194, 25.31331, 
    25.51457, 25.71571, 25.91673, 26.11763, 26.3184, 26.51904, 26.71955, 
    26.91992, 27.12016, 27.32025, 27.5202, 27.72001, 27.91966, 28.11917, 
    28.31852, 28.51771, 28.71674, 28.9156, 29.1143, 29.31284, 29.51119, 
    29.70938, 29.90739, 30.10522, 30.30286, 30.50033, 30.6976, 30.89468, 
    31.09158, 31.28827, 31.48477, 31.68107, 31.87716, 32.07306, 32.26874, 
    32.46421, 32.65947, 32.85452, 33.04934, 33.24395, 33.43834, 33.6325, 
    33.82644, 34.02015, 34.21362, 34.40686, 34.59987, 34.79264, 34.98517, 
    35.17746, 35.36951, 35.56131, 35.75286, 35.94416, 36.13521, 36.326, 
    36.51654, 36.70683, 36.89685, 37.08661, 37.2761, 37.46533, 37.6543, 
    37.84299, 38.03141, 38.21956, 38.40744, 38.59504, 38.78236, 38.96941, 
    39.15617, 39.34265, 39.52884, 39.71476, 39.90038, 40.08571, 40.27075, 
    40.45551, 40.63997, 40.82413, 41.008, 41.19156, 41.37484, 41.5578, 
    41.74047, 41.92284, 42.1049, 42.28666, 42.46811, 42.64926, 42.83009, 
    43.01062, 43.19083, 43.37073, 43.55032, 43.72959, 43.90855, 44.08719, 
    44.26551, 44.44352, 44.62121, 44.79857, 44.97562, 45.15234, 45.32874, 
    45.50482, 45.68057, 45.856, 46.0311, 46.20587, 46.38032, 46.55443, 
    46.72822, 46.90168, 47.07481, 47.24761, 47.42007, 47.59221, 47.76401, 
    47.93547, 48.10661, 48.27741, 48.44788, 48.618, 48.7878, 48.95726, 
    49.12638, 49.29516, 49.46361, 49.63171, 49.79949, 49.96692, 50.13401, 
    50.30077, 50.46718,
  -28.54487, -28.40909, -28.273, -28.1366, -27.99989, -27.86287, -27.72554, 
    -27.58789, -27.44993, -27.31166, -27.17307, -27.03416, -26.89494, 
    -26.7554, -26.61555, -26.47537, -26.33488, -26.19406, -26.05293, 
    -25.91147, -25.7697, -25.6276, -25.48517, -25.34243, -25.19936, 
    -25.05596, -24.91224, -24.76819, -24.62382, -24.47912, -24.33409, 
    -24.18873, -24.04304, -23.89703, -23.75068, -23.604, -23.457, -23.30966, 
    -23.16198, -23.01398, -22.86564, -22.71697, -22.56796, -22.41862, 
    -22.26895, -22.11894, -21.96859, -21.81791, -21.66689, -21.51554, 
    -21.36384, -21.21181, -21.05944, -20.90673, -20.75368, -20.6003, 
    -20.44657, -20.2925, -20.1381, -19.98335, -19.82826, -19.67283, 
    -19.51707, -19.36095, -19.2045, -19.0477, -18.89057, -18.73309, 
    -18.57527, -18.4171, -18.25859, -18.09974, -17.94055, -17.78101, 
    -17.62113, -17.46091, -17.30034, -17.13943, -16.97818, -16.81658, 
    -16.65464, -16.49236, -16.32973, -16.16676, -16.00344, -15.83979, 
    -15.67579, -15.51145, -15.34676, -15.18173, -15.01636, -14.85064, 
    -14.68459, -14.51819, -14.35145, -14.18437, -14.01695, -13.84918, 
    -13.68108, -13.51263, -13.34385, -13.17472, -13.00526, -12.83546, 
    -12.66532, -12.49484, -12.32402, -12.15287, -11.98138, -11.80955, 
    -11.63739, -11.46489, -11.29206, -11.1189, -10.9454, -10.77157, -10.5974, 
    -10.42291, -10.24809, -10.07293, -9.897447, -9.721634, -9.545494, 
    -9.369027, -9.192234, -9.015116, -8.837673, -8.659907, -8.481819, 
    -8.30341, -8.124679, -7.945629, -7.76626, -7.586573, -7.40657, -7.226251, 
    -7.045618, -6.864672, -6.683413, -6.501843, -6.319963, -6.137775, 
    -5.955279, -5.772477, -5.58937, -5.40596, -5.222247, -5.038232, 
    -4.853919, -4.669307, -4.484398, -4.299194, -4.113696, -3.927906, 
    -3.741824, -3.555454, -3.368795, -3.18185, -2.99462, -2.807107, 
    -2.619313, -2.431239, -2.242887, -2.054259, -1.865356, -1.676181, 
    -1.486734, -1.297018, -1.107035, -0.9167857, -0.7262732, -0.5354989, 
    -0.3444649, -0.153173, 0.0383747, 0.2301763, 0.4222297, 0.6145329, 
    0.8070839, 0.9998804, 1.192921, 1.386202, 1.579723, 1.77348, 1.967473, 
    2.161698, 2.356153, 2.550837, 2.745746, 2.940879, 3.136232, 3.331805, 
    3.527594, 3.723597, 3.919811, 4.116234, 4.312864, 4.509699, 4.706735, 
    4.903969, 5.101401, 5.299026, 5.496843, 5.694849, 5.89304, 6.091415, 
    6.289971, 6.488706, 6.687615, 6.886698, 7.08595, 7.285369, 7.484954, 
    7.6847, 7.884604, 8.084664, 8.284878, 8.485242, 8.685754, 8.88641, 
    9.087208, 9.288144, 9.489216, 9.690421, 9.891756, 10.09322, 10.2948, 
    10.49651, 10.69833, 10.90027, 11.10232, 11.30448, 11.50675, 11.70912, 
    11.91158, 12.11415, 12.3168, 12.51955, 12.72239, 12.9253, 13.1283, 
    13.33138, 13.53453, 13.73775, 13.94104, 14.14439, 14.34781, 14.55128, 
    14.75481, 14.9584, 15.16202, 15.3657, 15.56942, 15.77317, 15.97697, 
    16.18079, 16.38464, 16.58852, 16.79243, 16.99635, 17.20028, 17.40424, 
    17.6082, 17.81216, 18.01613, 18.2201, 18.42407, 18.62803, 18.83197, 
    19.03591, 19.23983, 19.44373, 19.6476, 19.85145, 20.05527, 20.25906, 
    20.46281, 20.66652, 20.87019, 21.07381, 21.27739, 21.48091, 21.68437, 
    21.88778, 22.09112, 22.2944, 22.49761, 22.70075, 22.90381, 23.1068, 
    23.3097, 23.51253, 23.71526, 23.9179, 24.12045, 24.3229, 24.52525, 
    24.7275, 24.92964, 25.13168, 25.3336, 25.5354, 25.73709, 25.93866, 
    26.1401, 26.34142, 26.5426, 26.74365, 26.94456, 27.14534, 27.34597, 
    27.54646, 27.7468, 27.94699, 28.14703, 28.34691, 28.54663, 28.74619, 
    28.94558, 29.14481, 29.34386, 29.54274, 29.74145, 29.93998, 30.13832, 
    30.33648, 30.53446, 30.73225, 30.92984, 31.12724, 31.32445, 31.52145, 
    31.71825, 31.91485, 32.11124, 32.30742, 32.50339, 32.69915, 32.89468, 
    33.09, 33.2851, 33.47997, 33.67462, 33.86904, 34.06323, 34.25718, 
    34.4509, 34.64439, 34.83763, 35.03063, 35.22339, 35.4159, 35.60817, 
    35.80018, 35.99194, 36.18345, 36.3747, 36.56569, 36.75643, 36.9469, 
    37.1371, 37.32705, 37.51672, 37.70612, 37.89526, 38.08411, 38.2727, 
    38.46101, 38.64904, 38.83679, 39.02426, 39.21144, 39.39834, 39.58495, 
    39.77128, 39.95731, 40.14306, 40.32851, 40.51367, 40.69853, 40.88309, 
    41.06736, 41.25133, 41.43499, 41.61835, 41.80141, 41.98417, 42.16661, 
    42.34875, 42.53059, 42.7121, 42.89331, 43.07421, 43.2548, 43.43507, 
    43.61502, 43.79465, 43.97397, 44.15297, 44.33165, 44.51001, 44.68805, 
    44.86576, 45.04316, 45.22022, 45.39696, 45.57338, 45.74947, 45.92523, 
    46.10066, 46.27576, 46.45053, 46.62498, 46.79909, 46.97287, 47.14631, 
    47.31942, 47.4922, 47.66465, 47.83675, 48.00853, 48.17997, 48.35107, 
    48.52183, 48.69225, 48.86234, 49.03209, 49.2015, 49.37057, 49.5393, 
    49.70769, 49.87574, 50.04345, 50.21082, 50.37785, 50.54453,
  -28.63888, -28.503, -28.36681, -28.23032, -28.09351, -27.95638, -27.81894, 
    -27.68119, -27.54313, -27.40475, -27.26605, -27.12703, -26.9877, 
    -26.84804, -26.70807, -26.56778, -26.42717, -26.28623, -26.14498, 
    -26.0034, -25.86149, -25.71927, -25.57672, -25.43384, -25.29064, 
    -25.14711, -25.00325, -24.85907, -24.71456, -24.56972, -24.42455, 
    -24.27905, -24.13321, -23.98705, -23.84056, -23.69373, -23.54657, 
    -23.39908, -23.25125, -23.10309, -22.95459, -22.80576, -22.65659, 
    -22.50709, -22.35724, -22.20707, -22.05655, -21.90569, -21.7545, 
    -21.60297, -21.4511, -21.29889, -21.14634, -20.99344, -20.84021, 
    -20.68664, -20.53272, -20.37846, -20.22386, -20.06892, -19.91364, 
    -19.75801, -19.60204, -19.44572, -19.28906, -19.13206, -18.97471, 
    -18.81702, -18.65899, -18.50061, -18.34188, -18.18281, -18.02339, 
    -17.86363, -17.70353, -17.54308, -17.38228, -17.22113, -17.05965, 
    -16.89781, -16.73563, -16.57311, -16.41023, -16.24702, -16.08346, 
    -15.91955, -15.75529, -15.5907, -15.42575, -15.26046, -15.09483, 
    -14.92885, -14.76253, -14.59586, -14.42885, -14.2615, -14.0938, 
    -13.92576, -13.75737, -13.58865, -13.41958, -13.25016, -13.08041, 
    -12.91032, -12.73988, -12.56911, -12.39799, -12.22653, -12.05474, 
    -11.88261, -11.71014, -11.53733, -11.36419, -11.1907, -11.01689, 
    -10.84274, -10.66825, -10.49343, -10.31828, -10.14279, -9.966974, 
    -9.790826, -9.614348, -9.437541, -9.260406, -9.082943, -8.905153, 
    -8.727037, -8.548596, -8.369832, -8.190744, -8.011334, -7.831604, 
    -7.651552, -7.471182, -7.290494, -7.109489, -6.928168, -6.746533, 
    -6.564584, -6.382323, -6.19975, -6.016868, -5.833677, -5.650179, 
    -5.466375, -5.282266, -5.097854, -4.913139, -4.728124, -4.54281, 
    -4.357198, -4.171289, -3.985086, -3.79859, -3.611802, -3.424723, 
    -3.237356, -3.049702, -2.861762, -2.673539, -2.485034, -2.296248, 
    -2.107183, -1.917842, -1.728226, -1.538336, -1.348175, -1.157744, 
    -0.9670459, -0.7760816, -0.5848532, -0.3933629, -0.2016125, -0.009604137, 
    0.1826603, 0.3751787, 0.5679491, 0.7609693, 0.9542372, 1.147751, 
    1.341508, 1.535506, 1.729743, 1.924218, 2.118927, 2.313868, 2.509039, 
    2.704438, 2.900062, 3.09591, 3.291978, 3.488264, 3.684767, 3.881482, 
    4.078409, 4.275544, 4.472885, 4.670429, 4.868175, 5.066118, 5.264257, 
    5.46259, 5.661112, 5.859823, 6.058719, 6.257797, 6.457055, 6.65649, 
    6.8561, 7.055881, 7.25583, 7.455946, 7.656225, 7.856664, 8.057261, 
    8.258011, 8.458914, 8.659966, 8.861163, 9.062503, 9.263984, 9.465601, 
    9.667353, 9.869235, 10.07125, 10.27338, 10.47564, 10.67801, 10.88051, 
    11.08311, 11.28583, 11.48865, 11.69157, 11.8946, 12.09772, 12.30094, 
    12.50425, 12.70764, 12.91112, 13.11469, 13.31833, 13.52204, 13.72583, 
    13.92968, 14.1336, 14.33759, 14.54163, 14.74572, 14.94987, 15.15407, 
    15.35832, 15.5626, 15.76693, 15.97129, 16.17569, 16.38011, 16.58457, 
    16.78904, 16.99353, 17.19804, 17.40257, 17.6071, 17.81164, 18.01618, 
    18.22072, 18.42526, 18.62979, 18.83431, 19.03882, 19.24331, 19.44778, 
    19.65222, 19.85664, 20.06104, 20.26539, 20.46971, 20.67399, 20.87823, 
    21.08242, 21.28656, 21.49065, 21.69468, 21.89866, 22.10257, 22.30641, 
    22.51019, 22.71389, 22.91752, 23.12107, 23.32454, 23.52792, 23.73121, 
    23.93441, 24.13752, 24.34053, 24.54344, 24.74625, 24.94894, 25.15153, 
    25.35401, 25.55636, 25.7586, 25.96072, 26.16271, 26.36457, 26.5663, 
    26.7679, 26.96935, 27.17067, 27.37185, 27.57288, 27.77375, 27.97448, 
    28.17505, 28.37547, 28.57572, 28.77581, 28.97573, 29.17549, 29.37507, 
    29.57448, 29.77371, 29.97276, 30.17162, 30.3703, 30.5688, 30.7671, 
    30.96521, 31.16312, 31.36083, 31.55835, 31.75565, 31.95275, 32.14965, 
    32.34633, 32.5428, 32.73905, 32.93509, 33.1309, 33.32648, 33.52185, 
    33.71698, 33.91189, 34.10656, 34.301, 34.4952, 34.68916, 34.88288, 
    35.07635, 35.26958, 35.46256, 35.65529, 35.84777, 36.03999, 36.23196, 
    36.42367, 36.61512, 36.8063, 36.99723, 37.18789, 37.37827, 37.56839, 
    37.75824, 37.94781, 38.13711, 38.32613, 38.51487, 38.70333, 38.89151, 
    39.0794, 39.26701, 39.45433, 39.64137, 39.82811, 40.01456, 40.20072, 
    40.38658, 40.57214, 40.75741, 40.94238, 41.12704, 41.31141, 41.49547, 
    41.67923, 41.86267, 42.04582, 42.22865, 42.41117, 42.59339, 42.77528, 
    42.95687, 43.13814, 43.3191, 43.49974, 43.68005, 43.86005, 44.03973, 
    44.21909, 44.39813, 44.57684, 44.75523, 44.9333, 45.11104, 45.28845, 
    45.46553, 45.64229, 45.81871, 45.99481, 46.17057, 46.346, 46.52111, 
    46.69587, 46.8703, 47.0444, 47.21817, 47.3916, 47.56469, 47.73744, 
    47.90986, 48.08194, 48.25368, 48.42508, 48.59614, 48.76686, 48.93724, 
    49.10728, 49.27699, 49.44634, 49.61536, 49.78403, 49.95236, 50.12035, 
    50.28799, 50.4553, 50.62225,
  -28.73322, -28.59725, -28.46097, -28.32437, -28.18746, -28.05024, 
    -27.91269, -27.77484, -27.63667, -27.49818, -27.35937, -27.22024, 
    -27.0808, -26.94103, -26.80094, -26.66054, -26.5198, -26.37875, 
    -26.23737, -26.09567, -25.95364, -25.81129, -25.66861, -25.52561, 
    -25.38227, -25.23861, -25.09462, -24.9503, -24.80565, -24.66067, 
    -24.51536, -24.36972, -24.22374, -24.07743, -23.93079, -23.78381, 
    -23.6365, -23.48886, -23.34087, -23.19256, -23.0439, -22.89491, 
    -22.74558, -22.59591, -22.4459, -22.29556, -22.14487, -21.99384, 
    -21.84248, -21.69077, -21.53872, -21.38633, -21.2336, -21.08052, 
    -20.9271, -20.77334, -20.61924, -20.46479, -20.31, -20.15486, -19.99938, 
    -19.84355, -19.68738, -19.53086, -19.374, -19.21679, -19.05923, 
    -18.90133, -18.74308, -18.58448, -18.42554, -18.26625, -18.10661, 
    -17.94662, -17.78629, -17.62561, -17.46458, -17.30321, -17.14148, 
    -16.97941, -16.81699, -16.65422, -16.49111, -16.32765, -16.16384, 
    -15.99968, -15.83517, -15.67032, -15.50512, -15.33957, -15.17367, 
    -15.00743, -14.84084, -14.6739, -14.50662, -14.33899, -14.17102, 
    -14.0027, -13.83403, -13.66502, -13.49567, -13.32597, -13.15593, 
    -12.98554, -12.81481, -12.64374, -12.47232, -12.30056, -12.12846, 
    -11.95603, -11.78325, -11.61013, -11.43667, -11.26287, -11.08873, 
    -10.91426, -10.73945, -10.5643, -10.38882, -10.213, -10.03685, -9.86037, 
    -9.683554, -9.506406, -9.328926, -9.151117, -8.97298, -8.794513, 
    -8.615719, -8.436598, -8.257152, -8.077381, -7.897287, -7.716871, 
    -7.536132, -7.355074, -7.173696, -6.992, -6.809986, -6.627657, -6.445013, 
    -6.262055, -6.078785, -5.895205, -5.711314, -5.527114, -5.342608, 
    -5.157795, -4.972679, -4.787259, -4.601538, -4.415516, -4.229196, 
    -4.042578, -3.855665, -3.668458, -3.480958, -3.293167, -3.105086, 
    -2.916718, -2.728064, -2.539125, -2.349904, -2.160401, -1.97062, 
    -1.780561, -1.590227, -1.399618, -1.208738, -1.017588, -0.8261696, 
    -0.6344851, -0.4425364, -0.2503254, -0.05785418, 0.1348753, 0.3278609, 
    0.5211006, 0.7145923, 0.908334, 1.102323, 1.296558, 1.491037, 1.685756, 
    1.880714, 2.075909, 2.271339, 2.467, 2.662892, 2.85901, 3.055354, 
    3.25192, 3.448707, 3.645711, 3.84293, 4.040363, 4.238005, 4.435856, 
    4.633912, 4.83217, 5.030628, 5.229284, 5.428135, 5.627178, 5.82641, 
    6.025829, 6.225433, 6.425218, 6.625181, 6.82532, 7.025633, 7.226116, 
    7.426765, 7.627581, 7.828557, 8.029693, 8.230984, 8.432428, 8.634023, 
    8.835765, 9.037651, 9.239678, 9.441844, 9.644145, 9.846579, 10.04914, 
    10.25183, 10.45464, 10.65757, 10.86062, 11.06379, 11.26706, 11.47044, 
    11.67393, 11.87751, 12.0812, 12.28498, 12.48885, 12.69281, 12.89686, 
    13.10098, 13.30519, 13.50947, 13.71383, 13.91825, 14.12274, 14.3273, 
    14.53191, 14.73658, 14.9413, 15.14607, 15.35089, 15.55575, 15.76065, 
    15.96559, 16.17056, 16.37556, 16.58058, 16.78563, 16.9907, 17.19579, 
    17.40088, 17.60599, 17.81111, 18.01622, 18.22134, 18.42645, 18.63156, 
    18.83666, 19.04174, 19.24681, 19.45185, 19.65687, 19.86187, 20.06683, 
    20.27176, 20.47666, 20.68151, 20.88632, 21.09109, 21.2958, 21.50046, 
    21.70506, 21.90961, 22.11409, 22.3185, 22.52284, 22.72712, 22.93131, 
    23.13543, 23.33946, 23.54341, 23.74726, 23.95103, 24.1547, 24.35827, 
    24.56174, 24.7651, 24.96836, 25.1715, 25.37453, 25.57745, 25.78024, 
    25.98291, 26.18545, 26.38787, 26.59015, 26.79229, 26.99429, 27.19616, 
    27.39788, 27.59945, 27.80087, 28.00213, 28.20325, 28.4042, 28.60498, 
    28.80561, 29.00607, 29.20635, 29.40646, 29.6064, 29.80615, 30.00573, 
    30.20512, 30.40432, 30.60333, 30.80215, 31.00078, 31.19921, 31.39743, 
    31.59546, 31.79327, 31.99088, 32.18828, 32.38547, 32.58244, 32.77919, 
    32.97572, 33.17203, 33.36811, 33.56396, 33.75959, 33.95498, 34.15014, 
    34.34506, 34.53974, 34.73418, 34.92838, 35.12233, 35.31603, 35.50948, 
    35.70268, 35.89563, 36.08832, 36.28075, 36.47292, 36.66483, 36.85647, 
    37.04784, 37.23895, 37.42979, 37.62035, 37.81064, 38.00066, 38.1904, 
    38.37985, 38.56903, 38.75792, 38.94653, 39.13486, 39.32289, 39.51064, 
    39.69809, 39.88525, 40.07212, 40.25869, 40.44496, 40.63094, 40.81661, 
    41.00198, 41.18705, 41.37181, 41.55627, 41.74042, 41.92426, 42.1078, 
    42.29102, 42.47393, 42.65652, 42.8388, 43.02076, 43.20241, 43.38374, 
    43.56474, 43.74543, 43.9258, 44.10584, 44.28556, 44.46495, 44.64402, 
    44.82277, 45.00118, 45.17926, 45.35702, 45.53445, 45.71154, 45.88831, 
    46.06474, 46.24084, 46.4166, 46.59203, 46.76712, 46.94188, 47.1163, 
    47.29038, 47.46413, 47.63753, 47.8106, 47.98333, 48.15571, 48.32775, 
    48.49946, 48.67082, 48.84184, 49.01252, 49.18285, 49.35284, 49.52248, 
    49.69178, 49.86074, 50.02935, 50.19761, 50.36553, 50.53311, 50.70033,
  -28.82791, -28.69184, -28.55546, -28.41877, -28.28176, -28.14443, 
    -28.00679, -27.86883, -27.73055, -27.59195, -27.45304, -27.3138, 
    -27.17424, -27.03437, -26.89417, -26.75364, -26.61279, -26.47162, 
    -26.33012, -26.1883, -26.04615, -25.90367, -25.76086, -25.61773, 
    -25.47427, -25.33047, -25.18635, -25.04189, -24.89711, -24.75199, 
    -24.60654, -24.46075, -24.31463, -24.16818, -24.02139, -23.87426, 
    -23.7268, -23.579, -23.43086, -23.28239, -23.13358, -22.98442, -22.83493, 
    -22.6851, -22.53493, -22.38441, -22.23356, -22.08236, -21.93082, 
    -21.77894, -21.62671, -21.47414, -21.32123, -21.16797, -21.01437, 
    -20.86042, -20.70613, -20.55149, -20.3965, -20.24117, -20.08549, 
    -19.92946, -19.77309, -19.61637, -19.4593, -19.30188, -19.14412, -18.986, 
    -18.82754, -18.66873, -18.50957, -18.35006, -18.1902, -18.02999, 
    -17.86943, -17.70852, -17.54726, -17.38565, -17.22369, -17.06138, 
    -16.89873, -16.73572, -16.57236, -16.40865, -16.24459, -16.08018, 
    -15.91542, -15.75031, -15.58485, -15.41904, -15.25288, -15.08638, 
    -14.91952, -14.75232, -14.58476, -14.41686, -14.24861, -14.08001, 
    -13.91106, -13.74177, -13.57213, -13.40214, -13.23181, -13.06113, 
    -12.8901, -12.71873, -12.54702, -12.37496, -12.20255, -12.0298, 
    -11.85671, -11.68328, -11.50951, -11.33539, -11.16094, -10.98614, 
    -10.81101, -10.63553, -10.45972, -10.28357, -10.10709, -9.930268, 
    -9.753112, -9.575622, -9.397799, -9.219643, -9.041155, -8.862336, 
    -8.683188, -8.503711, -8.323905, -8.143773, -7.963315, -7.782531, 
    -7.601424, -7.419993, -7.238241, -7.056168, -6.873775, -6.691064, 
    -6.508037, -6.324692, -6.141033, -5.957061, -5.772776, -5.58818, 
    -5.403275, -5.218061, -5.03254, -4.846714, -4.660584, -4.474152, 
    -4.287417, -4.100384, -3.913052, -3.725424, -3.537501, -3.349284, 
    -3.160776, -2.971977, -2.78289, -2.593517, -2.403858, -2.213916, 
    -2.023692, -1.833189, -1.642407, -1.45135, -1.260018, -1.068414, 
    -0.8765399, -0.6843972, -0.491988, -0.2993142, -0.106378, 0.08681865, 
    0.2802737, 0.473985, 0.6679505, 0.8621681, 1.056635, 1.251351, 1.446311, 
    1.641515, 1.83696, 2.032644, 2.228564, 2.424718, 2.621104, 2.817719, 
    3.014562, 3.211629, 3.408918, 3.606427, 3.804153, 4.002094, 4.200247, 
    4.398609, 4.597179, 4.795953, 4.994929, 5.194105, 5.393476, 5.593042, 
    5.792799, 5.992745, 6.192877, 6.393191, 6.593686, 6.794358, 6.995205, 
    7.196224, 7.397411, 7.598765, 7.800282, 8.00196, 8.203794, 8.405784, 
    8.607924, 8.810214, 9.01265, 9.215227, 9.417945, 9.620798, 9.823786, 
    10.0269, 10.23015, 10.43352, 10.63701, 10.84062, 11.04434, 11.24818, 
    11.45212, 11.65617, 11.86032, 12.06457, 12.26892, 12.47336, 12.67789, 
    12.8825, 13.0872, 13.29198, 13.49683, 13.70176, 13.90676, 14.11182, 
    14.31695, 14.52213, 14.72738, 14.93268, 15.13802, 15.34342, 15.54885, 
    15.75433, 15.95985, 16.16539, 16.37097, 16.57658, 16.7822, 16.98785, 
    17.19351, 17.39919, 17.60488, 17.81057, 18.01627, 18.22197, 18.42766, 
    18.63334, 18.83902, 19.04468, 19.25033, 19.45595, 19.66155, 19.86712, 
    20.07266, 20.27817, 20.48364, 20.68908, 20.89446, 21.0998, 21.30509, 
    21.51033, 21.7155, 21.92062, 22.12568, 22.33066, 22.53558, 22.74042, 
    22.94518, 23.14987, 23.35447, 23.55899, 23.76341, 23.96774, 24.17198, 
    24.37611, 24.58015, 24.78407, 24.98789, 25.1916, 25.39519, 25.59866, 
    25.80201, 26.00524, 26.20833, 26.4113, 26.61413, 26.81683, 27.01938, 
    27.22179, 27.42406, 27.62618, 27.82814, 28.02995, 28.23161, 28.4331, 
    28.63442, 28.83559, 29.03658, 29.2374, 29.43804, 29.63851, 29.83879, 
    30.03889, 30.23881, 30.43854, 30.63807, 30.83741, 31.03656, 31.2355, 
    31.43424, 31.63278, 31.83111, 32.02923, 32.22714, 32.42483, 32.6223, 
    32.81956, 33.01659, 33.2134, 33.40998, 33.60633, 33.80244, 33.99833, 
    34.19397, 34.38938, 34.58455, 34.77946, 34.97414, 35.16857, 35.36275, 
    35.55667, 35.75034, 35.94376, 36.13691, 36.32981, 36.52244, 36.71481, 
    36.90691, 37.09874, 37.2903, 37.48159, 37.6726, 37.86334, 38.0538, 
    38.24398, 38.43388, 38.62349, 38.81282, 39.00186, 39.19061, 39.37908, 
    39.56725, 39.75512, 39.9427, 40.12999, 40.31697, 40.50366, 40.69005, 
    40.87613, 41.06191, 41.24738, 41.43254, 41.6174, 41.80195, 41.98618, 
    42.1701, 42.35371, 42.53701, 42.71999, 42.90265, 43.08499, 43.26701, 
    43.44872, 43.63009, 43.81115, 43.99188, 44.17229, 44.35237, 44.53212, 
    44.71155, 44.89064, 45.06941, 45.24784, 45.42595, 45.60372, 45.78116, 
    45.95826, 46.13503, 46.31146, 46.48756, 46.66331, 46.83873, 47.01381, 
    47.18856, 47.36296, 47.53702, 47.71074, 47.88412, 48.05715, 48.22985, 
    48.40219, 48.5742, 48.74586, 48.91718, 49.08815, 49.25877, 49.42905, 
    49.59899, 49.76857, 49.93781, 50.1067, 50.27525, 50.44344, 50.61129, 
    50.77879,
  -28.92294, -28.78677, -28.6503, -28.5135, -28.3764, -28.23897, -28.10123, 
    -27.96316, -27.82478, -27.68608, -27.54706, -27.40771, -27.26804, 
    -27.12805, -26.98774, -26.8471, -26.70613, -26.56484, -26.42322, 
    -26.28128, -26.139, -25.9964, -25.85347, -25.71021, -25.56661, -25.42269, 
    -25.27843, -25.13384, -24.98892, -24.84366, -24.69807, -24.55215, 
    -24.40588, -24.25928, -24.11234, -23.96507, -23.81746, -23.66951, 
    -23.52122, -23.37259, -23.22362, -23.0743, -22.92465, -22.77465, 
    -22.62432, -22.47364, -22.32261, -22.17124, -22.01953, -21.86747, 
    -21.71507, -21.56232, -21.40923, -21.25579, -21.102, -20.94787, 
    -20.79339, -20.63856, -20.48338, -20.32785, -20.17198, -20.01575, 
    -19.85918, -19.70225, -19.54498, -19.38736, -19.22938, -19.07106, 
    -18.91238, -18.75335, -18.59397, -18.43424, -18.27416, -18.11373, 
    -17.95294, -17.79181, -17.63032, -17.46847, -17.30628, -17.14373, 
    -16.98083, -16.81758, -16.65398, -16.49002, -16.32572, -16.16105, 
    -15.99604, -15.83068, -15.66496, -15.49889, -15.33247, -15.1657, 
    -14.99858, -14.8311, -14.66328, -14.4951, -14.32657, -14.15769, 
    -13.98847, -13.81889, -13.64896, -13.47868, -13.30806, -13.13708, 
    -12.96576, -12.79409, -12.62208, -12.44971, -12.27701, -12.10395, 
    -11.93055, -11.7568, -11.58272, -11.40828, -11.23351, -11.05839, 
    -10.88293, -10.70713, -10.53098, -10.3545, -10.17768, -10.00052, 
    -9.823027, -9.645194, -9.467026, -9.288522, -9.109683, -8.930512, 
    -8.751008, -8.571173, -8.391007, -8.210512, -8.029688, -7.848536, 
    -7.667059, -7.485255, -7.303128, -7.120677, -6.937904, -6.75481, 
    -6.571396, -6.387664, -6.203615, -6.019249, -5.834569, -5.649575, 
    -5.46427, -5.278653, -5.092727, -4.906493, -4.719953, -4.533107, 
    -4.345958, -4.158507, -3.970755, -3.782704, -3.594356, -3.405712, 
    -3.216774, -3.027543, -2.838022, -2.648211, -2.458113, -2.267729, 
    -2.077061, -1.886111, -1.694881, -1.503372, -1.311587, -1.119528, 
    -0.9271954, -0.7345922, -0.5417203, -0.3485817, -0.1551783, 0.0384878, 
    0.2324145, 0.4265997, 0.6210412, 0.8157371, 1.010685, 1.205883, 1.401328, 
    1.597019, 1.792953, 1.989128, 2.185541, 2.38219, 2.579073, 2.776188, 
    2.973532, 3.171102, 3.368897, 3.566913, 3.765148, 3.9636, 4.162266, 
    4.361144, 4.56023, 4.759523, 4.959019, 5.158717, 5.358613, 5.558704, 
    5.758989, 5.959464, 6.160126, 6.360973, 6.562003, 6.76321, 6.964595, 
    7.166152, 7.367881, 7.569777, 7.771838, 7.97406, 8.176441, 8.378979, 
    8.58167, 8.78451, 8.987497, 9.190628, 9.3939, 9.59731, 9.800855, 
    10.00453, 10.20834, 10.41227, 10.61632, 10.82049, 11.02478, 11.22918, 
    11.43369, 11.63831, 11.84303, 12.04784, 12.25276, 12.45777, 12.66287, 
    12.86806, 13.07333, 13.27868, 13.48411, 13.68962, 13.89519, 14.10083, 
    14.30653, 14.5123, 14.71812, 14.924, 15.12992, 15.3359, 15.54192, 
    15.74797, 15.95407, 16.1602, 16.36636, 16.57254, 16.77875, 16.98498, 
    17.19123, 17.39749, 17.60376, 17.81004, 18.01632, 18.22259, 18.42887, 
    18.63514, 18.8414, 19.04764, 19.25387, 19.46007, 19.66626, 19.87241, 
    20.07853, 20.28462, 20.49067, 20.69669, 20.90265, 21.10857, 21.31444, 
    21.52025, 21.72601, 21.9317, 22.13733, 22.3429, 22.54839, 22.75381, 
    22.95914, 23.1644, 23.36958, 23.57466, 23.77966, 23.98456, 24.18937, 
    24.39407, 24.59867, 24.80316, 25.00755, 25.21181, 25.41597, 25.62, 
    25.82391, 26.0277, 26.23135, 26.43488, 26.63826, 26.84151, 27.04462, 
    27.24759, 27.4504, 27.65307, 27.85558, 28.05794, 28.26014, 28.46217, 
    28.66404, 28.86574, 29.06727, 29.26863, 29.46981, 29.67081, 29.87163, 
    30.07226, 30.27271, 30.47296, 30.67302, 30.87288, 31.07255, 31.27202, 
    31.47128, 31.67033, 31.86917, 32.06781, 32.26622, 32.46442, 32.66241, 
    32.86016, 33.0577, 33.25501, 33.45209, 33.64893, 33.84554, 34.04192, 
    34.23806, 34.43395, 34.6296, 34.82501, 35.02017, 35.21508, 35.40973, 
    35.60413, 35.79828, 35.99216, 36.18579, 36.37915, 36.57225, 36.76508, 
    36.95764, 37.14993, 37.34194, 37.53368, 37.72515, 37.91634, 38.10724, 
    38.29786, 38.4882, 38.67825, 38.86802, 39.0575, 39.24668, 39.43557, 
    39.62417, 39.81247, 40.00047, 40.18818, 40.37558, 40.56268, 40.74948, 
    40.93597, 41.12216, 41.30804, 41.4936, 41.67886, 41.8638, 42.04844, 
    42.23275, 42.41675, 42.60043, 42.78379, 42.96684, 43.14956, 43.33196, 
    43.51403, 43.69579, 43.87721, 44.05832, 44.23909, 44.41953, 44.59964, 
    44.77943, 44.95888, 45.138, 45.31678, 45.49523, 45.67335, 45.85113, 
    46.02857, 46.20567, 46.38244, 46.55887, 46.73496, 46.91071, 47.08611, 
    47.26118, 47.4359, 47.61028, 47.78431, 47.958, 48.13135, 48.30435, 
    48.477, 48.64931, 48.82127, 48.99289, 49.16415, 49.33507, 49.50564, 
    49.67587, 49.84573, 50.01526, 50.18443, 50.35325, 50.52172, 50.68985, 
    50.85762,
  -29.0183, -28.88205, -28.74548, -28.60859, -28.47138, -28.33386, -28.19601, 
    -28.05785, -27.91936, -27.78055, -27.64142, -27.50197, -27.36219, 
    -27.22209, -27.08166, -26.94091, -26.79983, -26.65842, -26.51668, 
    -26.37461, -26.23222, -26.08949, -25.94643, -25.80305, -25.65932, 
    -25.51527, -25.37088, -25.22616, -25.0811, -24.9357, -24.78997, -24.6439, 
    -24.4975, -24.35075, -24.20367, -24.05625, -23.90849, -23.76038, 
    -23.61194, -23.46315, -23.31402, -23.16455, -23.01474, -22.86458, 
    -22.71408, -22.56323, -22.41204, -22.2605, -22.10862, -21.95638, 
    -21.80381, -21.65088, -21.49761, -21.34398, -21.19001, -21.03569, 
    -20.88102, -20.726, -20.57063, -20.41491, -20.25884, -20.10242, 
    -19.94564, -19.78852, -19.63104, -19.47321, -19.31502, -19.15649, 
    -18.9976, -18.83835, -18.67876, -18.51881, -18.3585, -18.19785, 
    -18.03683, -17.87547, -17.71375, -17.55167, -17.38924, -17.22646, 
    -17.06332, -16.89983, -16.73598, -16.57178, -16.40722, -16.24231, 
    -16.07704, -15.91142, -15.74545, -15.57912, -15.41244, -15.2454, 
    -15.07801, -14.91026, -14.74216, -14.57371, -14.40491, -14.23575, 
    -14.06624, -13.89638, -13.72617, -13.5556, -13.38468, -13.21342, 
    -13.0418, -12.86983, -12.69751, -12.52485, -12.35183, -12.17846, 
    -12.00475, -11.83069, -11.65629, -11.48154, -11.30644, -11.131, 
    -10.95521, -10.77908, -10.60261, -10.42579, -10.24864, -10.07114, 
    -9.893302, -9.715125, -9.53661, -9.357758, -9.178568, -8.999043, 
    -8.819182, -8.638988, -8.458461, -8.277601, -8.096411, -7.914891, 
    -7.733041, -7.550864, -7.368359, -7.185529, -7.002374, -6.818896, 
    -6.635096, -6.450974, -6.266533, -6.081773, -5.896696, -5.711303, 
    -5.525595, -5.339574, -5.153242, -4.966598, -4.779646, -4.592386, 
    -4.40482, -4.216949, -4.028776, -3.840301, -3.651526, -3.462453, 
    -3.273083, -3.083419, -2.893461, -2.703211, -2.512671, -2.321844, 
    -2.13073, -1.939332, -1.747651, -1.555689, -1.363449, -1.170931, 
    -0.9781384, -0.7850729, -0.5917361, -0.3981304, -0.2042576, -0.0101199, 
    0.1842807, 0.378942, 0.573862, 0.7690384, 0.964469, 1.160152, 1.356084, 
    1.552264, 1.74869, 1.945358, 2.142267, 2.339414, 2.536797, 2.734414, 
    2.932261, 3.130338, 3.32864, 3.527166, 3.725913, 3.924879, 4.124061, 
    4.323456, 4.523062, 4.722877, 4.922896, 5.123119, 5.323542, 5.524162, 
    5.724977, 5.925984, 6.127181, 6.328563, 6.530129, 6.731876, 6.933801, 
    7.135901, 7.338173, 7.540614, 7.743222, 7.945992, 8.148924, 8.352012, 
    8.555255, 8.758649, 8.962192, 9.165879, 9.36971, 9.573679, 9.777784, 
    9.982022, 10.18639, 10.39088, 10.5955, 10.80024, 11.0051, 11.21006, 
    11.41514, 11.62033, 11.82562, 12.03102, 12.23651, 12.44209, 12.64777, 
    12.85353, 13.05938, 13.26531, 13.47131, 13.6774, 13.88355, 14.08977, 
    14.29606, 14.5024, 14.70881, 14.91527, 15.12178, 15.32833, 15.53493, 
    15.74158, 15.94826, 16.15497, 16.36172, 16.56849, 16.77528, 16.9821, 
    17.18893, 17.39578, 17.60263, 17.8095, 18.01636, 18.22323, 18.43009, 
    18.63694, 18.84379, 19.05062, 19.25743, 19.46422, 19.67099, 19.87773, 
    20.08444, 20.29111, 20.49775, 20.70434, 20.91089, 21.1174, 21.32385, 
    21.53024, 21.73658, 21.94285, 22.14907, 22.35521, 22.56128, 22.76727, 
    22.97319, 23.17902, 23.38477, 23.59044, 23.79601, 24.00148, 24.20686, 
    24.41213, 24.6173, 24.82236, 25.02732, 25.23215, 25.43687, 25.64147, 
    25.84595, 26.05029, 26.25451, 26.4586, 26.66254, 26.86635, 27.07001, 
    27.27353, 27.4769, 27.68012, 27.88319, 28.08609, 28.28884, 28.49142, 
    28.69383, 28.89608, 29.09815, 29.30005, 29.50177, 29.7033, 29.90466, 
    30.10583, 30.3068, 30.50759, 30.70818, 30.90857, 31.10876, 31.30874, 
    31.50853, 31.7081, 31.90746, 32.10661, 32.30554, 32.50425, 32.70274, 
    32.90101, 33.09905, 33.29686, 33.49444, 33.69179, 33.8889, 34.08577, 
    34.2824, 34.47878, 34.67493, 34.87082, 35.06646, 35.26185, 35.45699, 
    35.65187, 35.84649, 36.04085, 36.23494, 36.42877, 36.62234, 36.81563, 
    37.00865, 37.2014, 37.39388, 37.58607, 37.77799, 37.96963, 38.16098, 
    38.35205, 38.54283, 38.73333, 38.92353, 39.11344, 39.30306, 39.49238, 
    39.68141, 39.87014, 40.05856, 40.24669, 40.43451, 40.62203, 40.80924, 
    40.99614, 41.18274, 41.36902, 41.55499, 41.74065, 41.92599, 42.11102, 
    42.29573, 42.48012, 42.66419, 42.84794, 43.03137, 43.21447, 43.39725, 
    43.5797, 43.76183, 43.94363, 44.1251, 44.30623, 44.48704, 44.66751, 
    44.84766, 45.02746, 45.20694, 45.38607, 45.56487, 45.74333, 45.92146, 
    46.09924, 46.27668, 46.45378, 46.63055, 46.80696, 46.98304, 47.15877, 
    47.33416, 47.5092, 47.6839, 47.85825, 48.03225, 48.20591, 48.37922, 
    48.55218, 48.72479, 48.89706, 49.06897, 49.24053, 49.41174, 49.5826, 
    49.75311, 49.92327, 50.09308, 50.26253, 50.43163, 50.60038, 50.76878, 
    50.93682,
  -29.11402, -28.97767, -28.841, -28.70402, -28.56672, -28.42909, -28.29115, 
    -28.15288, -28.01429, -27.87538, -27.73614, -27.59658, -27.4567, 
    -27.31648, -27.17594, -27.03507, -26.89388, -26.75235, -26.6105, 
    -26.46831, -26.32579, -26.18294, -26.03976, -25.89624, -25.75239, 
    -25.60821, -25.46369, -25.31883, -25.17364, -25.0281, -24.88224, 
    -24.73603, -24.58948, -24.44259, -24.29536, -24.14779, -23.99988, 
    -23.85163, -23.70303, -23.55409, -23.4048, -23.25517, -23.1052, 
    -22.95488, -22.80421, -22.6532, -22.50184, -22.35013, -22.19807, 
    -22.04567, -21.89292, -21.73981, -21.58636, -21.43255, -21.2784, 
    -21.12389, -20.96904, -20.81383, -20.65826, -20.50235, -20.34608, 
    -20.18946, -20.03248, -19.87516, -19.71747, -19.55943, -19.40104, 
    -19.2423, -19.08319, -18.92374, -18.76392, -18.60375, -18.44323, 
    -18.28234, -18.12111, -17.95951, -17.79756, -17.63525, -17.47259, 
    -17.30957, -17.14619, -16.98245, -16.81836, -16.65391, -16.48911, 
    -16.32395, -16.15843, -15.99255, -15.82632, -15.65973, -15.49278, 
    -15.32548, -15.15782, -14.9898, -14.82143, -14.65271, -14.48362, 
    -14.31419, -14.14439, -13.97425, -13.80375, -13.63289, -13.46168, 
    -13.29012, -13.11821, -12.94594, -12.77332, -12.60035, -12.42703, 
    -12.25335, -12.07933, -11.90496, -11.73023, -11.55516, -11.37974, 
    -11.20398, -11.02786, -10.8514, -10.6746, -10.49745, -10.31996, 
    -10.14212, -9.963939, -9.785418, -9.606555, -9.427353, -9.24781, 
    -9.06793, -8.887713, -8.707159, -8.526269, -8.345044, -8.163486, 
    -7.981596, -7.799373, -7.61682, -7.433938, -7.250728, -7.06719, 
    -6.883326, -6.699138, -6.514626, -6.329791, -6.144635, -5.95916, 
    -5.773366, -5.587255, -5.400828, -5.214087, -5.027033, -4.839667, 
    -4.651991, -4.464007, -4.275715, -4.087118, -3.898217, -3.709014, 
    -3.51951, -3.329707, -3.139606, -2.94921, -2.758519, -2.567537, 
    -2.376264, -2.184702, -1.992853, -1.800719, -1.608303, -1.415604, 
    -1.222627, -1.029372, -0.8358418, -0.6420382, -0.4479631, -0.2536188, 
    -0.05900715, 0.1358696, 0.3310094, 0.52641, 0.7220694, 0.9179852, 
    1.114155, 1.310577, 1.507249, 1.704168, 1.901333, 2.09874, 2.296387, 
    2.494273, 2.692394, 2.890748, 3.089333, 3.288146, 3.487185, 3.686446, 
    3.885929, 4.085629, 4.285545, 4.485673, 4.686012, 4.886558, 5.087308, 
    5.288261, 5.489413, 5.690761, 5.892303, 6.094037, 6.295958, 6.498064, 
    6.700353, 6.902822, 7.105466, 7.308285, 7.511275, 7.714432, 7.917754, 
    8.121239, 8.324882, 8.52868, 8.732632, 8.936732, 9.140981, 9.345372, 
    9.549904, 9.754573, 9.959375, 10.16431, 10.36937, 10.57456, 10.77987, 
    10.98529, 11.19083, 11.39649, 11.60225, 11.80811, 12.01408, 12.22015, 
    12.42631, 12.63257, 12.83891, 13.04534, 13.25185, 13.45844, 13.6651, 
    13.87184, 14.07864, 14.28551, 14.49244, 14.69944, 14.90648, 15.11358, 
    15.32072, 15.52791, 15.73514, 15.94241, 16.14971, 16.35704, 16.56441, 
    16.77179, 16.97919, 17.18662, 17.39405, 17.6015, 17.80895, 18.01641, 
    18.22386, 18.43132, 18.63876, 18.84619, 19.05361, 19.26102, 19.4684, 
    19.67575, 19.88308, 20.09038, 20.29764, 20.50487, 20.71205, 20.91919, 
    21.12627, 21.33331, 21.54029, 21.74721, 21.95407, 22.16087, 22.36759, 
    22.57425, 22.78082, 22.98732, 23.19374, 23.40006, 23.60631, 23.81245, 
    24.01851, 24.22446, 24.43031, 24.63605, 24.84169, 25.04721, 25.25262, 
    25.45791, 25.66307, 25.86812, 26.07303, 26.27781, 26.48246, 26.68697, 
    26.89134, 27.09556, 27.29964, 27.50357, 27.70734, 27.91096, 28.11442, 
    28.31771, 28.52085, 28.72381, 28.9266, 29.12922, 29.33166, 29.53392, 
    29.736, 29.93789, 30.13959, 30.3411, 30.54242, 30.74354, 30.94446, 
    31.14518, 31.34569, 31.546, 31.74609, 31.94597, 32.14564, 32.34509, 
    32.54432, 32.74332, 32.9421, 33.14064, 33.33896, 33.53704, 33.73489, 
    33.9325, 34.12987, 34.327, 34.52388, 34.72051, 34.91689, 35.11302, 
    35.3089, 35.50452, 35.69987, 35.89497, 36.08981, 36.28438, 36.47868, 
    36.67271, 36.86647, 37.05996, 37.25317, 37.44611, 37.63876, 37.83113, 
    38.02322, 38.21502, 38.40654, 38.59777, 38.7887, 38.97935, 39.1697, 
    39.35975, 39.54951, 39.73896, 39.92812, 40.11697, 40.30552, 40.49376, 
    40.6817, 40.86933, 41.05664, 41.24365, 41.43034, 41.61671, 41.80278, 
    41.98852, 42.17395, 42.35905, 42.54383, 42.72829, 42.91243, 43.09624, 
    43.27973, 43.46289, 43.64572, 43.82822, 44.01039, 44.19223, 44.37373, 
    44.5549, 44.73574, 44.91624, 45.09641, 45.27623, 45.45572, 45.63487, 
    45.81368, 45.99215, 46.17027, 46.34806, 46.52549, 46.70259, 46.87934, 
    47.05574, 47.2318, 47.40752, 47.58288, 47.7579, 47.93256, 48.10688, 
    48.28085, 48.45447, 48.62774, 48.80065, 48.97321, 49.14542, 49.31728, 
    49.48879, 49.65994, 49.83074, 50.00119, 50.17128, 50.34101, 50.5104, 
    50.67942, 50.84809, 51.0164,
  -29.21008, -29.07364, -28.93688, -28.7998, -28.6624, -28.52468, -28.38663, 
    -28.24827, -28.10958, -27.97056, -27.83122, -27.69155, -27.55155, 
    -27.41123, -27.27058, -27.1296, -26.98829, -26.84665, -26.70467, 
    -26.56237, -26.41973, -26.27676, -26.13345, -25.98981, -25.84583, 
    -25.70152, -25.55686, -25.41187, -25.26654, -25.12088, -24.97487, 
    -24.82852, -24.68183, -24.5348, -24.38743, -24.23971, -24.09165, 
    -23.94324, -23.79449, -23.6454, -23.49596, -23.34617, -23.19604, 
    -23.04556, -22.89472, -22.74355, -22.59202, -22.44014, -22.28791, 
    -22.13533, -21.9824, -21.82912, -21.67549, -21.5215, -21.36717, 
    -21.21247, -21.05743, -20.90203, -20.74628, -20.59017, -20.4337, 
    -20.27688, -20.11971, -19.96218, -19.80429, -19.64605, -19.48745, 
    -19.32849, -19.16917, -19.0095, -18.84947, -18.68908, -18.52833, 
    -18.36723, -18.20576, -18.04394, -17.88176, -17.71922, -17.55632, 
    -17.39306, -17.22944, -17.06547, -16.90113, -16.73643, -16.57138, 
    -16.40596, -16.24019, -16.07406, -15.90757, -15.74072, -15.57351, 
    -15.40594, -15.23801, -15.06973, -14.90108, -14.73208, -14.56272, 
    -14.393, -14.22293, -14.0525, -13.88171, -13.71056, -13.53906, -13.36721, 
    -13.19499, -13.02243, -12.84951, -12.67623, -12.5026, -12.32862, 
    -12.15428, -11.97959, -11.80455, -11.62916, -11.45342, -11.27733, 
    -11.10089, -10.9241, -10.74696, -10.56947, -10.39164, -10.21346, 
    -10.03494, -9.856074, -9.676865, -9.497311, -9.317416, -9.137179, 
    -8.956604, -8.775688, -8.594435, -8.412845, -8.230917, -8.048656, 
    -7.866059, -7.683129, -7.499868, -7.316276, -7.132354, -6.948103, 
    -6.763525, -6.578621, -6.393392, -6.207839, -6.021964, -5.835768, 
    -5.649252, -5.462418, -5.275266, -5.0878, -4.900019, -4.711926, 
    -4.523521, -4.334807, -4.145784, -3.956456, -3.766822, -3.576886, 
    -3.386647, -3.196109, -3.005273, -2.81414, -2.622712, -2.430991, 
    -2.238979, -2.046678, -1.85409, -1.661216, -1.468058, -1.274618, 
    -1.080899, -0.886902, -0.6926292, -0.4980826, -0.3032644, -0.1081766, 
    0.08717857, 0.2827991, 0.4786828, 0.6748274, 0.8712308, 1.067891, 
    1.264805, 1.461971, 1.659386, 1.857049, 2.054957, 2.253108, 2.451498, 
    2.650126, 2.848989, 3.048086, 3.247412, 3.446966, 3.646745, 3.846747, 
    4.046968, 4.247407, 4.448061, 4.648927, 4.850001, 5.051283, 5.252768, 
    5.454455, 5.65634, 5.85842, 6.060693, 6.263155, 6.465805, 6.668639, 
    6.871654, 7.074848, 7.278216, 7.481757, 7.685468, 7.889345, 8.093385, 
    8.297585, 8.501943, 8.706455, 8.911118, 9.115929, 9.320885, 9.525983, 
    9.731218, 9.93659, 10.14209, 10.34773, 10.55349, 10.75937, 10.96537, 
    11.17148, 11.37771, 11.58405, 11.7905, 11.99705, 12.20369, 12.41044, 
    12.61727, 12.8242, 13.03121, 13.23831, 13.44548, 13.65273, 13.86005, 
    14.06745, 14.27491, 14.48243, 14.69, 14.89764, 15.10533, 15.31306, 
    15.52084, 15.72866, 15.93652, 16.14442, 16.35234, 16.5603, 16.76828, 
    16.97627, 17.18429, 17.39232, 17.60036, 17.8084, 18.01645, 18.2245, 
    18.43255, 18.64059, 18.84862, 19.05663, 19.26462, 19.4726, 19.68055, 
    19.88847, 20.09636, 20.30421, 20.51203, 20.7198, 20.92753, 21.13521, 
    21.34283, 21.55041, 21.75792, 21.96536, 22.17274, 22.38006, 22.5873, 
    22.79446, 23.00154, 23.20854, 23.41545, 23.62227, 23.829, 24.03563, 
    24.24217, 24.4486, 24.65492, 24.86113, 25.06723, 25.27321, 25.47907, 
    25.68481, 25.89042, 26.09591, 26.30126, 26.50647, 26.71155, 26.91648, 
    27.12127, 27.3259, 27.53039, 27.73473, 27.9389, 28.14292, 28.34677, 
    28.55045, 28.75397, 28.95731, 29.16047, 29.36346, 29.56626, 29.76888, 
    29.97132, 30.17356, 30.37561, 30.57746, 30.77912, 30.98057, 31.18182, 
    31.38286, 31.58369, 31.78431, 31.98472, 32.18491, 32.38487, 32.58461, 
    32.78413, 32.98343, 33.18248, 33.38131, 33.5799, 33.77825, 33.97636, 
    34.17423, 34.37186, 34.56923, 34.76636, 34.96323, 35.15985, 35.35622, 
    35.55232, 35.74816, 35.94374, 36.13905, 36.3341, 36.52887, 36.72338, 
    36.91761, 37.11156, 37.30524, 37.49863, 37.69175, 37.88457, 38.07712, 
    38.26937, 38.46134, 38.65301, 38.84439, 39.03548, 39.22627, 39.41676, 
    39.60695, 39.79684, 39.98642, 40.1757, 40.36468, 40.55334, 40.7417, 
    40.92974, 41.11747, 41.30489, 41.49199, 41.67878, 41.86524, 42.05139, 
    42.23721, 42.42271, 42.60789, 42.79274, 42.97727, 43.16147, 43.34534, 
    43.52888, 43.71209, 43.89497, 44.07751, 44.25972, 44.44159, 44.62313, 
    44.80433, 44.98519, 45.16571, 45.34589, 45.52574, 45.70523, 45.88439, 
    46.06321, 46.24167, 46.4198, 46.59757, 46.775, 46.95208, 47.12882, 
    47.30521, 47.48124, 47.65693, 47.83226, 48.00725, 48.18188, 48.35616, 
    48.53009, 48.70366, 48.87688, 49.04975, 49.22226, 49.39442, 49.56622, 
    49.73766, 49.90875, 50.07948, 50.24986, 50.41988, 50.58953, 50.75884, 
    50.92778, 51.09637,
  -29.30649, -29.16996, -29.0331, -28.89593, -28.75843, -28.62062, -28.48247, 
    -28.34401, -28.20521, -28.0661, -27.92665, -27.78687, -27.64677, 
    -27.50634, -27.36558, -27.22449, -27.08306, -26.9413, -26.79921, 
    -26.65679, -26.51403, -26.37094, -26.2275, -26.08374, -25.93963, 
    -25.79519, -25.65041, -25.50528, -25.35982, -25.21402, -25.06787, 
    -24.92138, -24.77456, -24.62738, -24.47986, -24.332, -24.18379, 
    -24.03524, -23.88634, -23.73709, -23.58749, -23.43754, -23.28725, 
    -23.13661, -22.98561, -22.83427, -22.68258, -22.53053, -22.37813, 
    -22.22538, -22.07227, -21.91882, -21.765, -21.61084, -21.45632, 
    -21.30144, -21.14621, -20.99062, -20.83467, -20.67837, -20.52171, 
    -20.36469, -20.20732, -20.04959, -19.8915, -19.73305, -19.57424, 
    -19.41507, -19.25554, -19.09565, -18.93541, -18.7748, -18.61383, 
    -18.4525, -18.29081, -18.12876, -17.96634, -17.80357, -17.64044, 
    -17.47694, -17.31308, -17.14886, -16.98428, -16.81934, -16.65404, 
    -16.48837, -16.32234, -16.15595, -15.9892, -15.82209, -15.65462, 
    -15.48679, -15.31859, -15.15003, -14.98112, -14.81184, -14.6422, 
    -14.47221, -14.30185, -14.13113, -13.96006, -13.78862, -13.61683, 
    -13.44467, -13.27216, -13.0993, -12.92607, -12.75249, -12.57855, 
    -12.40426, -12.22961, -12.0546, -11.87925, -11.70353, -11.52747, 
    -11.35105, -11.17428, -10.99716, -10.81969, -10.64187, -10.4637, 
    -10.28518, -10.10631, -9.9271, -9.74754, -9.567636, -9.387386, -9.206793, 
    -9.025858, -8.84458, -8.662962, -8.481004, -8.298707, -8.116073, 
    -7.933101, -7.749794, -7.566152, -7.382176, -7.197869, -7.01323, 
    -6.828261, -6.642963, -6.457338, -6.271387, -6.085111, -5.898511, 
    -5.711588, -5.524345, -5.336783, -5.148902, -4.960704, -4.772192, 
    -4.583365, -4.394227, -4.204778, -4.01502, -3.824955, -3.634583, 
    -3.443908, -3.25293, -3.061651, -2.870074, -2.678199, -2.486029, 
    -2.293566, -2.10081, -1.907765, -1.714431, -1.520812, -1.326908, 
    -1.132722, -0.938256, -0.7435119, -0.5484916, -0.3531973, -0.1576311, 
    0.03820484, 0.2343084, 0.4306775, 0.6273098, 0.8242031, 1.021355, 
    1.218764, 1.416426, 1.614341, 1.812505, 2.010916, 2.209572, 2.40847, 
    2.607608, 2.806983, 3.006593, 3.206436, 3.406508, 3.606807, 3.807331, 
    4.008076, 4.209042, 4.410223, 4.611619, 4.813225, 5.015041, 5.217062, 
    5.419286, 5.62171, 5.824331, 6.027147, 6.230155, 6.433351, 6.636733, 
    6.840298, 7.044042, 7.247964, 7.45206, 7.656326, 7.860761, 8.06536, 
    8.270122, 8.475041, 8.680118, 8.885345, 9.090723, 9.296247, 9.501914, 
    9.707721, 9.913665, 10.11974, 10.32595, 10.53228, 10.73874, 10.94532, 
    11.15201, 11.35882, 11.56574, 11.77277, 11.9799, 12.18713, 12.39446, 
    12.60188, 12.8094, 13.017, 13.22468, 13.43244, 13.64028, 13.8482, 
    14.05618, 14.26423, 14.47234, 14.68052, 14.88874, 15.09702, 15.30535, 
    15.51373, 15.72215, 15.9306, 16.13909, 16.34761, 16.55617, 16.76474, 
    16.97334, 17.18195, 17.39058, 17.59921, 17.80786, 18.0165, 18.22515, 
    18.43379, 18.64243, 18.85105, 19.05966, 19.26826, 19.47683, 19.68537, 
    19.89389, 20.10238, 20.31082, 20.51924, 20.7276, 20.93592, 21.1442, 
    21.35242, 21.56058, 21.76868, 21.97672, 22.1847, 22.3926, 22.60043, 
    22.80818, 23.01585, 23.22343, 23.43093, 23.63834, 23.84565, 24.05287, 
    24.25998, 24.467, 24.6739, 24.88069, 25.08737, 25.29393, 25.50036, 
    25.70668, 25.91286, 26.11892, 26.32484, 26.53063, 26.73627, 26.94177, 
    27.14713, 27.35233, 27.55738, 27.76228, 27.96701, 28.17159, 28.376, 
    28.58024, 28.78431, 28.9882, 29.19192, 29.39545, 29.5988, 29.80197, 
    30.00495, 30.20773, 30.41032, 30.61272, 30.81491, 31.0169, 31.21868, 
    31.42025, 31.62161, 31.82276, 32.02369, 32.2244, 32.42489, 32.62516, 
    32.82519, 33.025, 33.22457, 33.42391, 33.62301, 33.82187, 34.02048, 
    34.21886, 34.41698, 34.61486, 34.81248, 35.00985, 35.20696, 35.40381, 
    35.6004, 35.79673, 35.99279, 36.18858, 36.38411, 36.57936, 36.77433, 
    36.96904, 37.16346, 37.3576, 37.55146, 37.74503, 37.93832, 38.13132, 
    38.32403, 38.51645, 38.70857, 38.9004, 39.09193, 39.28316, 39.47409, 
    39.66472, 39.85504, 40.04506, 40.23477, 40.42417, 40.61325, 40.80203, 
    40.99049, 41.17864, 41.36647, 41.55399, 41.74118, 41.92805, 42.1146, 
    42.30082, 42.48672, 42.6723, 42.85754, 43.04246, 43.22705, 43.4113, 
    43.59522, 43.77881, 43.96207, 44.14499, 44.32756, 44.50981, 44.69172, 
    44.87328, 45.0545, 45.23538, 45.41592, 45.59612, 45.77597, 45.95547, 
    46.13463, 46.31344, 46.49191, 46.67002, 46.84779, 47.0252, 47.20227, 
    47.37898, 47.55534, 47.73135, 47.90701, 48.08231, 48.25726, 48.43185, 
    48.60609, 48.77997, 48.9535, 49.12666, 49.29948, 49.47193, 49.64402, 
    49.81576, 49.98714, 50.15816, 50.32882, 50.49912, 50.66906, 50.83864, 
    51.00786, 51.17672,
  -29.40325, -29.26662, -29.12968, -28.99241, -28.85482, -28.71691, 
    -28.57867, -28.4401, -28.30121, -28.16199, -28.02244, -27.88256, 
    -27.74235, -27.60181, -27.46094, -27.31973, -27.1782, -27.03632, 
    -26.89412, -26.75157, -26.6087, -26.46548, -26.32193, -26.17803, 
    -26.0338, -25.88923, -25.74432, -25.59907, -25.45347, -25.30753, 
    -25.16125, -25.01462, -24.86765, -24.72034, -24.57267, -24.42467, 
    -24.27631, -24.12761, -23.97855, -23.82915, -23.6794, -23.5293, 
    -23.37885, -23.22804, -23.07689, -22.92537, -22.77351, -22.6213, 
    -22.46873, -22.31581, -22.16253, -22.00889, -21.8549, -21.70055, 
    -21.54585, -21.39079, -21.23537, -21.07959, -20.92346, -20.76696, 
    -20.61011, -20.45289, -20.29532, -20.13738, -19.97909, -19.82043, 
    -19.66142, -19.50204, -19.3423, -19.18219, -19.02173, -18.8609, 
    -18.69971, -18.53816, -18.37624, -18.21396, -18.05132, -17.88832, 
    -17.72495, -17.56121, -17.39711, -17.23265, -17.06783, -16.90264, 
    -16.73708, -16.57117, -16.40489, -16.23824, -16.07123, -15.90386, 
    -15.73612, -15.56802, -15.39956, -15.23073, -15.06154, -14.89199, 
    -14.72207, -14.55179, -14.38115, -14.21015, -14.03879, -13.86706, 
    -13.69497, -13.52252, -13.34972, -13.17655, -13.00302, -12.82913, 
    -12.65489, -12.48028, -12.30532, -12.13, -11.95432, -11.77829, -11.6019, 
    -11.42515, -11.24806, -11.0706, -10.8928, -10.71464, -10.53613, 
    -10.35727, -10.17806, -9.998497, -9.818587, -9.63833, -9.457725, 
    -9.276773, -9.095477, -8.913836, -8.731853, -8.549526, -8.366858, 
    -8.18385, -8.000503, -7.816816, -7.632792, -7.448433, -7.263739, 
    -7.07871, -6.893349, -6.707657, -6.521635, -6.335283, -6.148604, 
    -5.961599, -5.774269, -5.586615, -5.398639, -5.210343, -5.021727, 
    -4.832794, -4.643544, -4.453979, -4.264102, -4.073913, -3.883413, 
    -3.692606, -3.501492, -3.310072, -3.11835, -2.926326, -2.734002, 
    -2.541381, -2.348463, -2.155251, -1.961747, -1.767952, -1.573869, 
    -1.379499, -1.184844, -0.9899068, -0.7946891, -0.5991929, -0.4034203, 
    -0.2073734, -0.01105434, 0.1855347, 0.3823915, 0.5795139, 0.7768996, 
    0.9745463, 1.172452, 1.370614, 1.56903, 1.767697, 1.966614, 2.165778, 
    2.365187, 2.564837, 2.764727, 2.964853, 3.165215, 3.365807, 3.566629, 
    3.767678, 3.968951, 4.170445, 4.372158, 4.574086, 4.776227, 4.97858, 
    5.181139, 5.383904, 5.58687, 5.790036, 5.993397, 6.196953, 6.400698, 
    6.604631, 6.808749, 7.013049, 7.217526, 7.42218, 7.627007, 7.832002, 
    8.037164, 8.24249, 8.447975, 8.653618, 8.859415, 9.065362, 9.271458, 
    9.477697, 9.684077, 9.890596, 10.09725, 10.30404, 10.51095, 10.71799, 
    10.92515, 11.13242, 11.33982, 11.54732, 11.75493, 11.96265, 12.17047, 
    12.37839, 12.5864, 12.7945, 13.00269, 13.21097, 13.41932, 13.62776, 
    13.83627, 14.04484, 14.25349, 14.4622, 14.67097, 14.87979, 15.08867, 
    15.2976, 15.50657, 15.71559, 15.92464, 16.13373, 16.34286, 16.55201, 
    16.76118, 16.97038, 17.17959, 17.38882, 17.59806, 17.8073, 18.01655, 
    18.2258, 18.43504, 18.64428, 18.8535, 19.06272, 19.27191, 19.48108, 
    19.69023, 19.89934, 20.10843, 20.31748, 20.52649, 20.73545, 20.94437, 
    21.15324, 21.36206, 21.57082, 21.77952, 21.98815, 22.19672, 22.40522, 
    22.61364, 22.82198, 23.03024, 23.23842, 23.44651, 23.65451, 23.86241, 
    24.07021, 24.27791, 24.48551, 24.693, 24.90037, 25.10763, 25.31477, 
    25.52179, 25.72868, 25.93545, 26.14208, 26.34858, 26.55494, 26.76115, 
    26.96723, 27.17315, 27.37892, 27.58454, 27.79, 27.9953, 28.20044, 
    28.40541, 28.6102, 28.81483, 29.01928, 29.22355, 29.42764, 29.63154, 
    29.83526, 30.03878, 30.24212, 30.44525, 30.64818, 30.85092, 31.05344, 
    31.25576, 31.45787, 31.65977, 31.86144, 32.0629, 32.26414, 32.46515, 
    32.66594, 32.86649, 33.06682, 33.26691, 33.46676, 33.66637, 33.86574, 
    34.06487, 34.26374, 34.46237, 34.66075, 34.85887, 35.05674, 35.25434, 
    35.45169, 35.64877, 35.84558, 36.04213, 36.2384, 36.43441, 36.63013, 
    36.82559, 37.02076, 37.21565, 37.41026, 37.60459, 37.79863, 37.99237, 
    38.18583, 38.379, 38.57187, 38.76445, 38.95672, 39.1487, 39.34037, 
    39.53174, 39.72281, 39.91357, 40.10402, 40.29416, 40.48399, 40.6735, 
    40.8627, 41.05158, 41.24015, 41.42839, 41.61632, 41.80392, 41.9912, 
    42.17815, 42.36478, 42.55108, 42.73705, 42.92269, 43.108, 43.29298, 
    43.47762, 43.66193, 43.84589, 44.02953, 44.21282, 44.39577, 44.57839, 
    44.76066, 44.94259, 45.12418, 45.30542, 45.48632, 45.66687, 45.84707, 
    46.02692, 46.20643, 46.38559, 46.56439, 46.74284, 46.92095, 47.0987, 
    47.27609, 47.45314, 47.62983, 47.80616, 47.98213, 48.15775, 48.33302, 
    48.50792, 48.68247, 48.85666, 49.03049, 49.20396, 49.37708, 49.54983, 
    49.72222, 49.89425, 50.06592, 50.23722, 50.40817, 50.57875, 50.74897, 
    50.91883, 51.08833, 51.25746,
  -29.50036, -29.36365, -29.22661, -29.08925, -28.95157, -28.81356, 
    -28.67522, -28.53656, -28.39757, -28.25824, -28.11859, -27.97861, 
    -27.83829, -27.69764, -27.55666, -27.41535, -27.2737, -27.13171, 
    -26.98939, -26.84673, -26.70373, -26.56039, -26.41672, -26.2727, 
    -26.12835, -25.98365, -25.8386, -25.69322, -25.54749, -25.40142, -25.255, 
    -25.10824, -24.96113, -24.81367, -24.66586, -24.51771, -24.36921, 
    -24.22035, -24.07115, -23.9216, -23.77169, -23.62143, -23.47082, 
    -23.31986, -23.16854, -23.01686, -22.86484, -22.71245, -22.55972, 
    -22.40662, -22.25317, -22.09935, -21.94519, -21.79066, -21.63577, 
    -21.48053, -21.32492, -21.16895, -21.01263, -20.85594, -20.69889, 
    -20.54148, -20.38371, -20.22557, -20.06707, -19.90821, -19.74899, 
    -19.5894, -19.42945, -19.26913, -19.10845, -18.9474, -18.78599, 
    -18.62421, -18.46207, -18.29956, -18.13669, -17.97345, -17.80984, 
    -17.64587, -17.48154, -17.31683, -17.15176, -16.98633, -16.82052, 
    -16.65436, -16.48782, -16.32092, -16.15365, -15.98602, -15.81802, 
    -15.64965, -15.48092, -15.31182, -15.14236, -14.97253, -14.80233, 
    -14.63177, -14.46085, -14.28956, -14.11791, -13.94589, -13.77351, 
    -13.60076, -13.42766, -13.25419, -13.08035, -12.90616, -12.73161, 
    -12.55669, -12.38141, -12.20578, -12.02978, -11.85342, -11.67671, 
    -11.49964, -11.32221, -11.14443, -10.96628, -10.78779, -10.60894, 
    -10.42973, -10.25018, -10.07027, -9.890007, -9.709395, -9.528435, 
    -9.347125, -9.165467, -8.983462, -8.801111, -8.618415, -8.435375, 
    -8.251991, -8.068266, -7.8842, -7.699794, -7.515049, -7.329966, 
    -7.144547, -6.958792, -6.772704, -6.586283, -6.399529, -6.212447, 
    -6.025035, -5.837295, -5.64923, -5.460839, -5.272125, -5.08309, 
    -4.893734, -4.704059, -4.514067, -4.323759, -4.133136, -3.942202, 
    -3.750956, -3.559401, -3.367539, -3.175371, -2.982898, -2.790124, 
    -2.597049, -2.403675, -2.210005, -2.016039, -1.821781, -1.627232, 
    -1.432393, -1.237268, -1.041857, -0.8461638, -0.6501894, -0.4539362, 
    -0.2574062, -0.06060177, 0.1364751, 0.333822, 0.5314369, 0.7293174, 
    0.9274613, 1.125866, 1.32453, 1.52345, 1.722624, 1.922049, 2.121724, 
    2.321645, 2.521811, 2.722218, 2.922863, 3.123746, 3.324862, 3.52621, 
    3.727787, 3.929589, 4.131615, 4.333862, 4.536326, 4.739005, 4.941897, 
    5.144998, 5.348306, 5.551818, 5.755531, 5.959442, 6.163548, 6.367846, 
    6.572334, 6.777008, 6.981865, 7.186902, 7.392117, 7.597506, 7.803066, 
    8.008794, 8.214686, 8.420741, 8.626954, 8.833323, 9.039844, 9.246513, 
    9.453329, 9.660288, 9.867385, 10.07462, 10.28199, 10.48948, 10.6971, 
    10.90485, 11.11271, 11.32069, 11.52878, 11.73699, 11.94529, 12.1537, 
    12.36221, 12.57082, 12.77951, 12.9883, 13.19717, 13.40612, 13.61515, 
    13.82426, 14.03344, 14.24268, 14.45199, 14.66136, 14.87078, 15.08026, 
    15.28979, 15.49937, 15.70899, 15.91865, 16.12834, 16.33807, 16.54782, 
    16.7576, 16.9674, 17.17722, 17.38705, 17.5969, 17.80674, 18.0166, 
    18.22645, 18.4363, 18.64614, 18.85597, 19.06579, 19.27559, 19.48536, 
    19.69511, 19.90483, 20.11452, 20.32417, 20.53378, 20.74335, 20.95288, 
    21.16235, 21.37177, 21.58112, 21.79042, 21.99966, 22.20882, 22.41792, 
    22.62693, 22.83587, 23.04473, 23.2535, 23.46219, 23.67078, 23.87927, 
    24.08767, 24.29596, 24.50414, 24.71222, 24.92018, 25.12802, 25.33575, 
    25.54335, 25.75083, 25.95817, 26.16538, 26.37246, 26.5794, 26.78619, 
    26.99283, 27.19933, 27.40568, 27.61186, 27.81789, 28.02376, 28.22946, 
    28.435, 28.64036, 28.84554, 29.05055, 29.25538, 29.46003, 29.66448, 
    29.86875, 30.07283, 30.27671, 30.48039, 30.68387, 30.88714, 31.09021, 
    31.29307, 31.49571, 31.69814, 31.90036, 32.10235, 32.30412, 32.50565, 
    32.70697, 32.90805, 33.10889, 33.3095, 33.50987, 33.71, 33.90988, 
    34.10951, 34.3089, 34.50803, 34.70691, 34.90554, 35.1039, 35.302, 
    35.49984, 35.69741, 35.89472, 36.09175, 36.28851, 36.485, 36.68121, 
    36.87714, 37.07279, 37.26815, 37.46323, 37.65802, 37.85253, 38.04674, 
    38.24066, 38.43428, 38.62761, 38.82064, 39.01336, 39.20579, 39.39791, 
    39.58972, 39.78123, 39.97242, 40.16331, 40.35388, 40.54414, 40.73409, 
    40.92371, 41.11301, 41.302, 41.49066, 41.679, 41.86702, 42.0547, 
    42.24206, 42.42909, 42.6158, 42.80216, 42.9882, 43.1739, 43.35926, 
    43.5443, 43.72898, 43.91334, 44.09735, 44.28102, 44.46435, 44.64734, 
    44.82998, 45.01228, 45.19423, 45.37583, 45.55708, 45.73799, 45.91854, 
    46.09875, 46.2786, 46.4581, 46.63725, 46.81605, 46.99449, 47.17257, 
    47.3503, 47.52767, 47.70469, 47.88134, 48.05764, 48.23358, 48.40916, 
    48.58438, 48.75924, 48.93374, 49.10788, 49.28165, 49.45506, 49.62811, 
    49.8008, 49.97313, 50.14508, 50.31668, 50.48791, 50.65878, 50.82928, 
    50.99942, 51.16919, 51.33859,
  -29.59783, -29.46103, -29.3239, -29.18645, -29.04868, -28.91057, -28.77214, 
    -28.63338, -28.49428, -28.35486, -28.21511, -28.07502, -27.9346, 
    -27.79384, -27.65275, -27.51133, -27.36957, -27.22747, -27.08503, 
    -26.94225, -26.79914, -26.65568, -26.51188, -26.36774, -26.22326, 
    -26.07844, -25.93327, -25.78775, -25.64189, -25.49569, -25.34913, 
    -25.20223, -25.05498, -24.90738, -24.75943, -24.61114, -24.46249, 
    -24.31348, -24.16413, -24.01443, -23.86436, -23.71395, -23.56318, 
    -23.41206, -23.26058, -23.10874, -22.95655, -22.804, -22.65109, 
    -22.49782, -22.34419, -22.19021, -22.03586, -21.88115, -21.72609, 
    -21.57066, -21.41486, -21.25871, -21.10219, -20.94531, -20.78807, 
    -20.63046, -20.47249, -20.31415, -20.15545, -19.99639, -19.83695, 
    -19.67715, -19.51699, -19.35646, -19.19556, -19.03429, -18.87266, 
    -18.71066, -18.54829, -18.38556, -18.22245, -18.05898, -17.89514, 
    -17.73093, -17.56636, -17.40141, -17.2361, -17.07041, -16.90436, 
    -16.73794, -16.57115, -16.40399, -16.23647, -16.06857, -15.90031, 
    -15.73167, -15.56267, -15.3933, -15.22357, -15.05346, -14.88299, 
    -14.71215, -14.54094, -14.36936, -14.19742, -14.02511, -13.85244, 
    -13.6794, -13.50599, -13.33222, -13.15808, -12.98358, -12.80871, 
    -12.63348, -12.45789, -12.28194, -12.10562, -11.92894, -11.75191, 
    -11.57451, -11.39675, -11.21863, -11.04015, -10.86132, -10.68213, 
    -10.50258, -10.32267, -10.14242, -9.961803, -9.780838, -9.59952, 
    -9.41785, -9.235829, -9.053459, -8.87074, -8.687674, -8.50426, -8.3205, 
    -8.136396, -7.951949, -7.767159, -7.582026, -7.396554, -7.210743, 
    -7.024594, -6.838108, -6.651286, -6.46413, -6.276642, -6.088822, 
    -5.900671, -5.712192, -5.523386, -5.334253, -5.144795, -4.955016, 
    -4.764914, -4.574492, -4.383752, -4.192695, -4.001323, -3.809638, 
    -3.61764, -3.425333, -3.232717, -3.039794, -2.846567, -2.653036, 
    -2.459205, -2.265074, -2.070645, -1.875921, -1.680904, -1.485595, 
    -1.289997, -1.09411, -0.8979389, -0.701484, -0.5047478, -0.3077325, 
    -0.1104403, 0.08712672, 0.2849663, 0.4830761, 0.6814539, 0.8800974, 
    1.079004, 1.278172, 1.477599, 1.677281, 1.877218, 2.077406, 2.277843, 
    2.478526, 2.679453, 2.880621, 3.082028, 3.283671, 3.485547, 3.687654, 
    3.88999, 4.09255, 4.295333, 4.498336, 4.701557, 4.904991, 5.108637, 
    5.312491, 5.516551, 5.720815, 5.925278, 6.129938, 6.334792, 6.539837, 
    6.74507, 6.950489, 7.156089, 7.361868, 7.567823, 7.773951, 7.980247, 
    8.186711, 8.393338, 8.600125, 8.807069, 9.014167, 9.221415, 9.42881, 
    9.636349, 9.844028, 10.05185, 10.2598, 10.46788, 10.67609, 10.88442, 
    11.09287, 11.30145, 11.51013, 11.71892, 11.92783, 12.13683, 12.34594, 
    12.55514, 12.76443, 12.97382, 13.18329, 13.39284, 13.60247, 13.81218, 
    14.02196, 14.2318, 14.44172, 14.65169, 14.86172, 15.0718, 15.28194, 
    15.49212, 15.70235, 15.91261, 16.12291, 16.33325, 16.54361, 16.754, 
    16.96441, 17.17483, 17.38527, 17.59573, 17.80618, 18.01665, 18.22711, 
    18.43756, 18.64802, 18.85846, 19.06888, 19.27929, 19.48967, 19.70003, 
    19.91035, 20.12065, 20.33091, 20.54113, 20.7513, 20.96143, 21.17151, 
    21.38153, 21.59149, 21.8014, 22.01123, 22.221, 22.43069, 22.64031, 
    22.84985, 23.05931, 23.26868, 23.47796, 23.68715, 23.89624, 24.10523, 
    24.31411, 24.52289, 24.73156, 24.94011, 25.14854, 25.35686, 25.56504, 
    25.77311, 25.98104, 26.18883, 26.39649, 26.60401, 26.81138, 27.0186, 
    27.22568, 27.4326, 27.63936, 27.84596, 28.0524, 28.25867, 28.46477, 
    28.67069, 28.87645, 29.08202, 29.28741, 29.49261, 29.69763, 29.90245, 
    30.10708, 30.31151, 30.51574, 30.71977, 30.92359, 31.1272, 31.3306, 
    31.53379, 31.73676, 31.93951, 32.14203, 32.34433, 32.5464, 32.74824, 
    32.94985, 33.15121, 33.35235, 33.55323, 33.75388, 33.95428, 34.15443, 
    34.35432, 34.55396, 34.75335, 34.95248, 35.15134, 35.34995, 35.54828, 
    35.74635, 35.94415, 36.14167, 36.33892, 36.53589, 36.73258, 36.92899, 
    37.12511, 37.32096, 37.51651, 37.71177, 37.90674, 38.10142, 38.2958, 
    38.48989, 38.68367, 38.87715, 39.07033, 39.26321, 39.45577, 39.64803, 
    39.83998, 40.03162, 40.22294, 40.41394, 40.60463, 40.79501, 40.98506, 
    41.17479, 41.36419, 41.55327, 41.74203, 41.93045, 42.11855, 42.30632, 
    42.49376, 42.68086, 42.86763, 43.05406, 43.24016, 43.42591, 43.61134, 
    43.79641, 43.98115, 44.16554, 44.34959, 44.53329, 44.71666, 44.89967, 
    45.08233, 45.26464, 45.44661, 45.62822, 45.80949, 45.9904, 46.17095, 
    46.35115, 46.531, 46.71049, 46.88963, 47.06841, 47.24683, 47.42489, 
    47.60259, 47.77993, 47.95692, 48.13354, 48.3098, 48.48569, 48.66123, 
    48.8364, 49.01121, 49.18565, 49.35973, 49.53344, 49.70679, 49.87978, 
    50.05239, 50.22464, 50.39653, 50.56804, 50.73919, 50.90998, 51.08039, 
    51.25044, 51.42012,
  -29.69565, -29.55877, -29.42155, -29.28401, -29.14614, -29.00794, 
    -28.86941, -28.73055, -28.59136, -28.45184, -28.31199, -28.17179, 
    -28.03127, -27.89041, -27.74921, -27.60768, -27.46581, -27.32359, 
    -27.18104, -27.03815, -26.89492, -26.75134, -26.60742, -26.46316, 
    -26.31855, -26.1736, -26.02831, -25.88266, -25.73667, -25.59033, 
    -25.44364, -25.2966, -25.14922, -25.00148, -24.85339, -24.70494, 
    -24.55615, -24.407, -24.2575, -24.10764, -23.95743, -23.80686, -23.65593, 
    -23.50465, -23.35301, -23.20101, -23.04865, -22.89593, -22.74285, 
    -22.58941, -22.43561, -22.28145, -22.12693, -21.97204, -21.81679, 
    -21.66118, -21.5052, -21.34886, -21.19215, -21.03508, -20.87764, 
    -20.71984, -20.56167, -20.40313, -20.24423, -20.08496, -19.92531, 
    -19.76531, -19.60493, -19.44418, -19.28307, -19.12159, -18.95973, 
    -18.79751, -18.63491, -18.47195, -18.30862, -18.14491, -17.98084, 
    -17.81639, -17.65158, -17.48639, -17.32083, -17.1549, -16.9886, 
    -16.82192, -16.65488, -16.48747, -16.31968, -16.15152, -15.983, -15.8141, 
    -15.64482, -15.47518, -15.30517, -15.13479, -14.96404, -14.79292, 
    -14.62142, -14.44956, -14.27733, -14.10473, -13.93176, -13.75842, 
    -13.58471, -13.41064, -13.2362, -13.06139, -12.88621, -12.71067, 
    -12.53477, -12.35849, -12.18186, -12.00485, -11.82749, -11.64976, 
    -11.47167, -11.29322, -11.11441, -10.93523, -10.7557, -10.57581, 
    -10.39555, -10.21495, -10.03398, -9.852659, -9.670982, -9.488952, 
    -9.306567, -9.123831, -8.940743, -8.757304, -8.573517, -8.38938, 
    -8.204896, -8.020065, -7.83489, -7.64937, -7.463507, -7.277302, 
    -7.090756, -6.903872, -6.716649, -6.529088, -6.341193, -6.152963, 
    -5.9644, -5.775506, -5.586281, -5.396729, -5.206848, -5.016642, 
    -4.826112, -4.635259, -4.444085, -4.252592, -4.060781, -3.868653, 
    -3.676212, -3.483457, -3.290391, -3.097017, -2.903334, -2.709347, 
    -2.515055, -2.320461, -2.125568, -1.930376, -1.734889, -1.539107, 
    -1.343033, -1.146669, -0.9500172, -0.7530795, -0.5558581, -0.3583551, 
    -0.1605727, 0.03748685, 0.2358214, 0.4344286, 0.6333061, 0.8324518, 
    1.031863, 1.231538, 1.431474, 1.631668, 1.832118, 2.032822, 2.233777, 
    2.434981, 2.636431, 2.838124, 3.040058, 3.24223, 3.444638, 3.647278, 
    3.850149, 4.053247, 4.25657, 4.460115, 4.663879, 4.867859, 5.072052, 
    5.276457, 5.481069, 5.685885, 5.890904, 6.096121, 6.301534, 6.50714, 
    6.712936, 6.918918, 7.125084, 7.331431, 7.537955, 7.744654, 7.951524, 
    8.158562, 8.365765, 8.573129, 8.780651, 8.988329, 9.196158, 9.404137, 
    9.612261, 9.820526, 10.02893, 10.23747, 10.44614, 10.65494, 10.86387, 
    11.07291, 11.28208, 11.49136, 11.70075, 11.91025, 12.11985, 12.32956, 
    12.53936, 12.74925, 12.95924, 13.16931, 13.37947, 13.58971, 13.80002, 
    14.0104, 14.22086, 14.43138, 14.64196, 14.8526, 15.06329, 15.27404, 
    15.48483, 15.69566, 15.90654, 16.11745, 16.3284, 16.53937, 16.75037, 
    16.96139, 17.17243, 17.38348, 17.59455, 17.80562, 18.0167, 18.22777, 
    18.43884, 18.6499, 18.86095, 19.07199, 19.28301, 19.494, 19.70497, 
    19.91591, 20.12682, 20.33769, 20.54852, 20.7593, 20.97004, 21.18073, 
    21.39136, 21.60193, 21.81244, 22.02288, 22.23326, 22.44356, 22.65378, 
    22.86392, 23.07398, 23.28395, 23.49384, 23.70362, 23.91331, 24.1229, 
    24.33238, 24.54175, 24.75102, 24.96016, 25.16919, 25.3781, 25.58688, 
    25.79553, 26.00405, 26.21243, 26.42067, 26.62877, 26.83673, 27.04453, 
    27.25219, 27.45968, 27.66702, 27.8742, 28.08121, 28.28805, 28.49472, 
    28.70122, 28.90754, 29.11368, 29.31963, 29.5254, 29.73097, 29.93635, 
    30.14154, 30.34653, 30.55131, 30.75589, 30.96026, 31.16442, 31.36837, 
    31.5721, 31.77561, 31.9789, 32.18196, 32.38479, 32.58739, 32.78976, 
    32.9919, 33.1938, 33.39545, 33.59686, 33.79803, 33.99894, 34.19961, 
    34.40002, 34.60017, 34.80006, 34.9997, 35.19907, 35.39817, 35.59701, 
    35.79557, 35.99386, 36.19188, 36.38961, 36.58707, 36.78425, 36.98114, 
    37.17775, 37.37407, 37.5701, 37.76583, 37.96127, 38.15642, 38.35126, 
    38.54581, 38.74005, 38.93399, 39.12762, 39.32095, 39.51397, 39.70667, 
    39.89907, 40.09114, 40.28291, 40.47435, 40.66547, 40.85627, 41.04675, 
    41.2369, 41.42673, 41.61623, 41.80541, 41.99425, 42.18276, 42.37094, 
    42.55878, 42.74629, 42.93346, 43.12029, 43.30678, 43.49293, 43.67874, 
    43.8642, 44.04932, 44.2341, 44.41853, 44.60261, 44.78635, 44.96973, 
    45.15276, 45.33544, 45.51777, 45.69975, 45.88136, 46.06263, 46.24354, 
    46.42409, 46.60429, 46.78412, 46.9636, 47.14272, 47.32147, 47.49987, 
    47.6779, 47.85557, 48.03288, 48.20982, 48.3864, 48.56261, 48.73846, 
    48.91395, 49.08907, 49.26382, 49.4382, 49.61222, 49.78587, 49.95914, 
    50.13206, 50.3046, 50.47677, 50.64857, 50.82001, 50.99107, 51.16177, 
    51.33209, 51.50204,
  -29.79384, -29.65686, -29.51956, -29.38193, -29.24397, -29.10568, 
    -28.96705, -28.8281, -28.68881, -28.54919, -28.40923, -28.26894, 
    -28.12831, -27.98735, -27.84604, -27.7044, -27.56242, -27.42009, 
    -27.27743, -27.13442, -26.99107, -26.84738, -26.70334, -26.55896, 
    -26.41422, -26.26915, -26.12372, -25.97795, -25.83183, -25.68536, 
    -25.53854, -25.39136, -25.24384, -25.09596, -24.94773, -24.79914, 
    -24.6502, -24.5009, -24.35125, -24.20124, -24.05088, -23.90015, 
    -23.74907, -23.59763, -23.44583, -23.29366, -23.14114, -22.98826, 
    -22.83501, -22.6814, -22.52743, -22.37309, -22.21839, -22.06333, 
    -21.9079, -21.7521, -21.59594, -21.43941, -21.28251, -21.12525, 
    -20.96762, -20.80962, -20.65125, -20.49251, -20.3334, -20.17393, 
    -20.01408, -19.85386, -19.69327, -19.53231, -19.37098, -19.20928, 
    -19.0472, -18.88476, -18.72194, -18.55875, -18.39518, -18.23125, 
    -18.06694, -17.90225, -17.7372, -17.57177, -17.40596, -17.23979, 
    -17.07324, -16.90631, -16.73901, -16.57134, -16.4033, -16.23488, 
    -16.06609, -15.89692, -15.72738, -15.55747, -15.38718, -15.21652, 
    -15.04549, -14.87408, -14.70231, -14.53016, -14.35764, -14.18474, 
    -14.01148, -13.83784, -13.66384, -13.48946, -13.31471, -13.1396, 
    -12.96411, -12.78826, -12.61203, -12.43544, -12.25848, -12.08116, 
    -11.90347, -11.72541, -11.54699, -11.3682, -11.18905, -11.00953, 
    -10.82966, -10.64942, -10.46882, -10.28786, -10.10654, -9.924862, 
    -9.742826, -9.560434, -9.377686, -9.194581, -9.011123, -8.827312, 
    -8.643148, -8.458633, -8.273767, -8.088553, -7.902991, -7.717082, 
    -7.530827, -7.344227, -7.157284, -6.969999, -6.782373, -6.594407, 
    -6.406103, -6.217462, -6.028485, -5.839174, -5.64953, -5.459555, 
    -5.26925, -5.078617, -4.887656, -4.696371, -4.504761, -4.312829, 
    -4.120577, -3.928006, -3.735118, -3.541915, -3.348398, -3.154569, 
    -2.96043, -2.765982, -2.571229, -2.37617, -2.18081, -1.985148, -1.789188, 
    -1.592931, -1.39638, -1.199536, -1.002402, -0.804979, -0.60727, 
    -0.4092769, -0.211002, -0.01244745, 0.1863845, 0.3854915, 0.5848714, 
    0.7845218, 0.9844402, 1.184624, 1.385072, 1.58578, 1.786747, 1.98797, 
    2.189446, 2.391173, 2.593148, 2.795369, 2.997833, 3.200537, 3.403479, 
    3.606656, 3.810065, 4.013704, 4.21757, 4.421659, 4.62597, 4.830499, 
    5.035244, 5.240201, 5.445367, 5.65074, 5.856317, 6.062095, 6.26807, 
    6.47424, 6.680602, 6.887152, 7.093887, 7.300805, 7.507902, 7.715175, 
    7.922621, 8.130236, 8.338017, 8.545963, 8.754067, 8.962329, 9.170744, 
    9.379309, 9.58802, 9.796875, 10.00587, 10.215, 10.42427, 10.63366, 
    10.84318, 11.05282, 11.26259, 11.47247, 11.68246, 11.89256, 12.10276, 
    12.31307, 12.52348, 12.73398, 12.94457, 13.15525, 13.36602, 13.57686, 
    13.78778, 13.99878, 14.20984, 14.42097, 14.63216, 14.84342, 15.05472, 
    15.26608, 15.47749, 15.68894, 15.90043, 16.11196, 16.32351, 16.5351, 
    16.74672, 16.95836, 17.17001, 17.38168, 17.59336, 17.80505, 18.01674, 
    18.22843, 18.44012, 18.6518, 18.86347, 19.07512, 19.28675, 19.49837, 
    19.70995, 19.92151, 20.13303, 20.34451, 20.55596, 20.76735, 20.97871, 
    21.19, 21.40125, 21.61243, 21.82355, 22.0346, 22.24559, 22.4565, 
    22.66733, 22.87808, 23.08875, 23.29932, 23.50981, 23.7202, 23.93049, 
    24.14068, 24.35077, 24.56074, 24.7706, 24.98034, 25.18997, 25.39947, 
    25.60884, 25.81809, 26.0272, 26.23617, 26.445, 26.65369, 26.86223, 
    27.07063, 27.27886, 27.48694, 27.69486, 27.90262, 28.1102, 28.31762, 
    28.52487, 28.73194, 28.93883, 29.14553, 29.35205, 29.55839, 29.76452, 
    29.97047, 30.17622, 30.38176, 30.5871, 30.79223, 30.99716, 31.20187, 
    31.40636, 31.61064, 31.81469, 32.01852, 32.22213, 32.4255, 32.62864, 
    32.83154, 33.03421, 33.23664, 33.43882, 33.64075, 33.84244, 34.04388, 
    34.24506, 34.44598, 34.64665, 34.84706, 35.0472, 35.24708, 35.44669, 
    35.64602, 35.84509, 36.04387, 36.24239, 36.44062, 36.63857, 36.83623, 
    37.0336, 37.23069, 37.42749, 37.624, 37.82021, 38.01612, 38.21173, 
    38.40705, 38.60205, 38.79676, 38.99116, 39.18525, 39.37903, 39.5725, 
    39.76565, 39.95849, 40.15101, 40.34321, 40.53509, 40.72665, 40.91788, 
    41.1088, 41.29937, 41.48963, 41.67955, 41.86914, 42.0584, 42.24733, 
    42.43591, 42.62416, 42.81208, 42.99965, 43.18688, 43.37377, 43.56031, 
    43.74651, 43.93237, 44.11787, 44.30303, 44.48784, 44.6723, 44.85641, 
    45.04016, 45.22357, 45.40662, 45.58931, 45.77164, 45.95362, 46.13525, 
    46.31651, 46.49741, 46.67795, 46.85814, 47.03795, 47.21741, 47.3965, 
    47.57523, 47.7536, 47.9316, 48.10923, 48.2865, 48.4634, 48.63993, 
    48.8161, 48.99189, 49.16732, 49.34238, 49.51707, 49.69139, 49.86533, 
    50.03891, 50.21212, 50.38495, 50.55742, 50.7295, 50.90122, 51.07257, 
    51.24354, 51.41414, 51.58437,
  -29.89238, -29.75532, -29.61793, -29.48021, -29.34216, -29.20378, 
    -29.06506, -28.92601, -28.78663, -28.64691, -28.50685, -28.36646, 
    -28.22573, -28.08466, -27.94325, -27.8015, -27.6594, -27.51697, 
    -27.37419, -27.23107, -27.0876, -26.94379, -26.79963, -26.65513, 
    -26.51028, -26.36508, -26.21953, -26.07363, -25.92737, -25.78077, 
    -25.63381, -25.48651, -25.33884, -25.19083, -25.04245, -24.89372, 
    -24.74464, -24.5952, -24.4454, -24.29524, -24.14472, -23.99384, -23.8426, 
    -23.691, -23.53904, -23.38672, -23.23403, -23.08098, -22.92756, 
    -22.77378, -22.61964, -22.46513, -22.31025, -22.15501, -21.9994, 
    -21.84342, -21.68707, -21.53036, -21.37327, -21.21581, -21.05799, 
    -20.89979, -20.74123, -20.58229, -20.42298, -20.2633, -20.10324, 
    -19.94282, -19.78202, -19.62084, -19.4593, -19.29738, -19.13508, 
    -18.97241, -18.80937, -18.64595, -18.48215, -18.31799, -18.15344, 
    -17.98852, -17.82322, -17.65755, -17.4915, -17.32508, -17.15828, 
    -16.9911, -16.82355, -16.65562, -16.48732, -16.31864, -16.14958, 
    -15.98015, -15.81034, -15.64015, -15.46959, -15.29866, -15.12734, 
    -14.95566, -14.7836, -14.61116, -14.43835, -14.26516, -14.0916, 
    -13.91767, -13.74336, -13.56868, -13.39363, -13.2182, -13.0424, 
    -12.86624, -12.6897, -12.51279, -12.33551, -12.15786, -11.97984, 
    -11.80145, -11.62269, -11.44357, -11.26408, -11.08423, -10.90401, 
    -10.72342, -10.54247, -10.36116, -10.17949, -9.997452, -9.815056, 
    -9.6323, -9.449185, -9.265713, -9.081883, -8.897698, -8.713158, 
    -8.528263, -8.343016, -8.157416, -7.971466, -7.785166, -7.598518, 
    -7.411522, -7.22418, -7.036493, -6.848463, -6.660089, -6.471375, 
    -6.282322, -6.092929, -5.9032, -5.713136, -5.522737, -5.332005, 
    -5.140943, -4.94955, -4.75783, -4.565783, -4.373411, -4.180717, -3.9877, 
    -3.794364, -3.60071, -3.406739, -3.212454, -3.017856, -2.822947, 
    -2.627729, -2.432204, -2.236374, -2.040241, -1.843806, -1.647072, 
    -1.450041, -1.252715, -1.055096, -0.8571854, -0.6589864, -0.460501, 
    -0.2617311, -0.0626791, 0.1366528, 0.3362622, 0.5361468, 0.7363044, 
    0.9367325, 1.137429, 1.338391, 1.539616, 1.741102, 1.942846, 2.144845, 
    2.347099, 2.549602, 2.752353, 2.95535, 3.158589, 3.362068, 3.565785, 
    3.769736, 3.973918, 4.178329, 4.382967, 4.587828, 4.792909, 4.998207, 
    5.20372, 5.409444, 5.615377, 5.821516, 6.027857, 6.234398, 6.441135, 
    6.648066, 6.855186, 7.062495, 7.269987, 7.47766, 7.685511, 7.893536, 
    8.101732, 8.310097, 8.518626, 8.727317, 8.936166, 9.145169, 9.354324, 
    9.563627, 9.773075, 9.982664, 10.19239, 10.40225, 10.61224, 10.82236, 
    11.03261, 11.24297, 11.45346, 11.66405, 11.87476, 12.08557, 12.29648, 
    12.5075, 12.71861, 12.92981, 13.1411, 13.35248, 13.56393, 13.77547, 
    13.98708, 14.19875, 14.4105, 14.62231, 14.83418, 15.0461, 15.25808, 
    15.4701, 15.68217, 15.89428, 16.10642, 16.3186, 16.53081, 16.74305, 
    16.95531, 17.16758, 17.37987, 17.59217, 17.80448, 18.01679, 18.2291, 
    18.44141, 18.65371, 18.866, 19.07827, 19.29053, 19.50276, 19.71496, 
    19.92714, 20.13928, 20.35138, 20.56344, 20.77546, 20.98743, 21.19934, 
    21.4112, 21.623, 21.83473, 22.0464, 22.258, 22.46952, 22.68097, 22.89233, 
    23.10361, 23.31479, 23.52589, 23.73689, 23.94779, 24.15858, 24.36927, 
    24.57985, 24.79031, 25.00066, 25.21088, 25.42098, 25.63095, 25.84079, 
    26.0505, 26.26007, 26.46949, 26.67877, 26.8879, 27.09688, 27.30571, 
    27.51437, 27.72287, 27.93121, 28.13938, 28.34738, 28.5552, 28.76285, 
    28.97031, 29.17759, 29.38468, 29.59158, 29.79829, 30.0048, 30.21111, 
    30.41721, 30.62311, 30.8288, 31.03428, 31.23955, 31.44459, 31.64942, 
    31.85402, 32.0584, 32.26254, 32.46645, 32.67014, 32.87358, 33.07678, 
    33.27974, 33.48245, 33.68491, 33.88712, 34.08908, 34.29079, 34.49223, 
    34.69342, 34.89434, 35.09499, 35.29538, 35.49549, 35.69533, 35.8949, 
    36.09418, 36.29319, 36.49192, 36.69036, 36.88851, 37.08638, 37.28395, 
    37.48123, 37.67821, 37.8749, 38.07129, 38.26737, 38.46315, 38.65863, 
    38.8538, 39.04866, 39.24321, 39.43744, 39.63136, 39.82497, 40.01825, 
    40.21122, 40.40386, 40.59618, 40.78818, 40.97985, 41.17119, 41.3622, 
    41.55288, 41.74322, 41.93324, 42.12291, 42.31225, 42.50125, 42.68991, 
    42.87823, 43.0662, 43.25384, 43.44112, 43.62807, 43.81466, 44.0009, 
    44.1868, 44.37234, 44.55753, 44.74237, 44.92686, 45.11098, 45.29476, 
    45.47818, 45.66123, 45.84393, 46.02627, 46.20825, 46.38987, 46.57112, 
    46.75201, 46.93254, 47.1127, 47.2925, 47.47193, 47.65099, 47.82969, 
    48.00802, 48.18598, 48.36357, 48.54079, 48.71765, 48.89413, 49.07024, 
    49.24598, 49.42134, 49.59634, 49.77096, 49.94521, 50.11908, 50.29258, 
    50.46571, 50.63846, 50.81084, 50.98284, 51.15447, 51.32572, 51.4966, 
    51.6671,
  -29.99129, -29.85415, -29.71667, -29.57886, -29.44072, -29.30225, 
    -29.16344, -29.02429, -28.88482, -28.745, -28.60484, -28.46435, 
    -28.32351, -28.18234, -28.04082, -27.89897, -27.75677, -27.61422, 
    -27.47133, -27.3281, -27.18452, -27.04059, -26.89631, -26.75169, 
    -26.60671, -26.46139, -26.31571, -26.16969, -26.0233, -25.87657, 
    -25.72948, -25.58204, -25.43424, -25.28608, -25.13757, -24.9887, 
    -24.83947, -24.68988, -24.53994, -24.38963, -24.23896, -24.08792, 
    -23.93653, -23.78477, -23.63265, -23.48017, -23.32732, -23.1741, 
    -23.02052, -22.86657, -22.71225, -22.55757, -22.40252, -22.24709, 
    -22.0913, -21.93514, -21.77861, -21.62171, -21.46443, -21.30679, 
    -21.14877, -20.99038, -20.83161, -20.67247, -20.51296, -20.35308, 
    -20.19282, -20.03218, -19.87117, -19.70978, -19.54802, -19.38588, 
    -19.22337, -19.06047, -18.8972, -18.73356, -18.56953, -18.40513, 
    -18.24035, -18.0752, -17.90966, -17.74374, -17.57745, -17.41078, 
    -17.24373, -17.0763, -16.9085, -16.74031, -16.57175, -16.4028, -16.23348, 
    -16.06378, -15.8937, -15.72325, -15.55241, -15.3812, -15.20961, 
    -15.03764, -14.86529, -14.69256, -14.51946, -14.34598, -14.17213, 
    -13.9979, -13.82329, -13.6483, -13.47294, -13.29721, -13.1211, -12.94462, 
    -12.76776, -12.59053, -12.41293, -12.23495, -12.0566, -11.87789, 
    -11.6988, -11.51934, -11.33951, -11.15931, -10.97875, -10.79782, 
    -10.61652, -10.43485, -10.25282, -10.07043, -9.887673, -9.704554, 
    -9.521072, -9.33723, -9.153028, -8.968468, -8.783549, -8.598274, 
    -8.412643, -8.226658, -8.040318, -7.853626, -7.666583, -7.47919, 
    -7.291448, -7.103358, -6.914921, -6.72614, -6.537014, -6.347546, 
    -6.157737, -5.967587, -5.7771, -5.586276, -5.395116, -5.203623, 
    -5.011797, -4.81964, -4.627154, -4.43434, -4.241201, -4.047738, 
    -3.853951, -3.659844, -3.465418, -3.270675, -3.075616, -2.880244, 
    -2.68456, -2.488566, -2.292264, -2.095657, -1.898745, -1.701532, 
    -1.504019, -1.306208, -1.108102, -0.9097018, -0.7110106, -0.5120302, 
    -0.3127629, -0.1132111, 0.08662318, 0.2867375, 0.4871295, 0.6877969, 
    0.8887372, 1.089948, 1.291427, 1.493172, 1.695179, 1.897448, 2.099974, 
    2.302756, 2.50579, 2.709075, 2.912607, 3.116385, 3.320404, 3.524663, 
    3.729158, 3.933887, 4.138847, 4.344036, 4.549449, 4.755085, 4.96094, 
    5.167012, 5.373298, 5.579794, 5.786497, 5.993405, 6.200515, 6.407823, 
    6.615326, 6.823021, 7.030905, 7.238976, 7.447228, 7.65566, 7.864268, 
    8.07305, 8.282, 8.491117, 8.700397, 8.909836, 9.119431, 9.329181, 
    9.539079, 9.749124, 9.959311, 10.16964, 10.3801, 10.59069, 10.80142, 
    11.01226, 11.22324, 11.43432, 11.64553, 11.85684, 12.06826, 12.27979, 
    12.49141, 12.70314, 12.91495, 13.12686, 13.33885, 13.55092, 13.76307, 
    13.9753, 14.1876, 14.39996, 14.61239, 14.82488, 15.03742, 15.25002, 
    15.46266, 15.67535, 15.88809, 16.10085, 16.31366, 16.52649, 16.73935, 
    16.95223, 17.16513, 17.37805, 17.59097, 17.80391, 18.01684, 18.22978, 
    18.44271, 18.65563, 18.86855, 19.08144, 19.29432, 19.50718, 19.72001, 
    19.9328, 20.14557, 20.35829, 20.57098, 20.78361, 20.9962, 21.20874, 
    21.42122, 21.63364, 21.84599, 22.05828, 22.27049, 22.48263, 22.69469, 
    22.90667, 23.11856, 23.33036, 23.54207, 23.75368, 23.96519, 24.17659, 
    24.38789, 24.59908, 24.81014, 25.0211, 25.23193, 25.44263, 25.6532, 
    25.86364, 26.07395, 26.28411, 26.49413, 26.70401, 26.91373, 27.1233, 
    27.33272, 27.54197, 27.75106, 27.95999, 28.16874, 28.37732, 28.58573, 
    28.79395, 29.00199, 29.20984, 29.41751, 29.62498, 29.83226, 30.03934, 
    30.24621, 30.45288, 30.65935, 30.8656, 31.07164, 31.27746, 31.48306, 
    31.68844, 31.89359, 32.09851, 32.3032, 32.50766, 32.71188, 32.91587, 
    33.11961, 33.3231, 33.52634, 33.72934, 33.93208, 34.13456, 34.33679, 
    34.53876, 34.74046, 34.9419, 35.14307, 35.34396, 35.54459, 35.74493, 
    35.94501, 36.14479, 36.3443, 36.54353, 36.74246, 36.9411, 37.13946, 
    37.33752, 37.53528, 37.73275, 37.92991, 38.12678, 38.32334, 38.51959, 
    38.71553, 38.91117, 39.10649, 39.3015, 39.49619, 39.69057, 39.88463, 
    40.07836, 40.27177, 40.46486, 40.65762, 40.85006, 41.04216, 41.23394, 
    41.42538, 41.61648, 41.80725, 41.99769, 42.18778, 42.37754, 42.56695, 
    42.75602, 42.94475, 43.13313, 43.32117, 43.50885, 43.69619, 43.88318, 
    44.06982, 44.2561, 44.44203, 44.62761, 44.81282, 44.99768, 45.18219, 
    45.36633, 45.55012, 45.73354, 45.91661, 46.0993, 46.28164, 46.46362, 
    46.64522, 46.82646, 47.00734, 47.18784, 47.36798, 47.54775, 47.72715, 
    47.90618, 48.08484, 48.26313, 48.44105, 48.61859, 48.79576, 48.97256, 
    49.14898, 49.32504, 49.50071, 49.67601, 49.85093, 50.02548, 50.19965, 
    50.37345, 50.54687, 50.71991, 50.89258, 51.06487, 51.23677, 51.40831, 
    51.57946, 51.75024,
  -30.09057, -29.95334, -29.81578, -29.67788, -29.53965, -29.40109, 
    -29.26219, -29.12295, -28.98337, -28.84346, -28.70321, -28.56261, 
    -28.42168, -28.2804, -28.13878, -27.99682, -27.85451, -27.71186, 
    -27.56886, -27.42551, -27.28181, -27.13777, -26.99338, -26.84863, 
    -26.70354, -26.55809, -26.41229, -26.26613, -26.11962, -25.97276, 
    -25.82554, -25.67796, -25.53003, -25.38173, -25.23308, -25.08407, 
    -24.9347, -24.78497, -24.63487, -24.48441, -24.33359, -24.18241, 
    -24.03086, -23.87894, -23.72666, -23.57402, -23.421, -23.26762, 
    -23.11387, -22.95975, -22.80527, -22.65041, -22.49518, -22.33958, 
    -22.18361, -22.02727, -21.87055, -21.71346, -21.556, -21.39816, 
    -21.23995, -21.08137, -20.92241, -20.76307, -20.60336, -20.44327, 
    -20.2828, -20.12195, -19.96073, -19.79913, -19.63715, -19.4748, 
    -19.31206, -19.14895, -18.98545, -18.82158, -18.65732, -18.49269, 
    -18.32767, -18.16228, -17.99651, -17.83035, -17.66381, -17.49689, 
    -17.3296, -17.16191, -16.99385, -16.82541, -16.65659, -16.48738, 
    -16.3178, -16.14783, -15.97748, -15.80675, -15.63564, -15.46415, 
    -15.29228, -15.12003, -14.94739, -14.77438, -14.60099, -14.42721, 
    -14.25306, -14.07853, -13.90362, -13.72833, -13.55267, -13.37662, 
    -13.2002, -13.0234, -12.84623, -12.66868, -12.49075, -12.31245, 
    -12.13378, -11.95473, -11.7753, -11.59551, -11.41534, -11.2348, 
    -11.05389, -10.87261, -10.69096, -10.50894, -10.32655, -10.1438, 
    -9.960682, -9.777197, -9.593349, -9.409136, -9.224561, -9.039623, 
    -8.854326, -8.668669, -8.482654, -8.29628, -8.10955, -7.922465, 
    -7.735026, -7.547234, -7.35909, -7.170596, -6.981752, -6.79256, 
    -6.603022, -6.413137, -6.22291, -6.03234, -5.841428, -5.650177, 
    -5.458587, -5.266661, -5.0744, -4.881805, -4.688878, -4.495621, 
    -4.302035, -4.108122, -3.913884, -3.719322, -3.524439, -3.329235, 
    -3.133714, -2.937876, -2.741724, -2.545259, -2.348483, -2.1514, 
    -1.954009, -1.756314, -1.558317, -1.360019, -1.161423, -0.9625312, 
    -0.7633452, -0.5638676, -0.3641006, -0.1640463, 0.0362928, 0.2369145, 
    0.4378164, 0.6389962, 0.8404514, 1.04218, 1.244178, 1.446445, 1.648977, 
    1.851773, 2.054828, 2.258142, 2.46171, 2.665531, 2.869602, 3.07392, 
    3.278483, 3.483287, 3.688329, 3.893608, 4.09912, 4.304862, 4.510832, 
    4.717026, 4.923442, 5.130076, 5.336926, 5.543988, 5.75126, 5.958738, 
    6.16642, 6.374301, 6.58238, 6.790653, 6.999117, 7.207768, 7.416604, 
    7.62562, 7.834815, 8.044184, 8.253724, 8.463432, 8.673306, 8.883339, 
    9.093531, 9.303877, 9.514374, 9.725019, 9.935807, 10.14674, 10.3578, 
    10.569, 10.78033, 10.99179, 11.20337, 11.41507, 11.62688, 11.83881, 
    12.05085, 12.26299, 12.47523, 12.68757, 12.9, 13.11252, 13.32513, 
    13.53783, 13.7506, 13.96345, 14.17637, 14.38935, 14.60241, 14.81552, 
    15.02869, 15.24191, 15.45518, 15.6685, 15.88186, 16.09525, 16.30868, 
    16.52214, 16.73563, 16.94914, 17.16267, 17.37621, 17.58976, 17.80333, 
    18.01689, 18.23046, 18.44402, 18.65757, 18.87111, 19.08464, 19.29814, 
    19.51163, 19.72508, 19.93851, 20.1519, 20.36525, 20.57856, 20.79182, 
    21.00504, 21.2182, 21.4313, 21.64434, 21.85732, 22.07023, 22.28306, 
    22.49582, 22.7085, 22.9211, 23.13361, 23.34603, 23.55835, 23.77058, 
    23.9827, 24.19472, 24.40663, 24.61843, 24.83011, 25.04167, 25.2531, 
    25.46441, 25.67559, 25.88664, 26.09755, 26.30831, 26.51893, 26.72941, 
    26.93973, 27.14989, 27.3599, 27.56975, 27.77943, 27.98895, 28.19829, 
    28.40745, 28.61644, 28.82525, 29.03387, 29.2423, 29.45055, 29.6586, 
    29.86645, 30.07409, 30.28154, 30.48878, 30.69581, 30.90262, 31.10922, 
    31.31561, 31.52176, 31.7277, 31.9334, 32.13888, 32.34412, 32.54913, 
    32.75389, 32.95842, 33.16269, 33.36673, 33.57051, 33.77404, 33.97731, 
    34.18032, 34.38308, 34.58557, 34.78779, 34.98975, 35.19143, 35.39285, 
    35.59398, 35.79484, 35.99541, 36.19571, 36.39572, 36.59544, 36.79487, 
    36.99401, 37.19286, 37.39141, 37.58966, 37.78761, 37.98525, 38.18259, 
    38.37963, 38.57636, 38.77277, 38.96888, 39.16466, 39.36013, 39.55529, 
    39.75012, 39.94463, 40.13882, 40.33268, 40.52621, 40.71942, 40.91229, 
    41.10484, 41.29704, 41.48891, 41.68045, 41.87165, 42.06251, 42.25303, 
    42.4432, 42.63303, 42.82251, 43.01165, 43.20044, 43.38887, 43.57696, 
    43.7647, 43.95208, 44.13911, 44.32579, 44.5121, 44.69806, 44.88366, 
    45.0689, 45.25378, 45.4383, 45.62246, 45.80625, 45.98967, 46.17273, 
    46.35543, 46.53776, 46.71972, 46.90131, 47.08253, 47.26338, 47.44386, 
    47.62397, 47.80371, 47.98307, 48.16206, 48.34068, 48.51892, 48.69679, 
    48.87428, 49.0514, 49.22813, 49.4045, 49.58048, 49.75609, 49.93132, 
    50.10617, 50.28064, 50.45473, 50.62844, 50.80177, 50.97473, 51.1473, 
    51.31949, 51.4913, 51.66273, 51.83378,
  -30.19021, -30.0529, -29.91525, -29.77727, -29.63895, -29.5003, -29.36131, 
    -29.22198, -29.08231, -28.9423, -28.80195, -28.66126, -28.52022, 
    -28.37885, -28.23712, -28.09505, -27.95264, -27.80988, -27.66677, 
    -27.52331, -27.3795, -27.23534, -27.09083, -26.94596, -26.80075, 
    -26.65518, -26.50925, -26.36297, -26.21634, -26.06934, -25.92199, 
    -25.77428, -25.62621, -25.47778, -25.32899, -25.17984, -25.03032, 
    -24.88045, -24.7302, -24.5796, -24.42863, -24.27729, -24.12559, 
    -23.97352, -23.82108, -23.66827, -23.51509, -23.36155, -23.20763, 
    -23.05334, -22.89869, -22.74366, -22.58825, -22.43248, -22.27633, 
    -22.1198, -21.9629, -21.80563, -21.64798, -21.48995, -21.33155, 
    -21.17277, -21.01361, -20.85407, -20.69416, -20.53386, -20.37319, 
    -20.21214, -20.05071, -19.8889, -19.7267, -19.56413, -19.40117, 
    -19.23783, -19.07411, -18.91001, -18.74553, -18.58066, -18.41541, 
    -18.24978, -18.08377, -17.91737, -17.75059, -17.58342, -17.41587, 
    -17.24794, -17.07963, -16.91093, -16.74184, -16.57238, -16.40252, 
    -16.23229, -16.06167, -15.89067, -15.71929, -15.54752, -15.37536, 
    -15.20283, -15.02991, -14.85661, -14.68292, -14.50886, -14.33441, 
    -14.15958, -13.98437, -13.80877, -13.6328, -13.45645, -13.27971, 
    -13.1026, -12.92511, -12.74723, -12.56898, -12.39036, -12.21135, 
    -12.03197, -11.85221, -11.67208, -11.49157, -11.31069, -11.12943, 
    -10.9478, -10.7658, -10.58343, -10.40068, -10.21757, -10.03409, 
    -9.850235, -9.666018, -9.481433, -9.296483, -9.111169, -8.925491, 
    -8.739451, -8.55305, -8.366287, -8.179166, -7.991687, -7.80385, 
    -7.615658, -7.427111, -7.238211, -7.048958, -6.859354, -6.669402, 
    -6.479101, -6.288453, -6.097459, -5.906122, -5.714442, -5.522421, 
    -5.330061, -5.137362, -4.944328, -4.750958, -4.557255, -4.363221, 
    -4.168857, -3.974165, -3.779147, -3.583804, -3.388138, -3.192152, 
    -2.995846, -2.799224, -2.602286, -2.405035, -2.207472, -2.009601, 
    -1.811422, -1.612938, -1.414151, -1.215063, -1.015677, -0.8159937, 
    -0.6160164, -0.4157471, -0.215188, -0.0143414, 0.1867903, 0.3882047, 
    0.5898995, 0.7918722, 0.9941204, 1.196642, 1.399433, 1.602493, 1.805818, 
    2.009406, 2.213253, 2.417359, 2.621719, 2.826332, 3.031193, 3.236302, 
    3.441654, 3.647248, 3.853079, 4.059146, 4.265445, 4.471974, 4.67873, 
    4.885708, 5.092908, 5.300325, 5.507957, 5.715801, 5.923852, 6.13211, 
    6.340569, 6.549227, 6.758081, 6.967127, 7.176363, 7.385786, 7.59539, 
    7.805175, 8.015136, 8.225269, 8.435572, 8.646041, 8.856673, 9.067465, 
    9.278412, 9.489511, 9.70076, 9.912154, 10.12369, 10.33536, 10.54717, 
    10.75911, 10.97118, 11.18338, 11.39569, 11.60812, 11.82066, 12.03332, 
    12.24607, 12.45894, 12.6719, 12.88495, 13.0981, 13.31133, 13.52465, 
    13.73804, 13.95152, 14.16506, 14.37868, 14.59236, 14.8061, 15.0199, 
    15.23375, 15.44765, 15.6616, 15.87558, 16.08961, 16.30367, 16.51777, 
    16.73188, 16.94603, 17.16019, 17.37436, 17.58855, 17.80274, 18.01694, 
    18.23114, 18.44533, 18.65952, 18.87369, 19.08785, 19.30199, 19.5161, 
    19.73019, 19.94425, 20.15827, 20.37225, 20.58619, 20.80008, 21.01393, 
    21.22772, 21.44145, 21.65512, 21.86872, 22.08225, 22.29572, 22.5091, 
    22.72241, 22.93563, 23.14876, 23.3618, 23.57474, 23.78759, 24.00033, 
    24.21297, 24.42549, 24.6379, 24.8502, 25.06237, 25.27442, 25.48634, 
    25.69813, 25.90978, 26.12129, 26.33267, 26.54389, 26.75497, 26.96589, 
    27.17666, 27.38726, 27.59771, 27.80798, 28.01809, 28.22802, 28.43778, 
    28.64735, 28.85675, 29.06595, 29.27497, 29.48379, 29.69242, 29.90085, 
    30.10907, 30.31709, 30.5249, 30.7325, 30.93988, 31.14705, 31.35399, 
    31.56071, 31.7672, 31.97347, 32.1795, 32.38529, 32.59085, 32.79616, 
    33.00123, 33.20605, 33.41063, 33.61494, 33.81901, 34.02282, 34.22636, 
    34.42965, 34.63266, 34.83541, 35.03789, 35.24009, 35.44202, 35.64367, 
    35.84504, 36.04613, 36.24693, 36.44744, 36.64767, 36.8476, 37.04724, 
    37.24657, 37.44562, 37.64436, 37.84279, 38.04092, 38.23874, 38.43626, 
    38.63346, 38.83035, 39.02692, 39.22318, 39.41911, 39.61473, 39.81002, 
    40.00499, 40.19962, 40.39394, 40.58792, 40.78157, 40.97488, 41.16787, 
    41.36051, 41.55282, 41.74479, 41.93641, 42.12769, 42.31863, 42.50923, 
    42.69947, 42.88937, 43.07892, 43.26812, 43.45696, 43.64545, 43.83359, 
    44.02137, 44.20879, 44.39585, 44.58256, 44.76891, 44.95489, 45.14051, 
    45.32576, 45.51065, 45.69518, 45.87934, 46.06313, 46.24656, 46.42962, 
    46.6123, 46.79461, 46.97655, 47.15813, 47.33932, 47.52015, 47.7006, 
    47.88067, 48.06037, 48.23969, 48.41864, 48.59721, 48.77539, 48.95321, 
    49.13064, 49.30769, 49.48437, 49.66066, 49.83658, 50.01211, 50.18726, 
    50.36203, 50.53642, 50.71042, 50.88405, 51.05729, 51.23014, 51.40262, 
    51.57471, 51.74642, 51.91775,
  -30.29023, -30.15283, -30.0151, -29.87703, -29.73863, -29.59989, -29.4608, 
    -29.32138, -29.18162, -29.04152, -28.90107, -28.76028, -28.61915, 
    -28.47767, -28.33584, -28.19367, -28.05115, -27.90828, -27.76506, 
    -27.62149, -27.47757, -27.33329, -27.18867, -27.04369, -26.89835, 
    -26.75266, -26.60661, -26.4602, -26.31344, -26.16632, -26.01884, 
    -25.87099, -25.72279, -25.57422, -25.42529, -25.276, -25.12635, 
    -24.97632, -24.82594, -24.67518, -24.52406, -24.37258, -24.22072, 
    -24.06849, -23.9159, -23.76293, -23.60959, -23.45588, -23.3018, 
    -23.14734, -22.99252, -22.83731, -22.68174, -22.52578, -22.36945, 
    -22.21275, -22.05567, -21.89821, -21.74037, -21.58215, -21.42356, 
    -21.26458, -21.10523, -20.94549, -20.78538, -20.62488, -20.464, 
    -20.30274, -20.1411, -19.97907, -19.81666, -19.65387, -19.4907, 
    -19.32714, -19.16319, -18.99887, -18.83415, -18.66905, -18.50357, 
    -18.3377, -18.17145, -18.00481, -17.83778, -17.67037, -17.50257, 
    -17.33439, -17.16582, -16.99686, -16.82752, -16.65779, -16.48767, 
    -16.31717, -16.14628, -15.97501, -15.80335, -15.6313, -15.45887, 
    -15.28605, -15.11284, -14.93925, -14.76528, -14.59092, -14.41617, 
    -14.24104, -14.06553, -13.88963, -13.71335, -13.53668, -13.35964, 
    -13.18221, -13.00439, -12.8262, -12.64763, -12.46867, -12.28934, 
    -12.10962, -11.92953, -11.74905, -11.5682, -11.38698, -11.20537, 
    -11.02339, -10.84104, -10.65831, -10.47521, -10.29173, -10.10789, 
    -9.923671, -9.739083, -9.554126, -9.368801, -9.183108, -8.997049, 
    -8.810624, -8.623836, -8.436684, -8.249169, -8.061295, -7.873059, 
    -7.684465, -7.495514, -7.306206, -7.116543, -6.926527, -6.736158, 
    -6.545438, -6.354368, -6.162951, -5.971186, -5.779076, -5.586622, 
    -5.393825, -5.200688, -5.007212, -4.813397, -4.619247, -4.424763, 
    -4.229946, -4.034799, -3.839321, -3.643517, -3.447387, -3.250934, 
    -3.054158, -2.857063, -2.65965, -2.461921, -2.263878, -2.065523, 
    -1.866858, -1.667885, -1.468607, -1.269025, -1.069142, -0.8689591, 
    -0.6684796, -0.4677055, -0.266639, -0.06528247, 0.1363617, 0.3382913, 
    0.5405037, 0.7429966, 0.9457675, 1.148814, 1.352133, 1.555723, 1.75958, 
    1.963703, 2.168088, 2.372734, 2.577636, 2.782793, 2.988201, 3.193859, 
    3.399763, 3.60591, 3.812297, 4.018922, 4.225781, 4.432873, 4.640193, 
    4.847738, 5.055507, 5.263495, 5.4717, 5.680118, 5.888746, 6.097582, 
    6.306622, 6.515863, 6.725302, 6.934935, 7.144759, 7.354771, 7.564967, 
    7.775345, 7.985901, 8.196631, 8.407533, 8.618603, 8.829836, 9.041231, 
    9.252783, 9.464489, 9.676345, 9.888349, 10.10049, 10.31278, 10.5252, 
    10.73776, 10.95044, 11.16325, 11.37618, 11.58923, 11.8024, 12.01567, 
    12.22905, 12.44254, 12.65612, 12.8698, 13.08358, 13.29744, 13.51138, 
    13.72541, 13.93951, 14.15369, 14.36793, 14.58224, 14.79662, 15.01105, 
    15.22553, 15.44007, 15.65465, 15.86927, 16.08393, 16.29863, 16.51336, 
    16.72812, 16.94289, 17.15769, 17.3725, 17.58733, 17.80216, 18.01699, 
    18.23183, 18.44666, 18.66148, 18.87629, 19.09108, 19.30586, 19.52061, 
    19.73533, 19.95002, 20.16468, 20.3793, 20.59387, 20.8084, 21.02287, 
    21.2373, 21.45166, 21.66596, 21.8802, 22.09436, 22.30845, 22.52247, 
    22.7364, 22.95024, 23.164, 23.37767, 23.59124, 23.80471, 24.01807, 
    24.23133, 24.44448, 24.65751, 24.87042, 25.08321, 25.29587, 25.50841, 
    25.72081, 25.93307, 26.1452, 26.35718, 26.56901, 26.78069, 26.99222, 
    27.20359, 27.4148, 27.62584, 27.83671, 28.04742, 28.25794, 28.46829, 
    28.67846, 28.88844, 29.09824, 29.30784, 29.51725, 29.72646, 29.93547, 
    30.14427, 30.35287, 30.56125, 30.76942, 30.97737, 31.18511, 31.39262, 
    31.5999, 31.80696, 32.01378, 32.22037, 32.42672, 32.63282, 32.83869, 
    33.04431, 33.24968, 33.45479, 33.65966, 33.86426, 34.0686, 34.27269, 
    34.4765, 34.68005, 34.88332, 35.08633, 35.28905, 35.4915, 35.69367, 
    35.89555, 36.09715, 36.29846, 36.49949, 36.70021, 36.90065, 37.10078, 
    37.30062, 37.50015, 37.69938, 37.8983, 38.09692, 38.29523, 38.49322, 
    38.6909, 38.88826, 39.08531, 39.28203, 39.47843, 39.67451, 39.87027, 
    40.06569, 40.26078, 40.45555, 40.64998, 40.84408, 41.03784, 41.23126, 
    41.42435, 41.61709, 41.80949, 42.00154, 42.19325, 42.38462, 42.57563, 
    42.7663, 42.95661, 43.14657, 43.33617, 43.52542, 43.71432, 43.90286, 
    44.09104, 44.27885, 44.46631, 44.65341, 44.84014, 45.0265, 45.21251, 
    45.39814, 45.58341, 45.76831, 45.95284, 46.13699, 46.32078, 46.5042, 
    46.68724, 46.86991, 47.0522, 47.23413, 47.41567, 47.59684, 47.77763, 
    47.95804, 48.13807, 48.31773, 48.49701, 48.6759, 48.85441, 49.03255, 
    49.2103, 49.38767, 49.56466, 49.74126, 49.91748, 50.09332, 50.26877, 
    50.44384, 50.61852, 50.79282, 50.96674, 51.14027, 51.31341, 51.48617, 
    51.65854, 51.83052, 52.00212,
  -30.39061, -30.25314, -30.11532, -29.97717, -29.83868, -29.69985, 
    -29.56068, -29.42117, -29.28131, -29.14112, -29.00057, -28.85969, 
    -28.71845, -28.57688, -28.43495, -28.29267, -28.15005, -28.00707, 
    -27.86374, -27.72006, -27.57603, -27.43164, -27.2869, -27.1418, 
    -26.99635, -26.85053, -26.70436, -26.55783, -26.41094, -26.26369, 
    -26.11608, -25.96811, -25.81977, -25.67107, -25.522, -25.37257, 
    -25.22277, -25.07261, -24.92208, -24.77118, -24.61991, -24.46827, 
    -24.31626, -24.16388, -24.01112, -23.858, -23.7045, -23.55062, -23.39638, 
    -23.24175, -23.08676, -22.93138, -22.77563, -22.6195, -22.463, -22.30611, 
    -22.14884, -21.9912, -21.83318, -21.67477, -21.51598, -21.35681, 
    -21.19726, -21.03733, -20.87701, -20.71631, -20.55523, -20.39376, 
    -20.23191, -20.06967, -19.90705, -19.74404, -19.58064, -19.41686, 
    -19.25269, -19.08814, -18.92319, -18.75787, -18.59215, -18.42604, 
    -18.25955, -18.09267, -17.9254, -17.75774, -17.58969, -17.42126, 
    -17.25243, -17.08322, -16.91361, -16.74362, -16.57324, -16.40247, 
    -16.23131, -16.05976, -15.88783, -15.7155, -15.54279, -15.36969, 
    -15.19619, -15.02232, -14.84805, -14.67339, -14.49835, -14.32292, 
    -14.1471, -13.9709, -13.79431, -13.61734, -13.43997, -13.26223, -13.0841, 
    -12.90558, -12.72668, -12.5474, -12.36773, -12.18768, -12.00725, 
    -11.82644, -11.64525, -11.46368, -11.28173, -11.0994, -10.91669, 
    -10.7336, -10.55014, -10.36631, -10.18209, -9.997508, -9.812549, 
    -9.627218, -9.441516, -9.255444, -9.069002, -8.882193, -8.695015, 
    -8.507472, -8.319564, -8.131291, -7.942656, -7.753659, -7.564302, 
    -7.374586, -7.184511, -6.99408, -6.803294, -6.612154, -6.420661, 
    -6.228817, -6.036623, -5.844081, -5.651192, -5.457958, -5.26438, 
    -5.07046, -4.8762, -4.681601, -4.486664, -4.291392, -4.095787, -3.899849, 
    -3.703582, -3.506986, -3.310063, -3.112816, -2.915246, -2.717356, 
    -2.519146, -2.32062, -2.12178, -1.922626, -1.723162, -1.52339, -1.323312, 
    -1.122929, -0.9222444, -0.7212604, -0.5199789, -0.3184026, -0.1165335, 
    0.08562583, 0.2880731, 0.4908058, 0.6938215, 0.8971178, 1.100692, 
    1.304542, 1.508664, 1.713057, 1.917718, 2.122643, 2.327832, 2.533279, 
    2.738983, 2.944942, 3.151151, 3.357609, 3.564313, 3.771259, 3.978445, 
    4.185868, 4.393525, 4.601413, 4.809529, 5.017869, 5.226431, 5.435212, 
    5.644208, 5.853417, 6.062836, 6.27246, 6.482286, 6.692313, 6.902536, 
    7.112952, 7.323557, 7.534349, 7.745325, 7.956479, 8.16781, 8.379314, 
    8.590987, 8.802826, 9.014828, 9.226989, 9.439304, 9.651772, 9.864388, 
    10.07715, 10.29005, 10.50309, 10.71626, 10.92957, 11.143, 11.35655, 
    11.57023, 11.78401, 11.99791, 12.21192, 12.42603, 12.64025, 12.85456, 
    13.06896, 13.28345, 13.49803, 13.71269, 13.92743, 14.14224, 14.35712, 
    14.57206, 14.78707, 15.00214, 15.21726, 15.43244, 15.64766, 15.86292, 
    16.07822, 16.29356, 16.50893, 16.72432, 16.93974, 17.15518, 17.37063, 
    17.58609, 17.80157, 18.01704, 18.23252, 18.44799, 18.66345, 18.8789, 
    19.09434, 19.30975, 19.52514, 19.74051, 19.95584, 20.17113, 20.38639, 
    20.6016, 20.81677, 21.03188, 21.24694, 21.46194, 21.67688, 21.89175, 
    22.10655, 22.32127, 22.53592, 22.75048, 22.96496, 23.17935, 23.39364, 
    23.60784, 23.82194, 24.03593, 24.24981, 24.46358, 24.67724, 24.89077, 
    25.10418, 25.31746, 25.53062, 25.74364, 25.95652, 26.16925, 26.38185, 
    26.59429, 26.80658, 27.01872, 27.23069, 27.44251, 27.65415, 27.86563, 
    28.07693, 28.28806, 28.49901, 28.70977, 28.92035, 29.13073, 29.34092, 
    29.55092, 29.76071, 29.9703, 30.17969, 30.38886, 30.59783, 30.80657, 
    31.0151, 31.22341, 31.43149, 31.63934, 31.84696, 32.05434, 32.26149, 
    32.4684, 32.67506, 32.88148, 33.08765, 33.29357, 33.49924, 33.70464, 
    33.90979, 34.11467, 34.31929, 34.52364, 34.72772, 34.93153, 35.13506, 
    35.33831, 35.54128, 35.74397, 35.94637, 36.14849, 36.35031, 36.55184, 
    36.75307, 36.95401, 37.15465, 37.35498, 37.55501, 37.75473, 37.95415, 
    38.15326, 38.35204, 38.55052, 38.74868, 38.94652, 39.14404, 39.34124, 
    39.53811, 39.73465, 39.93087, 40.12675, 40.3223, 40.51752, 40.71241, 
    40.90695, 41.10116, 41.29502, 41.48855, 41.68173, 41.87456, 42.06705, 
    42.25919, 42.45097, 42.64241, 42.8335, 43.02423, 43.2146, 43.40462, 
    43.59428, 43.78358, 43.97252, 44.1611, 44.34931, 44.53716, 44.72465, 
    44.91177, 45.09852, 45.2849, 45.47092, 45.65656, 45.84183, 46.02673, 
    46.21126, 46.39541, 46.57919, 46.76259, 46.94561, 47.12826, 47.31053, 
    47.49242, 47.67393, 47.85507, 48.03582, 48.21619, 48.39618, 48.57578, 
    48.755, 48.93385, 49.1123, 49.29037, 49.46806, 49.64536, 49.82227, 
    49.9988, 50.17494, 50.3507, 50.52607, 50.70105, 50.87564, 51.04985, 
    51.22366, 51.39709, 51.57013, 51.74279, 51.91505, 52.08693,
  -30.49137, -30.35382, -30.21592, -30.07768, -29.93911, -29.80019, 
    -29.66093, -29.52133, -29.38139, -29.2411, -29.10046, -28.95948, 
    -28.81815, -28.67647, -28.53444, -28.39206, -28.24933, -28.10625, 
    -27.96281, -27.81903, -27.67488, -27.53038, -27.38552, -27.24031, 
    -27.09474, -26.9488, -26.80251, -26.65586, -26.50884, -26.36147, 
    -26.21373, -26.06562, -25.91715, -25.76831, -25.61911, -25.46954, 
    -25.3196, -25.1693, -25.01862, -24.86757, -24.71616, -24.56437, -24.4122, 
    -24.25967, -24.10676, -23.95347, -23.79982, -23.64578, -23.49137, 
    -23.33658, -23.18141, -23.02587, -22.86994, -22.71364, -22.55695, 
    -22.39989, -22.24244, -22.08461, -21.9264, -21.76781, -21.60883, 
    -21.44946, -21.28972, -21.12959, -20.96907, -20.80817, -20.64688, 
    -20.4852, -20.32314, -20.16069, -19.99785, -19.83463, -19.67101, 
    -19.50701, -19.34262, -19.17784, -19.01266, -18.8471, -18.68115, 
    -18.51481, -18.34808, -18.18095, -18.01344, -17.84553, -17.67723, 
    -17.50855, -17.33947, -17.17, -17.00013, -16.82988, -16.65923, -16.4882, 
    -16.31677, -16.14495, -15.97273, -15.80013, -15.62713, -15.45375, 
    -15.27997, -15.1058, -14.93124, -14.75629, -14.58095, -14.40522, 
    -14.2291, -14.05259, -13.8757, -13.69841, -13.52073, -13.34267, 
    -13.16422, -12.98538, -12.80615, -12.62654, -12.44654, -12.26616, 
    -12.08539, -11.90424, -11.72271, -11.54079, -11.35849, -11.17581, 
    -10.99275, -10.8093, -10.62548, -10.44128, -10.2567, -10.07175, 
    -9.886418, -9.700713, -9.514633, -9.32818, -9.141355, -8.954158, 
    -8.766592, -8.578656, -8.390352, -8.201681, -8.012645, -7.823244, 
    -7.633479, -7.443353, -7.252865, -7.062018, -6.870813, -6.679251, 
    -6.487333, -6.295061, -6.102437, -5.909461, -5.716136, -5.522462, 
    -5.328442, -5.134077, -4.939369, -4.744318, -4.548928, -4.353199, 
    -4.157134, -3.960734, -3.764001, -3.566937, -3.369543, -3.171822, 
    -2.973775, -2.775405, -2.576714, -2.377702, -2.178374, -1.97873, 
    -1.778772, -1.578504, -1.377926, -1.177042, -0.975853, -0.7743618, 
    -0.5725707, -0.3704818, -0.1680977, 0.03457943, 0.2375471, 0.4408028, 
    0.644344, 0.8481685, 1.052273, 1.256656, 1.461315, 1.666246, 1.871447, 
    2.076916, 2.28265, 2.488645, 2.6949, 2.901411, 3.108176, 3.315192, 
    3.522455, 3.729963, 3.937714, 4.145703, 4.353929, 4.562388, 4.771077, 
    4.979993, 5.189132, 5.398493, 5.608071, 5.817863, 6.027867, 6.238079, 
    6.448495, 6.659113, 6.86993, 7.080941, 7.292144, 7.503535, 7.715111, 
    7.926868, 8.138803, 8.350913, 8.563193, 8.775641, 8.988254, 9.201027, 
    9.413957, 9.62704, 9.840273, 10.05365, 10.26717, 10.48083, 10.69463, 
    10.90856, 11.12261, 11.33679, 11.55109, 11.76551, 11.98004, 12.19468, 
    12.40942, 12.62427, 12.83921, 13.05425, 13.26938, 13.48459, 13.69989, 
    13.91526, 14.13071, 14.34623, 14.56182, 14.77747, 14.99318, 15.20894, 
    15.42476, 15.64062, 15.85652, 16.07247, 16.28845, 16.50446, 16.7205, 
    16.93656, 17.15265, 17.36875, 17.58485, 17.80097, 18.01709, 18.23321, 
    18.44933, 18.66544, 18.88153, 19.09761, 19.31367, 19.52971, 19.74572, 
    19.96169, 20.17763, 20.39353, 20.60939, 20.82519, 21.04095, 21.25665, 
    21.47229, 21.68787, 21.90338, 22.11881, 22.33418, 22.54946, 22.76466, 
    22.97977, 23.1948, 23.40972, 23.62455, 23.83928, 24.0539, 24.26842, 
    24.48281, 24.69709, 24.91125, 25.12529, 25.3392, 25.55297, 25.76661, 
    25.98011, 26.19347, 26.40668, 26.61974, 26.83264, 27.04539, 27.25797, 
    27.4704, 27.68265, 27.89473, 28.10664, 28.31837, 28.52992, 28.74128, 
    28.95245, 29.16343, 29.37422, 29.5848, 29.79519, 30.00537, 30.21534, 
    30.42509, 30.63464, 30.84397, 31.05307, 31.26195, 31.4706, 31.67902, 
    31.88721, 32.09517, 32.30288, 32.51035, 32.71757, 32.92455, 33.13127, 
    33.33774, 33.54396, 33.74991, 33.9556, 34.16103, 34.36619, 34.57108, 
    34.77569, 34.98003, 35.18409, 35.38787, 35.59137, 35.79458, 35.9975, 
    36.20013, 36.40247, 36.60451, 36.80626, 37.0077, 37.20884, 37.40968, 
    37.6102, 37.81042, 38.01033, 38.20993, 38.4092, 38.60817, 38.8068, 
    39.00512, 39.20312, 39.40079, 39.59813, 39.79514, 39.99183, 40.18817, 
    40.38418, 40.57986, 40.7752, 40.97019, 41.16484, 41.35916, 41.55312, 
    41.74674, 41.94001, 42.13293, 42.3255, 42.51772, 42.70958, 42.90108, 
    43.09223, 43.28302, 43.47345, 43.66352, 43.85323, 44.04257, 44.23155, 
    44.42016, 44.60841, 44.79629, 44.9838, 45.17093, 45.3577, 45.54409, 
    45.73011, 45.91576, 46.10103, 46.28593, 46.47044, 46.65458, 46.83834, 
    47.02173, 47.20473, 47.38735, 47.56959, 47.75145, 47.93292, 48.11401, 
    48.29472, 48.47504, 48.65498, 48.83453, 49.01369, 49.19247, 49.37086, 
    49.54886, 49.72648, 49.9037, 50.08054, 50.25699, 50.43305, 50.60872, 
    50.78399, 50.95888, 51.13338, 51.30748, 51.4812, 51.65453, 51.82746, 52, 
    52.17215,
  -30.59251, -30.45487, -30.3169, -30.17858, -30.03992, -29.90092, -29.76157, 
    -29.62188, -29.48185, -29.34146, -29.20074, -29.05966, -28.91823, 
    -28.77645, -28.63433, -28.49184, -28.34901, -28.20582, -28.06228, 
    -27.91838, -27.77413, -27.62952, -27.48455, -27.33922, -27.19353, 
    -27.04748, -26.90106, -26.75429, -26.60715, -26.45964, -26.31178, 
    -26.16354, -26.01494, -25.86597, -25.71663, -25.56692, -25.41685, 
    -25.2664, -25.11558, -24.96438, -24.81282, -24.66088, -24.50856, 
    -24.35588, -24.20281, -24.04937, -23.89555, -23.74135, -23.58677, 
    -23.43182, -23.27648, -23.12077, -22.96467, -22.80819, -22.65133, 
    -22.49408, -22.33645, -22.17844, -22.02004, -21.86126, -21.70209, 
    -21.54254, -21.3826, -21.22227, -21.06155, -20.90045, -20.73895, 
    -20.57707, -20.4148, -20.25214, -20.08908, -19.92564, -19.76181, 
    -19.59758, -19.43297, -19.26796, -19.10256, -18.93677, -18.77058, 
    -18.604, -18.43703, -18.26966, -18.10191, -17.93375, -17.76521, 
    -17.59627, -17.42693, -17.2572, -17.08708, -16.91656, -16.74565, 
    -16.57435, -16.40265, -16.23055, -16.05807, -15.88518, -15.71191, 
    -15.53824, -15.36417, -15.18971, -15.01486, -14.83962, -14.66398, 
    -14.48795, -14.31153, -14.13471, -13.9575, -13.7799, -13.60191, 
    -13.42353, -13.24476, -13.0656, -12.88605, -12.7061, -12.52577, 
    -12.34506, -12.16395, -11.98246, -11.80058, -11.61832, -11.43567, 
    -11.25263, -11.06922, -10.88542, -10.70123, -10.51667, -10.33172, 
    -10.1464, -9.960696, -9.774614, -9.588156, -9.40132, -9.21411, -9.026525, 
    -8.838569, -8.650239, -8.461538, -8.272468, -8.083029, -7.893222, 
    -7.703049, -7.512511, -7.321609, -7.130344, -6.938719, -6.746733, 
    -6.554389, -6.361688, -6.168631, -5.97522, -5.781457, -5.587342, 
    -5.392878, -5.198066, -5.002907, -4.807404, -4.611558, -4.41537, 
    -4.218843, -4.021979, -3.824779, -3.627244, -3.429377, -3.23118, 
    -3.032655, -2.833803, -2.634626, -2.435128, -2.235309, -2.035172, 
    -1.834718, -1.633951, -1.432872, -1.231484, -1.029788, -0.8277874, 
    -0.6254839, -0.42288, -0.2199781, -0.01678063, 0.18671, 0.3904914, 
    0.594561, 0.7989163, 1.003555, 1.208474, 1.413671, 1.619143, 1.824888, 
    2.030903, 2.237185, 2.443732, 2.65054, 2.857607, 3.06493, 3.272506, 
    3.480333, 3.688406, 3.896725, 4.105284, 4.314082, 4.523115, 4.73238, 
    4.941875, 5.151596, 5.361539, 5.571702, 5.782082, 5.992675, 6.203477, 
    6.414487, 6.6257, 6.837114, 7.048724, 7.260528, 7.472521, 7.684701, 
    7.897065, 8.109608, 8.322327, 8.535219, 8.748281, 8.961508, 9.174896, 
    9.388444, 9.602146, 9.816, 10.03, 10.24415, 10.45843, 10.67285, 10.88741, 
    11.10209, 11.3169, 11.53183, 11.74688, 11.96205, 12.17732, 12.3927, 
    12.60818, 12.82376, 13.03944, 13.25521, 13.47106, 13.687, 13.90302, 
    14.11911, 14.33527, 14.5515, 14.7678, 14.98415, 15.20056, 15.41702, 
    15.63353, 15.85009, 16.06668, 16.28331, 16.49997, 16.71666, 16.93337, 
    17.1501, 17.36685, 17.58361, 17.80037, 18.01715, 18.23392, 18.45068, 
    18.66744, 18.88418, 19.10091, 19.31762, 19.53431, 19.75096, 19.96758, 
    20.18417, 20.40072, 20.61722, 20.83367, 21.05008, 21.26642, 21.48271, 
    21.69893, 21.91508, 22.13116, 22.34716, 22.56309, 22.77893, 22.99468, 
    23.21034, 23.42591, 23.64138, 23.85674, 24.07199, 24.28714, 24.50217, 
    24.71708, 24.93187, 25.14654, 25.36107, 25.57547, 25.78974, 26.00386, 
    26.21784, 26.43167, 26.64535, 26.85887, 27.07223, 27.28543, 27.49847, 
    27.71133, 27.92402, 28.13654, 28.34888, 28.56103, 28.77299, 28.98476, 
    29.19634, 29.40772, 29.6189, 29.82988, 30.04065, 30.25121, 30.46156, 
    30.67169, 30.88159, 31.09128, 31.30074, 31.50997, 31.71896, 31.92772, 
    32.13625, 32.34452, 32.55256, 32.76035, 32.96788, 33.17516, 33.38219, 
    33.58896, 33.79546, 34.0017, 34.20768, 34.41338, 34.6188, 34.82396, 
    35.02884, 35.23343, 35.43774, 35.64176, 35.8455, 36.04894, 36.25209, 
    36.45495, 36.65751, 36.85976, 37.06171, 37.26336, 37.4647, 37.66573, 
    37.86645, 38.06685, 38.26694, 38.46671, 38.66615, 38.86528, 39.06408, 
    39.26255, 39.4607, 39.65851, 39.856, 40.05314, 40.24995, 40.44643, 
    40.64256, 40.83835, 41.0338, 41.2289, 41.42366, 41.61807, 41.81213, 
    42.00584, 42.19919, 42.39219, 42.58484, 42.77713, 42.96906, 43.16063, 
    43.35183, 43.54268, 43.73315, 43.92327, 44.11302, 44.3024, 44.49141, 
    44.68005, 44.86832, 45.05622, 45.24375, 45.4309, 45.61768, 45.80407, 
    45.9901, 46.17574, 46.361, 46.54589, 46.73039, 46.91452, 47.09826, 
    47.28161, 47.46458, 47.64717, 47.82938, 48.0112, 48.19263, 48.37367, 
    48.55433, 48.7346, 48.91447, 49.09396, 49.27306, 49.45177, 49.63009, 
    49.80802, 49.98556, 50.1627, 50.33946, 50.51582, 50.69179, 50.86737, 
    51.04255, 51.21734, 51.39173, 51.56573, 51.73934, 51.91256, 52.08538, 
    52.2578,
  -30.69403, -30.55631, -30.41825, -30.27985, -30.14111, -30.00203, 
    -29.86259, -29.72282, -29.58269, -29.44222, -29.3014, -29.16022, 
    -29.0187, -28.87683, -28.7346, -28.59202, -28.44908, -28.30579, 
    -28.16214, -28.01814, -27.87378, -27.72905, -27.58397, -27.43852, 
    -27.29272, -27.14655, -27.00002, -26.85312, -26.70586, -26.55823, 
    -26.41023, -26.26187, -26.11313, -25.96403, -25.81456, -25.66471, 
    -25.5145, -25.36391, -25.21294, -25.06161, -24.90989, -24.7578, 
    -24.60534, -24.4525, -24.29928, -24.14568, -23.9917, -23.83734, -23.6826, 
    -23.52748, -23.37198, -23.21609, -23.05982, -22.90317, -22.74613, 
    -22.5887, -22.43089, -22.2727, -22.11411, -21.95514, -21.79579, 
    -21.63604, -21.4759, -21.31538, -21.15446, -20.99315, -20.83146, 
    -20.66937, -20.50689, -20.34401, -20.18075, -20.01709, -19.85303, 
    -19.68859, -19.52375, -19.35851, -19.19288, -19.02686, -18.86044, 
    -18.69363, -18.52641, -18.35881, -18.19081, -18.02241, -17.85361, 
    -17.68442, -17.51483, -17.34484, -17.17446, -17.00368, -16.83251, 
    -16.66093, -16.48896, -16.3166, -16.14383, -15.97067, -15.79711, 
    -15.62316, -15.4488, -15.27406, -15.09891, -14.92337, -14.74744, 
    -14.5711, -14.39438, -14.21725, -14.03974, -13.86183, -13.68352, 
    -13.50482, -13.32573, -13.14624, -12.96636, -12.78609, -12.60543, 
    -12.42438, -12.24293, -12.0611, -11.87888, -11.69626, -11.51326, 
    -11.32988, -11.1461, -10.96194, -10.7774, -10.59247, -10.40716, 
    -10.22146, -10.03538, -9.848926, -9.662086, -9.474869, -9.287272, 
    -9.099299, -8.91095, -8.722225, -8.533127, -8.343656, -8.153812, 
    -7.963599, -7.773015, -7.582064, -7.390747, -7.199063, -7.007015, 
    -6.814605, -6.621832, -6.4287, -6.235209, -6.041362, -5.847158, 
    -5.652601, -5.457691, -5.26243, -5.066819, -4.870862, -4.674558, 
    -4.47791, -4.280919, -4.083588, -3.885918, -3.687911, -3.489569, 
    -3.290894, -3.091887, -2.892551, -2.692888, -2.4929, -2.292588, 
    -2.091956, -1.891004, -1.689736, -1.488153, -1.286258, -1.084053, 
    -0.8815402, -0.6787218, -0.4756003, -0.2721781, -0.06845753, 0.1355589, 
    0.3398686, 0.5444693, 0.7493582, 0.954533, 1.159991, 1.365729, 1.571746, 
    1.778037, 1.984601, 2.191435, 2.398536, 2.605901, 2.813526, 3.021411, 
    3.229551, 3.437944, 3.646586, 3.855475, 4.064608, 4.273981, 4.483592, 
    4.693437, 4.903513, 5.113818, 5.324348, 5.5351, 5.74607, 5.957256, 
    6.168653, 6.38026, 6.592072, 6.804086, 7.016298, 7.228706, 7.441306, 
    7.654095, 7.867068, 8.080223, 8.293555, 8.507063, 8.72074, 8.934587, 
    9.148595, 9.362764, 9.57709, 9.791568, 10.0062, 10.22097, 10.43588, 
    10.65094, 10.86612, 11.08144, 11.29688, 11.51245, 11.72814, 11.94394, 
    12.15985, 12.37587, 12.59199, 12.80822, 13.02453, 13.24094, 13.45744, 
    13.67403, 13.89069, 14.10743, 14.32424, 14.54112, 14.75806, 14.97507, 
    15.19213, 15.40924, 15.6264, 15.84361, 16.06085, 16.27813, 16.49545, 
    16.71279, 16.93015, 17.14754, 17.36494, 17.58235, 17.79977, 18.0172, 
    18.23462, 18.45204, 18.66945, 18.88685, 19.10423, 19.32159, 19.53893, 
    19.75624, 19.97352, 20.19076, 20.40795, 20.62511, 20.84221, 21.05926, 
    21.27626, 21.49319, 21.71006, 21.92686, 22.14359, 22.36024, 22.57681, 
    22.79329, 23.00969, 23.22599, 23.4422, 23.65831, 23.87431, 24.09021, 
    24.30599, 24.52166, 24.73721, 24.95263, 25.16792, 25.38309, 25.59812, 
    25.81301, 26.02777, 26.24237, 26.45682, 26.67112, 26.88527, 27.09925, 
    27.31307, 27.52672, 27.7402, 27.95351, 28.16663, 28.37958, 28.59234, 
    28.80491, 29.01728, 29.22947, 29.44145, 29.65323, 29.8648, 30.07616, 
    30.28732, 30.49825, 30.70897, 30.91946, 31.12973, 31.33977, 31.54958, 
    31.75916, 31.96849, 32.17759, 32.38643, 32.59504, 32.80339, 33.01149, 
    33.21933, 33.42692, 33.63424, 33.8413, 34.04809, 34.25461, 34.46086, 
    34.66683, 34.87253, 35.07794, 35.28307, 35.48792, 35.69247, 35.89673, 
    36.1007, 36.30437, 36.50775, 36.71082, 36.91359, 37.11606, 37.31821, 
    37.52006, 37.7216, 37.92281, 38.12371, 38.3243, 38.52456, 38.72449, 
    38.9241, 39.12339, 39.32234, 39.52097, 39.71925, 39.91721, 40.11483, 
    40.3121, 40.50904, 40.70563, 40.90188, 41.09779, 41.29334, 41.48854, 
    41.6834, 41.8779, 42.07205, 42.26584, 42.45927, 42.65235, 42.84507, 
    43.03742, 43.22941, 43.42104, 43.61229, 43.80319, 43.99371, 44.18387, 
    44.37365, 44.56306, 44.7521, 44.94077, 45.12906, 45.31697, 45.50451, 
    45.69167, 45.87844, 46.06484, 46.25086, 46.4365, 46.62175, 46.80662, 
    46.9911, 47.1752, 47.35891, 47.54224, 47.72518, 47.90773, 48.08989, 
    48.27166, 48.45304, 48.63403, 48.81463, 48.99484, 49.17466, 49.35408, 
    49.53312, 49.71175, 49.89, 50.06784, 50.2453, 50.42236, 50.59902, 
    50.77529, 50.95117, 51.12664, 51.30173, 51.47641, 51.6507, 51.82459, 
    51.99809, 52.17118, 52.34389,
  -30.79592, -30.65813, -30.51999, -30.38151, -30.24269, -30.10352, -29.964, 
    -29.82414, -29.68393, -29.54336, -29.40245, -29.26118, -29.11957, 
    -28.9776, -28.83527, -28.69259, -28.54955, -28.40616, -28.26241, 
    -28.11829, -27.97382, -27.82899, -27.68379, -27.53823, -27.39231, 
    -27.24603, -27.09937, -26.95236, -26.80497, -26.65722, -26.50909, 
    -26.3606, -26.21174, -26.0625, -25.9129, -25.76291, -25.61256, -25.46183, 
    -25.31072, -25.15924, -25.00739, -24.85515, -24.70253, -24.54954, 
    -24.39616, -24.24241, -24.08827, -23.93375, -23.77885, -23.62356, 
    -23.46789, -23.31184, -23.15539, -22.99857, -22.84135, -22.68375, 
    -22.52576, -22.36738, -22.20861, -22.04946, -21.88991, -21.72997, 
    -21.56964, -21.40891, -21.2478, -21.08629, -20.92439, -20.76209, 
    -20.5994, -20.43632, -20.27284, -20.10896, -19.94469, -19.78003, 
    -19.61496, -19.4495, -19.28365, -19.11739, -18.95074, -18.78369, 
    -18.61624, -18.44839, -18.28014, -18.11149, -17.94245, -17.77301, 
    -17.60316, -17.43292, -17.26228, -17.09124, -16.91979, -16.74795, 
    -16.57571, -16.40307, -16.23003, -16.05659, -15.88275, -15.70851, 
    -15.53387, -15.35883, -15.1834, -15.00756, -14.83132, -14.65469, 
    -14.47766, -14.30023, -14.1224, -13.94418, -13.76556, -13.58654, 
    -13.40712, -13.22731, -13.04711, -12.86651, -12.68551, -12.50412, 
    -12.32234, -12.14016, -11.95759, -11.77464, -11.59128, -11.40754, 
    -11.22341, -11.03889, -10.85398, -10.66869, -10.48301, -10.29694, 
    -10.11049, -9.92365, -9.73643, -9.548828, -9.360845, -9.172482, 
    -8.983739, -8.794618, -8.605121, -8.415247, -8.224998, -8.034376, 
    -7.843382, -7.652016, -7.460281, -7.268177, -7.075706, -6.882868, 
    -6.689667, -6.496102, -6.302176, -6.107889, -5.913244, -5.718242, 
    -5.522884, -5.327172, -5.131108, -4.934694, -4.73793, -4.54082, 
    -4.343364, -4.145564, -3.947423, -3.748941, -3.550122, -3.350966, 
    -3.151476, -2.951654, -2.751502, -2.551022, -2.350215, -2.149085, 
    -1.947633, -1.745861, -1.543772, -1.341368, -1.138651, -0.9356236, 
    -0.7322877, -0.528646, -0.3247008, -0.1204545, 0.08409029, 0.2889312, 
    0.4940657, 0.6994911, 0.905205, 1.111205, 1.317488, 1.524051, 1.730892, 
    1.938008, 2.145396, 2.353054, 2.560979, 2.769167, 2.977616, 3.186323, 
    3.395285, 3.604499, 3.813962, 4.023671, 4.233623, 4.443815, 4.654243, 
    4.864905, 5.075798, 5.286918, 5.498261, 5.709826, 5.921607, 6.133604, 
    6.34581, 6.558225, 6.770843, 6.983662, 7.196678, 7.409888, 7.623288, 
    7.836875, 8.050646, 8.264596, 8.478722, 8.693021, 8.907488, 9.122121, 
    9.336916, 9.551868, 9.766975, 9.982233, 10.19764, 10.41319, 10.62887, 
    10.84469, 11.06065, 11.27673, 11.49294, 11.70926, 11.92571, 12.14226, 
    12.35892, 12.57569, 12.79256, 13.00953, 13.22659, 13.44374, 13.66097, 
    13.87828, 14.09567, 14.31314, 14.53067, 14.74826, 14.96592, 15.18364, 
    15.4014, 15.61922, 15.83708, 16.05498, 16.27292, 16.49089, 16.70889, 
    16.92691, 17.14496, 17.36302, 17.58109, 17.79917, 18.01725, 18.23533, 
    18.45341, 18.67148, 18.88954, 19.10758, 19.3256, 19.54359, 19.76155, 
    19.97949, 20.19738, 20.41524, 20.63305, 20.85081, 21.06851, 21.28616, 
    21.50375, 21.72127, 21.93872, 22.1561, 22.3734, 22.59062, 22.80775, 
    23.0248, 23.24175, 23.4586, 23.67536, 23.892, 24.10854, 24.32496, 
    24.54127, 24.75746, 24.97352, 25.18946, 25.40525, 25.62092, 25.83644, 
    26.05183, 26.26706, 26.48214, 26.69707, 26.91184, 27.12645, 27.34089, 
    27.55516, 27.76926, 27.98318, 28.19692, 28.41048, 28.62385, 28.83703, 
    29.05002, 29.2628, 29.47539, 29.68777, 29.89994, 30.11191, 30.32365, 
    30.53518, 30.74649, 30.95758, 31.16843, 31.37906, 31.58945, 31.7996, 
    32.00952, 32.21919, 32.42861, 32.63779, 32.84671, 33.05537, 33.26378, 
    33.47193, 33.67981, 33.88743, 34.09477, 34.30185, 34.50864, 34.71516, 
    34.9214, 35.12735, 35.33302, 35.5384, 35.74349, 35.94828, 36.15278, 
    36.35698, 36.56088, 36.76447, 36.96776, 37.17074, 37.37341, 37.57576, 
    37.7778, 37.97952, 38.18092, 38.382, 38.58276, 38.78318, 38.98328, 
    39.18306, 39.38249, 39.58159, 39.78036, 39.97879, 40.17688, 40.37462, 
    40.57202, 40.76908, 40.96579, 41.16215, 41.35815, 41.55381, 41.74911, 
    41.94406, 42.13865, 42.33287, 42.52674, 42.72025, 42.91339, 43.10617, 
    43.29859, 43.49063, 43.68231, 43.87362, 44.06456, 44.25512, 44.4453, 
    44.63512, 44.82456, 45.01362, 45.2023, 45.39061, 45.57853, 45.76607, 
    45.95323, 46.14001, 46.3264, 46.51241, 46.69802, 46.88326, 47.06811, 
    47.25256, 47.43663, 47.62031, 47.8036, 47.9865, 48.16901, 48.35112, 
    48.53284, 48.71417, 48.8951, 49.07564, 49.25578, 49.43553, 49.61488, 
    49.79384, 49.9724, 50.15056, 50.32832, 50.50569, 50.68266, 50.85923, 
    51.0354, 51.21117, 51.38655, 51.56152, 51.7361, 51.91027, 52.08405, 
    52.25743, 52.4304,
  -30.8982, -30.76033, -30.62212, -30.48356, -30.34466, -30.2054, -30.0658, 
    -29.92585, -29.78555, -29.6449, -29.5039, -29.36254, -29.22083, 
    -29.07876, -28.93634, -28.79356, -28.65042, -28.50693, -28.36307, 
    -28.21885, -28.07427, -27.92933, -27.78402, -27.63835, -27.49232, 
    -27.34591, -27.19914, -27.052, -26.9045, -26.75662, -26.60837, -26.45975, 
    -26.31076, -26.16139, -26.01165, -25.86153, -25.71104, -25.56017, 
    -25.40892, -25.2573, -25.1053, -24.95291, -24.80015, -24.647, -24.49347, 
    -24.33956, -24.18526, -24.03059, -23.87552, -23.72007, -23.56423, 
    -23.40801, -23.2514, -23.09439, -22.93701, -22.77923, -22.62106, 
    -22.46249, -22.30354, -22.1442, -21.98446, -21.82433, -21.6638, 
    -21.50288, -21.34157, -21.17986, -21.01776, -20.85526, -20.69236, 
    -20.52906, -20.36537, -20.20128, -20.03679, -19.8719, -19.70662, 
    -19.54093, -19.37484, -19.20835, -19.04147, -18.87418, -18.70649, 
    -18.5384, -18.36991, -18.20102, -18.03173, -17.86203, -17.69193, 
    -17.52143, -17.35053, -17.17923, -17.00752, -16.83541, -16.6629, 
    -16.48998, -16.31667, -16.14295, -15.96883, -15.7943, -15.61937, 
    -15.44405, -15.26832, -15.09218, -14.91565, -14.73871, -14.56138, 
    -14.38364, -14.2055, -14.02697, -13.84803, -13.66869, -13.48895, 
    -13.30882, -13.12828, -12.94735, -12.76602, -12.5843, -12.40217, 
    -12.21965, -12.03674, -11.85343, -11.66973, -11.48563, -11.30114, 
    -11.11626, -10.93099, -10.74533, -10.55928, -10.37284, -10.18601, 
    -9.998793, -9.811191, -9.623203, -9.434832, -9.246077, -9.05694, 
    -8.867421, -8.677524, -8.487246, -8.296591, -8.105559, -7.914152, 
    -7.722371, -7.530216, -7.33769, -7.144794, -6.951529, -6.757896, 
    -6.563897, -6.369534, -6.174807, -5.979718, -5.784269, -5.588462, 
    -5.392298, -5.195778, -4.998905, -4.80168, -4.604105, -4.406181, 
    -4.207911, -4.009296, -3.810338, -3.611039, -3.411401, -3.211426, 
    -3.011115, -2.810472, -2.609497, -2.408194, -2.206563, -2.004608, 
    -1.802331, -1.599733, -1.396817, -1.193586, -0.9900409, -0.786185, 
    -0.5820204, -0.3775496, -0.1727749, 0.03230109, 0.2376759, 0.443347, 
    0.6493118, 0.8555676, 1.062112, 1.268942, 1.476055, 1.683449, 1.89112, 
    2.099066, 2.307284, 2.515771, 2.724525, 2.933542, 3.142819, 3.352354, 
    3.562143, 3.772183, 3.982472, 4.193006, 4.403782, 4.614798, 4.826048, 
    5.037532, 5.249245, 5.461185, 5.673347, 5.885728, 6.098326, 6.311137, 
    6.524157, 6.737383, 6.950812, 7.164441, 7.378264, 7.59228, 7.806485, 
    8.020874, 8.235445, 8.450194, 8.665118, 8.880212, 9.095472, 9.310897, 
    9.526481, 9.74222, 9.958112, 10.17415, 10.39034, 10.60666, 10.82312, 
    11.03972, 11.25644, 11.47329, 11.69026, 11.90735, 12.12456, 12.34187, 
    12.55929, 12.7768, 12.99442, 13.21213, 13.42993, 13.64782, 13.86579, 
    14.08384, 14.30196, 14.52014, 14.7384, 14.95672, 15.17509, 15.39352, 
    15.61199, 15.83051, 16.04908, 16.26768, 16.48631, 16.70497, 16.92365, 
    17.14236, 17.36108, 17.57981, 17.79856, 18.0173, 18.23605, 18.45479, 
    18.67352, 18.89224, 19.11094, 19.32962, 19.54828, 19.7669, 19.9855, 
    20.20406, 20.42257, 20.64104, 20.85946, 21.07782, 21.29613, 21.51437, 
    21.73255, 21.95066, 22.1687, 22.38665, 22.60452, 22.82231, 23.04001, 
    23.25761, 23.47511, 23.69251, 23.90981, 24.12699, 24.34406, 24.56102, 
    24.77785, 24.99455, 25.21113, 25.42757, 25.64387, 25.86003, 26.07605, 
    26.29192, 26.50763, 26.72319, 26.93859, 27.15382, 27.36889, 27.58379, 
    27.79851, 28.01305, 28.22741, 28.44159, 28.65557, 28.86937, 29.08296, 
    29.29636, 29.50955, 29.72254, 29.93532, 30.14788, 30.36023, 30.57236, 
    30.78426, 30.99594, 31.20738, 31.4186, 31.62958, 31.84031, 32.05081, 
    32.26106, 32.47106, 32.68081, 32.8903, 33.09954, 33.30851, 33.51723, 
    33.72567, 33.93385, 34.14175, 34.34938, 34.55672, 34.76379, 34.97058, 
    35.17708, 35.38329, 35.58921, 35.79483, 36.00016, 36.20519, 36.40991, 
    36.61434, 36.81845, 37.02226, 37.22575, 37.42894, 37.6318, 37.83435, 
    38.03658, 38.23848, 38.44006, 38.64131, 38.84223, 39.04282, 39.24308, 
    39.443, 39.64259, 39.84183, 40.04074, 40.2393, 40.43751, 40.63538, 
    40.8329, 41.03007, 41.22689, 41.42335, 41.61946, 41.81521, 42.0106, 
    42.20564, 42.4003, 42.59461, 42.78855, 42.98212, 43.17533, 43.36817, 
    43.56064, 43.75273, 43.94445, 44.1358, 44.32677, 44.51737, 44.70759, 
    44.89743, 45.08688, 45.27596, 45.46465, 45.65297, 45.84089, 46.02843, 
    46.21559, 46.40236, 46.58873, 46.77472, 46.96032, 47.14553, 47.33035, 
    47.51478, 47.69881, 47.88245, 48.0657, 48.24855, 48.43101, 48.61307, 
    48.79473, 48.976, 49.15687, 49.33734, 49.51741, 49.69709, 49.87636, 
    50.05523, 50.23371, 50.41178, 50.58946, 50.76673, 50.9436, 51.12007, 
    51.29614, 51.47181, 51.64707, 51.82193, 51.9964, 52.17045, 52.34411, 
    52.51736,
  -31.00087, -30.86293, -30.72463, -30.586, -30.44701, -30.30768, -30.16799, 
    -30.02796, -29.88757, -29.74683, -29.60574, -29.46429, -29.32249, 
    -29.18032, -29.03781, -28.89493, -28.75169, -28.60809, -28.46413, 
    -28.31981, -28.17513, -28.03008, -27.88466, -27.73888, -27.59273, 
    -27.44621, -27.29932, -27.15206, -27.00443, -26.85643, -26.70806, 
    -26.55931, -26.41019, -26.26069, -26.11082, -25.96057, -25.80994, 
    -25.65893, -25.50755, -25.35578, -25.20363, -25.0511, -24.89819, 
    -24.74489, -24.59121, -24.43714, -24.28269, -24.12785, -23.97262, 
    -23.81701, -23.661, -23.50461, -23.34783, -23.19065, -23.03309, 
    -22.87513, -22.71678, -22.55804, -22.3989, -22.23937, -22.07945, 
    -21.91912, -21.75841, -21.59729, -21.43578, -21.27387, -21.11156, 
    -20.94885, -20.78575, -20.62224, -20.45834, -20.29403, -20.12932, 
    -19.96422, -19.79871, -19.6328, -19.46648, -19.29976, -19.13264, 
    -18.96512, -18.79719, -18.62886, -18.46013, -18.29099, -18.12145, 
    -17.9515, -17.78115, -17.61039, -17.43923, -17.26766, -17.09569, 
    -16.92331, -16.75053, -16.57734, -16.40375, -16.22975, -16.05534, 
    -15.88053, -15.70532, -15.5297, -15.35368, -15.17725, -15.00041, 
    -14.82318, -14.64554, -14.46749, -14.28904, -14.11019, -13.93094, 
    -13.75128, -13.57122, -13.39076, -13.2099, -13.02863, -12.84697, 
    -12.6649, -12.48244, -12.29958, -12.11632, -11.93266, -11.7486, 
    -11.56415, -11.3793, -11.19406, -11.00843, -10.8224, -10.63597, 
    -10.44916, -10.26195, -10.07436, -9.886371, -9.697997, -9.509236, 
    -9.320088, -9.130556, -8.940639, -8.75034, -8.559657, -8.368594, 
    -8.177151, -7.98533, -7.793131, -7.600556, -7.407607, -7.214284, 
    -7.020589, -6.826523, -6.632089, -6.437286, -6.242117, -6.046584, 
    -5.850687, -5.654428, -5.45781, -5.260833, -5.063499, -4.865811, 
    -4.667769, -4.469376, -4.270633, -4.071542, -3.872105, -3.672325, 
    -3.472202, -3.271739, -3.070938, -2.869801, -2.668329, -2.466527, 
    -2.264394, -2.061933, -1.859148, -1.656039, -1.452609, -1.24886, 
    -1.044796, -0.840417, -0.6357269, -0.4307278, -0.225422, -0.01981207, 
    0.1860994, 0.3923099, 0.5988169, 0.8056177, 1.01271, 1.22009, 1.427756, 
    1.635705, 1.843935, 2.052442, 2.261223, 2.470276, 2.679598, 2.889186, 
    3.099036, 3.309147, 3.519514, 3.730135, 3.941007, 4.152127, 4.363491, 
    4.575097, 4.78694, 4.999018, 5.211328, 5.423867, 5.63663, 5.849615, 
    6.062819, 6.276237, 6.489867, 6.703705, 6.917747, 7.131991, 7.346433, 
    7.561068, 7.775894, 7.990907, 8.206103, 8.421479, 8.637031, 8.852755, 
    9.068647, 9.284705, 9.500924, 9.7173, 9.93383, 10.15051, 10.36734, 
    10.5843, 10.80141, 11.01865, 11.23602, 11.45352, 11.67114, 11.88888, 
    12.10673, 12.3247, 12.54277, 12.76094, 12.97922, 13.19758, 13.41604, 
    13.63459, 13.85321, 14.07192, 14.2907, 14.50955, 14.72847, 14.94745, 
    15.16648, 15.38558, 15.60472, 15.8239, 16.04313, 16.26239, 16.48169, 
    16.70102, 16.92037, 17.13974, 17.35913, 17.57853, 17.79794, 18.01735, 
    18.23677, 18.45617, 18.67557, 18.89496, 19.11433, 19.33368, 19.553, 
    19.77229, 19.99155, 20.21077, 20.42995, 20.64908, 20.86817, 21.08719, 
    21.30617, 21.52507, 21.74391, 21.96268, 22.18137, 22.39999, 22.61852, 
    22.83697, 23.05532, 23.27357, 23.49173, 23.70979, 23.92774, 24.14557, 
    24.36329, 24.58089, 24.79837, 25.01572, 25.23294, 25.45003, 25.66697, 
    25.88377, 26.10043, 26.31694, 26.53329, 26.74948, 26.96551, 27.18138, 
    27.39708, 27.6126, 27.82795, 28.04312, 28.2581, 28.4729, 28.6875, 
    28.90191, 29.11612, 29.33014, 29.54394, 29.75754, 29.97092, 30.18409, 
    30.39704, 30.60977, 30.82227, 31.03454, 31.24659, 31.45839, 31.66996, 
    31.88128, 32.09237, 32.3032, 32.51378, 32.72411, 32.93418, 33.14399, 
    33.35353, 33.56281, 33.77182, 33.98056, 34.18902, 34.39721, 34.60511, 
    34.81273, 35.02007, 35.22712, 35.43387, 35.64033, 35.84649, 36.05236, 
    36.25792, 36.46318, 36.66813, 36.87277, 37.0771, 37.28111, 37.48481, 
    37.68819, 37.89125, 38.09398, 38.29639, 38.49847, 38.70022, 38.90164, 
    39.10272, 39.30347, 39.50388, 39.70395, 39.90368, 40.10306, 40.30209, 
    40.50078, 40.69912, 40.89711, 41.09474, 41.29202, 41.48893, 41.6855, 
    41.8817, 42.07754, 42.27301, 42.46812, 42.66287, 42.85725, 43.05125, 
    43.24489, 43.43815, 43.63104, 43.82356, 44.0157, 44.20746, 44.39884, 
    44.58984, 44.78047, 44.97071, 45.16056, 45.35003, 45.53912, 45.72782, 
    45.91613, 46.10406, 46.29159, 46.47873, 46.66549, 46.85185, 47.03782, 
    47.22339, 47.40857, 47.59336, 47.77774, 47.96174, 48.14533, 48.32853, 
    48.51133, 48.69373, 48.87573, 49.05733, 49.23853, 49.41933, 49.59973, 
    49.77972, 49.95932, 50.13851, 50.3173, 50.49568, 50.67366, 50.85124, 
    51.02841, 51.20518, 51.38155, 51.55751, 51.73306, 51.90821, 52.08296, 
    52.2573, 52.43123, 52.60476,
  -31.10393, -30.96591, -30.82754, -30.68882, -30.54976, -30.41035, 
    -30.27058, -30.13046, -29.98999, -29.84916, -29.70798, -29.56644, 
    -29.42455, -29.28229, -29.13968, -28.9967, -28.85337, -28.70967, 
    -28.56561, -28.42118, -28.27639, -28.13123, -27.9857, -27.83981, 
    -27.69355, -27.54692, -27.39991, -27.25253, -27.10479, -26.95666, 
    -26.80817, -26.65929, -26.51004, -26.36042, -26.21041, -26.06003, 
    -25.90926, -25.75812, -25.60659, -25.45468, -25.30239, -25.14971, 
    -24.99665, -24.8432, -24.68937, -24.53515, -24.38054, -24.22554, 
    -24.07015, -23.91438, -23.75821, -23.60165, -23.44469, -23.28735, 
    -23.12961, -22.97148, -22.81295, -22.65402, -22.4947, -22.33499, 
    -22.17487, -22.01436, -21.85345, -21.69214, -21.53043, -21.36832, 
    -21.20581, -21.0429, -20.87958, -20.71587, -20.55175, -20.38723, 
    -20.2223, -20.05697, -19.89124, -19.72511, -19.55856, -19.39161, 
    -19.22426, -19.0565, -18.88834, -18.71977, -18.55079, -18.3814, 
    -18.21161, -18.04141, -17.87081, -17.69979, -17.52837, -17.35654, 
    -17.1843, -17.01166, -16.8386, -16.66514, -16.49127, -16.31699, 
    -16.14231, -15.96721, -15.79171, -15.6158, -15.43948, -15.26276, 
    -15.08562, -14.90808, -14.73014, -14.55178, -14.37302, -14.19386, 
    -14.01429, -13.83431, -13.65392, -13.47314, -13.29195, -13.11035, 
    -12.92835, -12.74595, -12.56314, -12.37994, -12.19633, -12.01232, 
    -11.82791, -11.6431, -11.4579, -11.27229, -11.08629, -10.89989, -10.7131, 
    -10.52591, -10.33832, -10.15034, -9.961975, -9.773214, -9.584063, 
    -9.394522, -9.204592, -9.014275, -8.823572, -8.632483, -8.441011, 
    -8.249156, -8.056919, -7.864301, -7.671305, -7.477931, -7.284179, 
    -7.090053, -6.895553, -6.700681, -6.505438, -6.309825, -6.113845, 
    -5.917498, -5.720786, -5.523712, -5.326275, -5.128479, -4.930326, 
    -4.731815, -4.53295, -4.333733, -4.134164, -3.934247, -3.733982, 
    -3.533373, -3.33242, -3.131126, -2.929493, -2.727523, -2.525218, 
    -2.32258, -2.119612, -1.916315, -1.712693, -1.508746, -1.304478, 
    -1.099891, -0.8949873, -0.689769, -0.4842388, -0.2783991, -0.07225253, 
    0.1341985, 0.3409513, 0.5480033, 0.7553518, 0.9629943, 1.170928, 1.37915, 
    1.587658, 1.796448, 2.005519, 2.214867, 2.424489, 2.634383, 2.844545, 
    3.054972, 3.265661, 3.476611, 3.687816, 3.899274, 4.110983, 4.322938, 
    4.535137, 4.747577, 4.960253, 5.173164, 5.386305, 5.599673, 5.813265, 
    6.027078, 6.241108, 6.455351, 6.669805, 6.884465, 7.099328, 7.314391, 
    7.52965, 7.745101, 7.960741, 8.176566, 8.392572, 8.608757, 8.825116, 
    9.041644, 9.25834, 9.475198, 9.692215, 9.909388, 10.12671, 10.34418, 
    10.5618, 10.77955, 10.99744, 11.21546, 11.43361, 11.65189, 11.87028, 
    12.08879, 12.30741, 12.52614, 12.74497, 12.96391, 13.18293, 13.40205, 
    13.62126, 13.84055, 14.05992, 14.27937, 14.49889, 14.71847, 14.93812, 
    15.15782, 15.37758, 15.59739, 15.81725, 16.03714, 16.25708, 16.47705, 
    16.69704, 16.91707, 17.13711, 17.35717, 17.57724, 17.79732, 18.01741, 
    18.23749, 18.45757, 18.67764, 18.8977, 19.11774, 19.33776, 19.55775, 
    19.77771, 19.99764, 20.21754, 20.43738, 20.65718, 20.87694, 21.09663, 
    21.31627, 21.53584, 21.75535, 21.97478, 22.19414, 22.41342, 22.63261, 
    22.85172, 23.07073, 23.28965, 23.50847, 23.72718, 23.94578, 24.16427, 
    24.38265, 24.6009, 24.81903, 25.03703, 25.2549, 25.47264, 25.69023, 
    25.90768, 26.12498, 26.34212, 26.55912, 26.77595, 26.99262, 27.20912, 
    27.42545, 27.64161, 27.85759, 28.07338, 28.28899, 28.50441, 28.71964, 
    28.93467, 29.1495, 29.36413, 29.57855, 29.79276, 30.00676, 30.22054, 
    30.43409, 30.64743, 30.86053, 31.0734, 31.28604, 31.49845, 31.71061, 
    31.92252, 32.13419, 32.34561, 32.55677, 32.76768, 32.97833, 33.18872, 
    33.39884, 33.60869, 33.81827, 34.02757, 34.2366, 34.44534, 34.6538, 
    34.86198, 35.06987, 35.27747, 35.48477, 35.69177, 35.89848, 36.10488, 
    36.31098, 36.51677, 36.72225, 36.92742, 37.13227, 37.33681, 37.54103, 
    37.74492, 37.94849, 38.15174, 38.35466, 38.55724, 38.75949, 38.96141, 
    39.16299, 39.36423, 39.56513, 39.76568, 39.96589, 40.16576, 40.36527, 
    40.56443, 40.76324, 40.96169, 41.15979, 41.35753, 41.55491, 41.75193, 
    41.94858, 42.14487, 42.34079, 42.53635, 42.73153, 42.92635, 43.12078, 
    43.31485, 43.50854, 43.70186, 43.89479, 44.08735, 44.27953, 44.47132, 
    44.66273, 44.85376, 45.04441, 45.23466, 45.42453, 45.61401, 45.8031, 
    45.9918, 46.18011, 46.36802, 46.55554, 46.74267, 46.9294, 47.11574, 
    47.30168, 47.48722, 47.67236, 47.85711, 48.04145, 48.2254, 48.40894, 
    48.59209, 48.77483, 48.95717, 49.1391, 49.32063, 49.50176, 49.68248, 
    49.8628, 50.04272, 50.22223, 50.40133, 50.58002, 50.75831, 50.9362, 
    51.11367, 51.29074, 51.4674, 51.64365, 51.8195, 51.99493, 52.16996, 
    52.34459, 52.5188, 52.6926,
  -31.20737, -31.06928, -30.93084, -30.79204, -30.6529, -30.51341, -30.37356, 
    -30.23336, -30.0928, -29.95189, -29.81062, -29.66899, -29.52701, 
    -29.38466, -29.24195, -29.09888, -28.95545, -28.81165, -28.66749, 
    -28.52296, -28.37806, -28.2328, -28.08716, -27.94116, -27.79478, 
    -27.64804, -27.50092, -27.35343, -27.20556, -27.05731, -26.90869, 
    -26.7597, -26.61032, -26.46056, -26.31042, -26.15991, -26.00901, 
    -25.85773, -25.70606, -25.55401, -25.40158, -25.24875, -25.09554, 
    -24.94195, -24.78796, -24.63359, -24.47882, -24.32367, -24.16812, 
    -24.01218, -23.85584, -23.69912, -23.542, -23.38448, -23.22657, 
    -23.06826, -22.90955, -22.75045, -22.59094, -22.43104, -22.27074, 
    -22.11004, -21.94893, -21.78743, -21.62552, -21.46321, -21.3005, 
    -21.13738, -20.97386, -20.80994, -20.64561, -20.48087, -20.31573, 
    -20.15018, -19.98422, -19.81786, -19.65109, -19.48392, -19.31633, 
    -19.14833, -18.97993, -18.81112, -18.6419, -18.47227, -18.30223, 
    -18.13177, -17.96091, -17.78964, -17.61796, -17.44587, -17.27337, 
    -17.10045, -16.92713, -16.75339, -16.57924, -16.40468, -16.22972, 
    -16.05434, -15.87855, -15.70234, -15.52573, -15.34871, -15.17128, 
    -14.99344, -14.81518, -14.63652, -14.45745, -14.27797, -14.09808, 
    -13.91778, -13.73707, -13.55596, -13.37444, -13.19251, -13.01018, 
    -12.82744, -12.64429, -12.46074, -12.27678, -12.09242, -11.90766, 
    -11.72249, -11.53693, -11.35096, -11.16459, -10.97782, -10.79065, 
    -10.60309, -10.41512, -10.22676, -10.03801, -9.848858, -9.659314, 
    -9.469378, -9.279051, -9.088333, -8.897225, -8.705729, -8.513846, 
    -8.321577, -8.128923, -7.935885, -7.742465, -7.548665, -7.354484, 
    -7.159925, -6.964989, -6.769678, -6.573992, -6.377934, -6.181505, 
    -5.984706, -5.78754, -5.590007, -5.39211, -5.19385, -4.995228, -4.796247, 
    -4.596909, -4.397215, -4.197166, -3.996766, -3.796016, -3.594917, 
    -3.393472, -3.191683, -2.989552, -2.78708, -2.584271, -2.381126, 
    -2.177648, -1.973838, -1.769699, -1.565233, -1.360443, -1.155331, 
    -0.9498992, -0.74415, -0.5380861, -0.3317097, -0.1250237, 0.08196963, 
    0.2892676, 0.4968675, 0.7047668, 0.9129628, 1.121453, 1.330234, 1.539303, 
    1.748658, 1.958296, 2.168213, 2.378408, 2.588876, 2.799615, 3.010623, 
    3.221895, 3.433429, 3.645222, 3.85727, 4.069571, 4.282121, 4.494917, 
    4.707956, 4.921235, 5.134749, 5.348497, 5.562474, 5.776677, 5.991102, 
    6.205747, 6.420608, 6.635681, 6.850962, 7.066449, 7.282137, 7.498023, 
    7.714104, 7.930375, 8.146832, 8.363474, 8.580296, 8.797292, 9.014461, 
    9.231797, 9.449299, 9.666961, 9.88478, 10.10275, 10.32087, 10.53914, 
    10.75754, 10.97609, 11.19477, 11.41357, 11.6325, 11.85155, 12.07072, 
    12.29001, 12.5094, 12.7289, 12.94849, 13.16819, 13.38797, 13.60785, 
    13.82781, 14.04785, 14.26796, 14.48815, 14.7084, 14.92872, 15.1491, 
    15.36953, 15.59001, 15.81054, 16.03112, 16.25173, 16.47237, 16.69304, 
    16.91374, 17.13446, 17.35519, 17.57594, 17.7967, 18.01746, 18.23822, 
    18.45898, 18.67972, 18.90046, 19.12117, 19.34187, 19.56254, 19.78317, 
    20.00378, 20.22434, 20.44487, 20.66534, 20.88577, 21.10613, 21.32644, 
    21.54668, 21.76686, 21.98697, 22.20699, 22.42694, 22.6468, 22.86657, 
    23.08625, 23.30583, 23.52531, 23.74469, 23.96395, 24.1831, 24.40214, 
    24.62105, 24.83983, 25.05849, 25.27701, 25.4954, 25.71364, 25.93174, 
    26.14968, 26.36748, 26.58512, 26.80259, 27.0199, 27.23705, 27.45401, 
    27.67081, 27.88742, 28.10385, 28.32009, 28.53614, 28.752, 28.96765, 
    29.18311, 29.39835, 29.61339, 29.82822, 30.04283, 30.25722, 30.47139, 
    30.68533, 30.89904, 31.11252, 31.32576, 31.53876, 31.75152, 31.96403, 
    32.17629, 32.3883, 32.60005, 32.81154, 33.02277, 33.23374, 33.44444, 
    33.65486, 33.86501, 34.07488, 34.28448, 34.49379, 34.70281, 34.91154, 
    35.11999, 35.32814, 35.53599, 35.74355, 35.95079, 36.15774, 36.36438, 
    36.5707, 36.77672, 36.98242, 37.1878, 37.39286, 37.5976, 37.80201, 
    38.0061, 38.20986, 38.41328, 38.61637, 38.81913, 39.02155, 39.22363, 
    39.42536, 39.62675, 39.82779, 40.02849, 40.22884, 40.42883, 40.62846, 
    40.82775, 41.02667, 41.22523, 41.42344, 41.62128, 41.81875, 42.01586, 
    42.2126, 42.40897, 42.60497, 42.8006, 42.99585, 43.19073, 43.38523, 
    43.57935, 43.77309, 43.96645, 44.15942, 44.35202, 44.54422, 44.73605, 
    44.92748, 45.11853, 45.30919, 45.49945, 45.68932, 45.8788, 46.06789, 
    46.25658, 46.44488, 46.63278, 46.82029, 47.00739, 47.1941, 47.3804, 
    47.56631, 47.75181, 47.93691, 48.12161, 48.30591, 48.4898, 48.67329, 
    48.85637, 49.03905, 49.22132, 49.40318, 49.58464, 49.76569, 49.94633, 
    50.12656, 50.30639, 50.4858, 50.66481, 50.84341, 51.0216, 51.19937, 
    51.37674, 51.5537, 51.73024, 51.90638, 52.08211, 52.25742, 52.43232, 
    52.60682, 52.7809,
  -31.31121, -31.17304, -31.03453, -30.89566, -30.75644, -30.61687, 
    -30.47694, -30.33666, -30.19602, -30.05502, -29.91367, -29.77195, 
    -29.62987, -29.48743, -29.34463, -29.20147, -29.05794, -28.91404, 
    -28.76978, -28.62515, -28.48015, -28.33478, -28.18904, -28.04292, 
    -27.89644, -27.74958, -27.60234, -27.45473, -27.30675, -27.15838, 
    -27.00964, -26.86052, -26.71102, -26.56113, -26.41087, -26.26022, 
    -26.10918, -25.95777, -25.80596, -25.65377, -25.50119, -25.34822, 
    -25.19487, -25.04112, -24.88699, -24.73246, -24.57754, -24.42223, 
    -24.26652, -24.11042, -23.95392, -23.79703, -23.63974, -23.48205, 
    -23.32397, -23.16548, -23.0066, -22.84731, -22.68763, -22.52754, 
    -22.36705, -22.20616, -22.04486, -21.88316, -21.72106, -21.55855, 
    -21.39564, -21.23232, -21.06859, -20.90445, -20.73991, -20.57496, 
    -20.4096, -20.24383, -20.07766, -19.91107, -19.74407, -19.57667, 
    -19.40885, -19.24062, -19.07198, -18.90292, -18.73346, -18.56358, 
    -18.39329, -18.22259, -18.05148, -17.87995, -17.708, -17.53565, 
    -17.36288, -17.1897, -17.0161, -16.84209, -16.66767, -16.49283, 
    -16.31758, -16.14191, -15.96584, -15.78934, -15.61244, -15.43512, 
    -15.25739, -15.07924, -14.90068, -14.72171, -14.54233, -14.36253, 
    -14.18232, -14.0017, -13.82067, -13.63923, -13.45738, -13.27512, 
    -13.09245, -12.90937, -12.72588, -12.54198, -12.35768, -12.17296, 
    -11.98785, -11.80232, -11.61639, -11.43006, -11.24332, -11.05618, 
    -10.86864, -10.6807, -10.49236, -10.30361, -10.11447, -9.924932, 
    -9.734996, -9.544664, -9.353937, -9.162817, -8.971304, -8.779399, 
    -8.587104, -8.39442, -8.201346, -8.007888, -7.814043, -7.619814, 
    -7.425202, -7.230208, -7.034835, -6.839083, -6.642953, -6.446448, 
    -6.249569, -6.052317, -5.854693, -5.656701, -5.458341, -5.259614, 
    -5.060524, -4.86107, -4.661256, -4.461082, -4.260552, -4.059667, 
    -3.858428, -3.656838, -3.454899, -3.252613, -3.049981, -2.847006, 
    -2.64369, -2.440035, -2.236044, -2.031719, -1.827061, -1.622074, 
    -1.416759, -1.211119, -1.005156, -0.7988735, -0.5922731, -0.3853574, 
    -0.178129, 0.02940953, 0.2372555, 0.4454063, 0.6538593, 0.8626117, 
    1.071661, 1.281004, 1.490638, 1.700561, 1.910769, 2.121259, 2.332029, 
    2.543075, 2.754395, 2.965986, 3.177844, 3.389967, 3.60235, 3.814992, 
    4.027889, 4.241037, 4.454434, 4.668076, 4.88196, 5.096082, 5.31044, 
    5.525029, 5.739847, 5.954889, 6.170153, 6.385634, 6.60133, 6.817237, 
    7.033351, 7.249668, 7.466186, 7.682899, 7.899806, 8.1169, 8.334181, 
    8.551642, 8.769281, 8.987095, 9.205077, 9.423226, 9.641538, 9.860007, 
    10.07863, 10.29741, 10.51633, 10.73539, 10.95459, 11.17393, 11.39339, 
    11.61299, 11.8327, 12.05254, 12.27249, 12.49254, 12.71271, 12.93297, 
    13.15334, 13.3738, 13.59434, 13.81497, 14.03569, 14.25648, 14.47734, 
    14.69827, 14.91926, 15.14032, 15.36143, 15.58259, 15.8038, 16.02505, 
    16.24634, 16.46766, 16.68901, 16.91039, 17.13179, 17.35321, 17.57463, 
    17.79607, 18.01751, 18.23895, 18.46039, 18.68182, 18.90323, 19.12463, 
    19.346, 19.56735, 19.78867, 20.00995, 20.2312, 20.4524, 20.67355, 
    20.89465, 21.1157, 21.33668, 21.5576, 21.77845, 21.99923, 22.21993, 
    22.44055, 22.66108, 22.88153, 23.10187, 23.32212, 23.54227, 23.76231, 
    23.98224, 24.20206, 24.42176, 24.64133, 24.86078, 25.08009, 25.29927, 
    25.51831, 25.73721, 25.95596, 26.17456, 26.39301, 26.61129, 26.82941, 
    27.04737, 27.26516, 27.48277, 27.7002, 27.91745, 28.13452, 28.35139, 
    28.56808, 28.78456, 29.00085, 29.21693, 29.4328, 29.64847, 29.86391, 
    30.07914, 30.29415, 30.50893, 30.72348, 30.9378, 31.15189, 31.36573, 
    31.57934, 31.7927, 32.00581, 32.21866, 32.43126, 32.6436, 32.85569, 
    33.0675, 33.27905, 33.49033, 33.70133, 33.91206, 34.1225, 34.33266, 
    34.54254, 34.75213, 34.96143, 35.17043, 35.37914, 35.58754, 35.79564, 
    36.00344, 36.21093, 36.41811, 36.62497, 36.83152, 37.03776, 37.24367, 
    37.44926, 37.65452, 37.85946, 38.06406, 38.26833, 38.47227, 38.67587, 
    38.87914, 39.08206, 39.28463, 39.48687, 39.68875, 39.89029, 40.09147, 
    40.2923, 40.49277, 40.69289, 40.89264, 41.09204, 41.29107, 41.48974, 
    41.68805, 41.88598, 42.08354, 42.28074, 42.47756, 42.674, 42.87007, 
    43.06577, 43.26108, 43.45601, 43.65056, 43.84473, 44.03852, 44.23191, 
    44.42492, 44.61755, 44.80978, 45.00163, 45.19307, 45.38413, 45.5748, 
    45.76507, 45.95494, 46.14442, 46.3335, 46.52217, 46.71046, 46.89833, 
    47.08581, 47.27289, 47.45956, 47.64583, 47.8317, 48.01715, 48.20221, 
    48.38686, 48.5711, 48.75493, 48.93835, 49.12137, 49.30398, 49.48617, 
    49.66796, 49.84933, 50.0303, 50.21086, 50.391, 50.57073, 50.75005, 
    50.92896, 51.10745, 51.28553, 51.4632, 51.64045, 51.81729, 51.99372, 
    52.16973, 52.34533, 52.52052, 52.69529, 52.86964,
  -31.41544, -31.2772, -31.13862, -30.99968, -30.86038, -30.72073, -30.58072, 
    -30.44036, -30.29964, -30.15856, -30.01711, -29.87531, -29.73315, 
    -29.59062, -29.44773, -29.30447, -29.16084, -29.01685, -28.87248, 
    -28.72775, -28.58265, -28.43718, -28.29133, -28.14511, -27.99851, 
    -27.85154, -27.70419, -27.55647, -27.40836, -27.25988, -27.11102, 
    -26.96177, -26.81214, -26.66213, -26.51174, -26.36095, -26.20979, 
    -26.05824, -25.90629, -25.75396, -25.60124, -25.44813, -25.29463, 
    -25.14074, -24.98645, -24.83177, -24.6767, -24.52123, -24.36536, 
    -24.2091, -24.05244, -23.89538, -23.73792, -23.58006, -23.42181, 
    -23.26315, -23.10409, -22.94462, -22.78476, -22.62449, -22.46381, 
    -22.30273, -22.14124, -21.97935, -21.81705, -21.65434, -21.49122, 
    -21.3277, -21.16376, -20.99942, -20.83467, -20.6695, -20.50393, 
    -20.33794, -20.17154, -20.00473, -19.83751, -19.66987, -19.50182, 
    -19.33336, -19.16448, -18.99518, -18.82548, -18.65535, -18.48482, 
    -18.31386, -18.14249, -17.97071, -17.79851, -17.62589, -17.45285, 
    -17.2794, -17.10554, -16.93125, -16.75655, -16.58143, -16.4059, 
    -16.22995, -16.05358, -15.8768, -15.6996, -15.52198, -15.34395, -15.1655, 
    -14.98663, -14.80735, -14.62766, -14.44755, -14.26702, -14.08608, 
    -13.90472, -13.72295, -13.54077, -13.35818, -13.17517, -12.99175, 
    -12.80791, -12.62367, -12.43902, -12.25395, -12.06848, -11.8826, 
    -11.69631, -11.50961, -11.3225, -11.13499, -10.94707, -10.75875, 
    -10.57003, -10.3809, -10.19137, -10.00144, -9.811111, -9.620382, 
    -9.429255, -9.23773, -9.045811, -8.853496, -8.660787, -8.467686, 
    -8.274194, -8.080312, -7.88604, -7.691382, -7.496337, -7.300908, 
    -7.105095, -6.9089, -6.712325, -6.515371, -6.318039, -6.120332, -5.92225, 
    -5.723796, -5.524971, -5.325776, -5.126214, -4.926286, -4.725994, 
    -4.525341, -4.324326, -4.122953, -3.921224, -3.719141, -3.516705, 
    -3.313919, -3.110784, -2.907303, -2.703478, -2.499311, -2.294805, 
    -2.089961, -1.884782, -1.679271, -1.473428, -1.267258, -1.060762, 
    -0.8539431, -0.6468033, -0.4393454, -0.2315719, -0.02348532, 0.1849116, 
    0.3936162, 0.6026258, 0.8119378, 1.021549, 1.231457, 1.441659, 1.652153, 
    1.862934, 2.074, 2.285349, 2.496977, 2.708881, 2.921058, 3.133506, 
    3.34622, 3.559198, 3.772437, 3.985933, 4.199683, 4.413684, 4.627933, 
    4.842426, 5.05716, 5.272131, 5.487336, 5.702772, 5.918435, 6.134321, 
    6.350428, 6.566751, 6.783287, 7.000032, 7.216982, 7.434135, 7.651486, 
    7.869031, 8.086767, 8.30469, 8.522797, 8.741082, 8.959544, 9.178177, 
    9.396977, 9.615942, 9.835067, 10.05435, 10.27378, 10.49336, 10.71308, 
    10.93295, 11.15295, 11.37308, 11.59334, 11.81372, 12.03423, 12.25485, 
    12.47558, 12.69641, 12.91735, 13.13839, 13.35952, 13.58075, 13.80205, 
    14.02345, 14.24491, 14.46645, 14.68807, 14.90974, 15.13148, 15.35327, 
    15.57511, 15.797, 16.01894, 16.24091, 16.46292, 16.68495, 16.90702, 
    17.1291, 17.3512, 17.57332, 17.79544, 18.01757, 18.23969, 18.46182, 
    18.68393, 18.90603, 19.12811, 19.35017, 19.5722, 19.7942, 20.01617, 
    20.2381, 20.45998, 20.68182, 20.9036, 21.12533, 21.34699, 21.56859, 
    21.79012, 22.01158, 22.23296, 22.45425, 22.67546, 22.89658, 23.11761, 
    23.33853, 23.55935, 23.78006, 24.00066, 24.22115, 24.44151, 24.66175, 
    24.88186, 25.10184, 25.32168, 25.54138, 25.76094, 25.98035, 26.19961, 
    26.4187, 26.63764, 26.85642, 27.07502, 27.29346, 27.51172, 27.72979, 
    27.94769, 28.16539, 28.38291, 28.60023, 28.81735, 29.03427, 29.25098, 
    29.46748, 29.68377, 29.89984, 30.11569, 30.33132, 30.54672, 30.76189, 
    30.97682, 31.19152, 31.40597, 31.62018, 31.83414, 32.04786, 32.26131, 
    32.47451, 32.68745, 32.90012, 33.11252, 33.32466, 33.53652, 33.7481, 
    33.9594, 34.17043, 34.38116, 34.59161, 34.80177, 35.01163, 35.22119, 
    35.43046, 35.63942, 35.84807, 36.05642, 36.26446, 36.47218, 36.67959, 
    36.88668, 37.09345, 37.29989, 37.50601, 37.7118, 37.91726, 38.12239, 
    38.32718, 38.53163, 38.73574, 38.93951, 39.14294, 39.34602, 39.54875, 
    39.75113, 39.95316, 40.15483, 40.35615, 40.55711, 40.7577, 40.95794, 
    41.15781, 41.35731, 41.55645, 41.75521, 41.95361, 42.15163, 42.34928, 
    42.54655, 42.74345, 42.93996, 43.13609, 43.33185, 43.52721, 43.7222, 
    43.9168, 44.11101, 44.30483, 44.49826, 44.6913, 44.88394, 45.07619, 
    45.26805, 45.45951, 45.65058, 45.84124, 46.03151, 46.22138, 46.41084, 
    46.59991, 46.78857, 46.97683, 47.16468, 47.35213, 47.53917, 47.7258, 
    47.91203, 48.09784, 48.28325, 48.46825, 48.65284, 48.83702, 49.02079, 
    49.20414, 49.38708, 49.56962, 49.75174, 49.93344, 50.11473, 50.2956, 
    50.47606, 50.65611, 50.83574, 51.01495, 51.19375, 51.37214, 51.5501, 
    51.72765, 51.90479, 52.08151, 52.25781, 52.43369, 52.60916, 52.78421, 
    52.95885,
  -31.52007, -31.38177, -31.2431, -31.10409, -30.96472, -30.82499, -30.68491, 
    -30.54447, -30.40366, -30.2625, -30.12097, -29.97908, -29.83683, 
    -29.69421, -29.55123, -29.40788, -29.26416, -29.12007, -28.97561, 
    -28.83077, -28.68557, -28.53999, -28.39404, -28.24771, -28.10101, 
    -27.95393, -27.80647, -27.65863, -27.5104, -27.3618, -27.21282, 
    -27.06345, -26.9137, -26.76356, -26.61304, -26.46213, -26.31083, 
    -26.15914, -26.00706, -25.85459, -25.70173, -25.54848, -25.39483, 
    -25.24079, -25.08636, -24.93153, -24.7763, -24.62067, -24.46465, 
    -24.30823, -24.1514, -23.99418, -23.83655, -23.67853, -23.5201, 
    -23.36126, -23.20203, -23.04238, -22.88234, -22.72188, -22.56102, 
    -22.39975, -22.23807, -22.07598, -21.91349, -21.75058, -21.58727, 
    -21.42354, -21.2594, -21.09485, -20.92988, -20.76451, -20.59871, 
    -20.43251, -20.26589, -20.09885, -19.9314, -19.76354, -19.59525, 
    -19.42655, -19.25744, -19.0879, -18.91795, -18.74759, -18.5768, 
    -18.40559, -18.23397, -18.06193, -17.88947, -17.71659, -17.54329, 
    -17.36957, -17.19543, -17.02087, -16.84589, -16.6705, -16.49468, 
    -16.31844, -16.14179, -15.96471, -15.78722, -15.6093, -15.43097, 
    -15.25222, -15.07304, -14.89345, -14.71344, -14.53302, -14.35217, 
    -14.17091, -13.98923, -13.80713, -13.62462, -13.44169, -13.25834, 
    -13.07458, -12.8904, -12.70581, -12.52081, -12.33539, -12.14956, 
    -11.96332, -11.77666, -11.5896, -11.40213, -11.21424, -11.02595, 
    -10.83725, -10.64814, -10.45863, -10.26871, -10.07839, -9.887664, 
    -9.696536, -9.505008, -9.313078, -9.120749, -8.928023, -8.7349, 
    -8.541381, -8.347467, -8.153161, -7.958462, -7.763372, -7.567894, 
    -7.372026, -7.175773, -6.979134, -6.782112, -6.584707, -6.386921, 
    -6.188757, -5.990215, -5.791297, -5.592005, -5.39234, -5.192305, -4.9919, 
    -4.791129, -4.589992, -4.388491, -4.186629, -3.984407, -3.781828, 
    -3.578893, -3.375605, -3.171965, -2.967976, -2.76364, -2.558958, 
    -2.353934, -2.14857, -1.942867, -1.736828, -1.530456, -1.323752, 
    -1.11672, -0.9093623, -0.7016804, -0.4936775, -0.2853559, -0.07671843, 
    0.1322324, 0.3414938, 0.5510631, 0.7609376, 0.9711144, 1.181591, 
    1.392364, 1.603431, 1.814789, 2.026434, 2.238365, 2.450578, 2.663069, 
    2.875837, 3.088877, 3.302186, 3.515763, 3.729602, 3.943701, 4.158056, 
    4.372665, 4.587524, 4.80263, 5.017979, 5.233568, 5.449393, 5.665451, 
    5.881738, 6.098251, 6.314986, 6.53194, 6.749109, 6.966489, 7.184077, 
    7.401869, 7.619861, 7.83805, 8.056431, 8.275002, 8.493756, 8.712693, 
    8.931807, 9.151093, 9.37055, 9.590173, 9.809957, 10.0299, 10.24999, 
    10.47024, 10.69063, 10.91116, 11.13183, 11.35263, 11.57356, 11.79461, 
    12.01579, 12.23708, 12.45849, 12.68, 12.90162, 13.12334, 13.34515, 
    13.56705, 13.78904, 14.01112, 14.23327, 14.4555, 14.67779, 14.90015, 
    15.12257, 15.34505, 15.56758, 15.79016, 16.01278, 16.23545, 16.45814, 
    16.68087, 16.90362, 17.1264, 17.34919, 17.57199, 17.79481, 18.01762, 
    18.24044, 18.46325, 18.68605, 18.90884, 19.13161, 19.35436, 19.57709, 
    19.79978, 20.02243, 20.24505, 20.46762, 20.69014, 20.91261, 21.13503, 
    21.35738, 21.57966, 21.80188, 22.02402, 22.24608, 22.46805, 22.68994, 
    22.91174, 23.13344, 23.35504, 23.57654, 23.79793, 24.0192, 24.24036, 
    24.4614, 24.68231, 24.90309, 25.12374, 25.34424, 25.56461, 25.78483, 
    26.0049, 26.22482, 26.44458, 26.66418, 26.88361, 27.10287, 27.32195, 
    27.54086, 27.75958, 27.97813, 28.19648, 28.41463, 28.6326, 28.85036, 
    29.06791, 29.28526, 29.50239, 29.71931, 29.93601, 30.15249, 30.36874, 
    30.58476, 30.80055, 31.0161, 31.23141, 31.44648, 31.6613, 31.87587, 
    32.09018, 32.30424, 32.51804, 32.73158, 32.94484, 33.15784, 33.37056, 
    33.58301, 33.79518, 34.00706, 34.21866, 34.42998, 34.641, 34.85172, 
    35.06215, 35.27228, 35.48211, 35.69163, 35.90084, 36.10974, 36.31833, 
    36.5266, 36.73455, 36.94218, 37.14949, 37.35647, 37.56312, 37.76944, 
    37.97543, 38.18108, 38.38639, 38.59136, 38.79599, 39.00027, 39.2042, 
    39.40778, 39.61102, 39.8139, 40.01642, 40.21859, 40.42039, 40.62183, 
    40.82291, 41.02362, 41.22397, 41.42395, 41.62355, 41.82279, 42.02164, 
    42.22013, 42.41823, 42.61596, 42.8133, 43.01027, 43.20684, 43.40303, 
    43.59884, 43.79426, 43.98928, 44.18392, 44.37817, 44.57202, 44.76548, 
    44.95854, 45.1512, 45.34346, 45.53533, 45.7268, 45.91786, 46.10852, 
    46.29878, 46.48864, 46.67808, 46.86713, 47.05576, 47.24399, 47.43181, 
    47.61922, 47.80622, 47.99281, 48.17898, 48.36475, 48.5501, 48.73504, 
    48.91956, 49.10368, 49.28737, 49.47065, 49.65351, 49.83596, 50.01799, 
    50.19961, 50.38081, 50.56158, 50.74195, 50.92189, 51.10141, 51.28052, 
    51.45921, 51.63747, 51.81532, 51.99275, 52.16976, 52.34635, 52.52252, 
    52.69827, 52.8736, 53.04851,
  -31.6251, -31.48672, -31.34799, -31.20891, -31.06946, -30.92966, -30.7895, 
    -30.64898, -30.5081, -30.36685, -30.22524, -30.08327, -29.94093, 
    -29.79822, -29.65515, -29.5117, -29.36789, -29.22371, -29.07915, 
    -28.93422, -28.78891, -28.64323, -28.49718, -28.35074, -28.20393, 
    -28.05674, -27.90916, -27.76121, -27.61287, -27.46416, -27.31505, 
    -27.16556, -27.01569, -26.86542, -26.71477, -26.56373, -26.4123, 
    -26.26048, -26.10827, -25.95566, -25.80266, -25.64927, -25.49547, 
    -25.34129, -25.1867, -25.03172, -24.87634, -24.72056, -24.56438, 
    -24.4078, -24.25081, -24.09343, -23.93563, -23.77744, -23.61884, 
    -23.45983, -23.30042, -23.1406, -22.98037, -22.81973, -22.65868, 
    -22.49722, -22.33536, -22.17308, -22.01039, -21.84728, -21.68377, 
    -21.51984, -21.35549, -21.19073, -21.02556, -20.85997, -20.69396, 
    -20.52753, -20.36069, -20.19344, -20.02576, -19.85766, -19.68915, 
    -19.52021, -19.35086, -19.18109, -19.01089, -18.84028, -18.66924, 
    -18.49779, -18.32591, -18.15361, -17.98089, -17.80775, -17.63418, 
    -17.4602, -17.28579, -17.11095, -16.9357, -16.76002, -16.58392, -16.4074, 
    -16.23046, -16.05309, -15.8753, -15.69709, -15.51845, -15.33939, 
    -15.15991, -14.98001, -14.79969, -14.61895, -14.43778, -14.2562, 
    -14.07419, -13.89177, -13.70892, -13.52566, -13.34197, -13.15787, 
    -12.97335, -12.78841, -12.60306, -12.41728, -12.2311, -12.04449, 
    -11.85748, -11.67004, -11.4822, -11.29394, -11.10527, -10.91619, 
    -10.7267, -10.5368, -10.3465, -10.15578, -9.964659, -9.773131, -9.5812, 
    -9.388864, -9.196126, -9.002987, -8.809447, -8.615509, -8.421173, 
    -8.22644, -8.031312, -7.83579, -7.639875, -7.443569, -7.246873, 
    -7.049788, -6.852317, -6.65446, -6.456219, -6.257595, -6.058591, 
    -5.859207, -5.659446, -5.45931, -5.258799, -5.057916, -4.856662, 
    -4.65504, -4.453052, -4.250698, -4.047982, -3.844904, -3.641468, 
    -3.437675, -3.233528, -3.029028, -2.824178, -2.618979, -2.413435, 
    -2.207547, -2.001318, -1.794749, -1.587845, -1.380606, -1.173035, 
    -0.9651347, -0.756908, -0.5483571, -0.3394847, -0.1302933, 0.07921428, 
    0.2890355, 0.4991675, 0.7096076, 0.9203529, 1.131401, 1.342748, 1.554392, 
    1.76633, 1.978558, 2.191074, 2.403875, 2.616957, 2.830318, 3.043954, 
    3.257863, 3.47204, 3.686483, 3.901189, 4.116154, 4.331374, 4.546847, 
    4.762569, 4.978537, 5.194747, 5.411196, 5.62788, 5.844795, 6.061938, 
    6.279306, 6.496895, 6.714701, 6.932721, 7.15095, 7.369385, 7.588023, 
    7.806859, 8.025889, 8.245111, 8.46452, 8.684111, 8.903881, 9.123827, 
    9.343944, 9.564228, 9.784675, 10.00528, 10.22604, 10.44696, 10.66802, 
    10.88922, 11.11056, 11.33204, 11.55364, 11.77537, 11.99723, 12.2192, 
    12.44129, 12.66348, 12.88578, 13.10818, 13.33068, 13.55327, 13.77595, 
    13.99871, 14.22155, 14.44446, 14.66745, 14.8905, 15.11361, 15.33678, 
    15.56, 15.78327, 16.00659, 16.22994, 16.45333, 16.67676, 16.9002, 
    17.12367, 17.34716, 17.57066, 17.79417, 18.01768, 18.24119, 18.4647, 
    18.68819, 18.91168, 19.13515, 19.35859, 19.582, 19.80539, 20.02874, 
    20.25205, 20.47531, 20.69853, 20.92169, 21.14479, 21.36783, 21.59081, 
    21.81371, 22.03654, 22.25928, 22.48195, 22.70452, 22.92701, 23.14939, 
    23.37167, 23.59385, 23.81592, 24.03787, 24.25971, 24.48142, 24.70301, 
    24.92446, 25.14578, 25.36696, 25.588, 25.80889, 26.02962, 26.25021, 
    26.47063, 26.69089, 26.91098, 27.1309, 27.35064, 27.5702, 27.78958, 
    28.00877, 28.22777, 28.44658, 28.66518, 28.88358, 29.10178, 29.31977, 
    29.53754, 29.75509, 29.97243, 30.18953, 30.40641, 30.62306, 30.83947, 
    31.05564, 31.27157, 31.48725, 31.70269, 31.91787, 32.13279, 32.34745, 
    32.56186, 32.77599, 32.98986, 33.20345, 33.41677, 33.62981, 33.84256, 
    34.05503, 34.26722, 34.47911, 34.6907, 34.902, 35.113, 35.3237, 35.53409, 
    35.74417, 35.95395, 36.16341, 36.37255, 36.58137, 36.78987, 36.99804, 
    37.20589, 37.41341, 37.62059, 37.82745, 38.03396, 38.24014, 38.44597, 
    38.65146, 38.85661, 39.0614, 39.26585, 39.46994, 39.67367, 39.87705, 
    40.08007, 40.28273, 40.48503, 40.68696, 40.88852, 41.08972, 41.29054, 
    41.49099, 41.69107, 41.89077, 42.0901, 42.28904, 42.4876, 42.68578, 
    42.88358, 43.08099, 43.27801, 43.47465, 43.67089, 43.86674, 44.06221, 
    44.25727, 44.45194, 44.64621, 44.84009, 45.03357, 45.22664, 45.41932, 
    45.61159, 45.80346, 45.99492, 46.18597, 46.37663, 46.56687, 46.7567, 
    46.94613, 47.13514, 47.32375, 47.51194, 47.69972, 47.88708, 48.07404, 
    48.26057, 48.4467, 48.6324, 48.81769, 49.00256, 49.18702, 49.37106, 
    49.55467, 49.73787, 49.92065, 50.10301, 50.28495, 50.46647, 50.64757, 
    50.82824, 51.0085, 51.18834, 51.36774, 51.54674, 51.7253, 51.90345, 
    52.08117, 52.25847, 52.43535, 52.61181, 52.78784, 52.96345, 53.13864,
  -31.73053, -31.59209, -31.45329, -31.31413, -31.17462, -31.03474, -30.8945, 
    -30.7539, -30.61294, -30.47162, -30.32992, -30.18787, -30.04544, 
    -29.90265, -29.75948, -29.61595, -29.47204, -29.32776, -29.18311, 
    -29.03808, -28.89268, -28.7469, -28.60074, -28.4542, -28.30728, 
    -28.15998, -28.01229, -27.86423, -27.71578, -27.56694, -27.41772, 
    -27.26811, -27.11811, -26.96772, -26.81695, -26.66578, -26.51422, 
    -26.36226, -26.20991, -26.05717, -25.90403, -25.75049, -25.59656, 
    -25.44223, -25.2875, -25.13237, -24.97683, -24.8209, -24.66456, 
    -24.50782, -24.35067, -24.19312, -24.03517, -23.8768, -23.71803, 
    -23.55885, -23.39926, -23.23927, -23.07886, -22.91804, -22.7568, 
    -22.59516, -22.4331, -22.27063, -22.10775, -21.94444, -21.78073, 
    -21.61659, -21.45205, -21.28708, -21.12169, -20.95589, -20.78967, 
    -20.62303, -20.45596, -20.28848, -20.12058, -19.95226, -19.78351, 
    -19.61434, -19.44475, -19.27474, -19.1043, -18.93344, -18.76216, 
    -18.59045, -18.41832, -18.24576, -18.07278, -17.89938, -17.72555, 
    -17.55129, -17.37661, -17.20151, -17.02597, -16.85002, -16.67363, 
    -16.49683, -16.31959, -16.14193, -15.96385, -15.78534, -15.6064, 
    -15.42704, -15.24725, -15.06704, -14.88641, -14.70535, -14.52386, 
    -14.34195, -14.15962, -13.97687, -13.79369, -13.61009, -13.42606, 
    -13.24162, -13.05675, -12.87147, -12.68576, -12.49963, -12.31309, 
    -12.12612, -11.93874, -11.75094, -11.56273, -11.37409, -11.18505, 
    -10.99559, -10.80571, -10.61543, -10.42473, -10.23362, -10.0421, 
    -9.850171, -9.657835, -9.465092, -9.271943, -9.07839, -8.884434, 
    -8.690074, -8.495314, -8.300154, -8.104595, -7.908638, -7.712286, 
    -7.515539, -7.318399, -7.120867, -6.922945, -6.724634, -6.525935, 
    -6.326851, -6.127382, -5.927531, -5.7273, -5.526689, -5.325701, 
    -5.124337, -4.9226, -4.72049, -4.518012, -4.315164, -4.111951, -3.908373, 
    -3.704434, -3.500134, -3.295477, -3.090464, -2.885097, -2.679379, 
    -2.473312, -2.266898, -2.060139, -1.853039, -1.645599, -1.437821, 
    -1.229709, -1.021264, -0.8124897, -0.6033881, -0.3939619, -0.1842137, 
    0.02585376, 0.2362377, 0.4469355, 0.6579443, 0.8692613, 1.080884, 
    1.292808, 1.505033, 1.717553, 1.930368, 2.143472, 2.356865, 2.570541, 
    2.784499, 2.998735, 3.213246, 3.428028, 3.643079, 3.858394, 4.073972, 
    4.289808, 4.505898, 4.722241, 4.938831, 5.155666, 5.372742, 5.590056, 
    5.807603, 6.025382, 6.243386, 6.461614, 6.680061, 6.898724, 7.117599, 
    7.336681, 7.555968, 7.775455, 7.99514, 8.215016, 8.435082, 8.655334, 
    8.875765, 9.096374, 9.317155, 9.538105, 9.75922, 9.980496, 10.20193, 
    10.42352, 10.64525, 10.86713, 11.08915, 11.3113, 11.53359, 11.756, 
    11.97854, 12.20119, 12.42396, 12.64684, 12.86983, 13.09292, 13.31611, 
    13.53939, 13.76276, 13.98621, 14.20974, 14.43335, 14.65703, 14.88077, 
    15.10458, 15.32845, 15.55237, 15.77634, 16.00035, 16.2244, 16.44849, 
    16.67261, 16.89676, 17.12093, 17.34511, 17.56931, 17.79352, 18.01773, 
    18.24195, 18.46615, 18.69035, 18.91453, 19.1387, 19.36284, 19.58696, 
    19.81104, 20.03509, 20.25909, 20.48306, 20.70697, 20.93082, 21.15462, 
    21.37836, 21.60203, 21.82562, 22.04914, 22.27258, 22.49594, 22.7192, 
    22.94238, 23.16545, 23.38842, 23.61128, 23.83404, 24.05667, 24.27919, 
    24.50159, 24.72385, 24.94598, 25.16798, 25.38984, 25.61155, 25.83311, 
    26.05452, 26.27577, 26.49686, 26.71778, 26.93854, 27.15912, 27.37952, 
    27.59974, 27.81978, 28.03962, 28.25928, 28.47873, 28.69799, 28.91704, 
    29.13588, 29.35451, 29.57292, 29.79111, 30.00908, 30.22682, 30.44434, 
    30.66161, 30.87865, 31.09545, 31.312, 31.5283, 31.74435, 31.96015, 
    32.17568, 32.39096, 32.60596, 32.82071, 33.03517, 33.24936, 33.46328, 
    33.67691, 33.89025, 34.10332, 34.31608, 34.52856, 34.74073, 34.95261, 
    35.16418, 35.37545, 35.58641, 35.79706, 36.0074, 36.21741, 36.42711, 
    36.63649, 36.84554, 37.05426, 37.26265, 37.47071, 37.67844, 37.88582, 
    38.09287, 38.29957, 38.50593, 38.71194, 38.91761, 39.12292, 39.32787, 
    39.53247, 39.73672, 39.9406, 40.14412, 40.34727, 40.55006, 40.75249, 
    40.95454, 41.15622, 41.35752, 41.55845, 41.759, 41.95917, 42.15896, 
    42.35837, 42.55739, 42.75603, 42.95428, 43.15214, 43.34961, 43.54669, 
    43.74337, 43.93966, 44.13556, 44.33105, 44.52615, 44.72084, 44.91514, 
    45.10904, 45.30252, 45.49561, 45.68829, 45.88056, 46.07242, 46.26387, 
    46.45492, 46.64555, 46.83578, 47.02559, 47.21498, 47.40396, 47.59253, 
    47.78068, 47.96841, 48.15573, 48.34262, 48.5291, 48.71516, 48.90081, 
    49.08603, 49.27082, 49.4552, 49.63916, 49.82269, 50.0058, 50.18849, 
    50.37076, 50.5526, 50.73402, 50.91501, 51.09558, 51.27572, 51.45544, 
    51.63474, 51.8136, 51.99205, 52.17006, 52.34766, 52.52482, 52.70156, 
    52.87788, 53.05377, 53.22923,
  -31.83637, -31.69786, -31.55899, -31.41976, -31.28017, -31.14023, 
    -30.99991, -30.85924, -30.7182, -30.5768, -30.43502, -30.29288, 
    -30.15037, -30.00749, -29.86424, -29.72062, -29.57662, -29.43225, 
    -29.2875, -29.14237, -28.99687, -28.85099, -28.70473, -28.55808, 
    -28.41106, -28.26365, -28.11586, -27.96768, -27.81911, -27.67016, 
    -27.52082, -27.37109, -27.22097, -27.07046, -26.91956, -26.76826, 
    -26.61657, -26.46449, -26.312, -26.15912, -26.00585, -25.85217, -25.6981, 
    -25.54362, -25.38874, -25.23346, -25.07778, -24.92169, -24.76519, 
    -24.6083, -24.45099, -24.29328, -24.13515, -23.97662, -23.81768, 
    -23.65833, -23.49857, -23.33839, -23.1778, -23.0168, -22.85539, 
    -22.69356, -22.53131, -22.36865, -22.20557, -22.04207, -21.87815, 
    -21.71382, -21.54906, -21.38389, -21.2183, -21.05228, -20.88584, 
    -20.71898, -20.5517, -20.384, -20.21587, -20.04732, -19.87834, -19.70894, 
    -19.53911, -19.36886, -19.19818, -19.02707, -18.85554, -18.68359, 
    -18.5112, -18.33839, -18.16515, -17.99148, -17.81738, -17.64286, 
    -17.46791, -17.29253, -17.11672, -16.94048, -16.76382, -16.58672, 
    -16.4092, -16.23125, -16.05287, -15.87406, -15.69482, -15.51516, 
    -15.33506, -15.15454, -14.97359, -14.79221, -14.61041, -14.42818, 
    -14.24552, -14.06243, -13.87892, -13.69499, -13.51062, -13.32584, 
    -13.14062, -12.95499, -12.76893, -12.58245, -12.39554, -12.20822, 
    -12.02047, -11.8323, -11.64371, -11.45471, -11.26528, -11.07544, 
    -10.88518, -10.6945, -10.50341, -10.31191, -10.11999, -9.927659, 
    -9.734918, -9.541766, -9.348206, -9.154237, -8.959862, -8.76508, 
    -8.569895, -8.374306, -8.178314, -7.981922, -7.785131, -7.587942, 
    -7.390356, -7.192375, -6.993999, -6.795232, -6.596075, -6.396528, 
    -6.196594, -5.996274, -5.795569, -5.594482, -5.393015, -5.191168, 
    -4.988945, -4.786346, -4.583375, -4.380032, -4.176319, -3.972239, 
    -3.767793, -3.562985, -3.357815, -3.152286, -2.946401, -2.74016, 
    -2.533568, -2.326626, -2.119336, -1.9117, -1.703722, -1.495403, 
    -1.286747, -1.077754, -0.8684294, -0.658774, -0.4487911, -0.2384831, 
    -0.02785284, 0.183097, 0.3943636, 0.6059442, 0.817836, 1.030036, 
    1.242541, 1.455349, 1.668456, 1.88186, 2.095557, 2.309544, 2.523818, 
    2.738376, 2.953215, 3.168332, 3.383723, 3.599385, 3.815314, 4.031508, 
    4.247963, 4.464675, 4.681642, 4.898859, 5.116323, 5.33403, 5.551977, 
    5.770161, 5.988577, 6.207222, 6.426093, 6.645185, 6.864496, 7.08402, 
    7.303754, 7.523695, 7.743838, 7.96418, 8.184717, 8.405444, 8.626358, 
    8.847455, 9.068731, 9.290182, 9.511803, 9.733591, 9.955541, 10.17765, 
    10.39991, 10.62232, 10.84488, 11.06758, 11.29042, 11.51339, 11.73649, 
    11.95972, 12.18306, 12.40652, 12.63009, 12.85377, 13.07755, 13.30143, 
    13.52541, 13.74947, 13.97362, 14.19785, 14.42216, 14.64654, 14.87099, 
    15.09549, 15.32006, 15.54468, 15.76935, 15.99407, 16.21883, 16.44362, 
    16.66844, 16.89329, 17.11816, 17.34306, 17.56796, 17.79287, 18.01779, 
    18.24271, 18.46762, 18.69252, 18.91741, 19.14228, 19.36712, 19.59194, 
    19.81673, 20.04148, 20.26619, 20.49085, 20.71547, 20.94002, 21.16452, 
    21.38896, 21.61333, 21.83762, 22.06184, 22.28597, 22.51003, 22.73399, 
    22.95785, 23.18162, 23.40528, 23.62883, 23.85228, 24.0756, 24.29881, 
    24.52189, 24.74484, 24.96765, 25.19033, 25.41287, 25.63526, 25.85749, 
    26.07958, 26.3015, 26.52327, 26.74486, 26.96628, 27.18753, 27.4086, 
    27.62948, 27.85018, 28.07069, 28.291, 28.51111, 28.73102, 28.95072, 
    29.17021, 29.38949, 29.60854, 29.82738, 30.04599, 30.26437, 30.48251, 
    30.70042, 30.91809, 31.13552, 31.3527, 31.56962, 31.78629, 32.00271, 
    32.21886, 32.43475, 32.65037, 32.86572, 33.08079, 33.29558, 33.51009, 
    33.72432, 33.93827, 34.15192, 34.36527, 34.57833, 34.79109, 35.00355, 
    35.2157, 35.42754, 35.63908, 35.85029, 36.06119, 36.27177, 36.48203, 
    36.69196, 36.90156, 37.11084, 37.31977, 37.52838, 37.73664, 37.94457, 
    38.15215, 38.35938, 38.56627, 38.77281, 38.97899, 39.18482, 39.39029, 
    39.59541, 39.80016, 40.00455, 40.20857, 40.41222, 40.61551, 40.81842, 
    41.02096, 41.22312, 41.42491, 41.62632, 41.82734, 42.02798, 42.22824, 
    42.42812, 42.62761, 42.8267, 43.02541, 43.22372, 43.42164, 43.61916, 
    43.81629, 44.01302, 44.20934, 44.40527, 44.6008, 44.79592, 44.99063, 
    45.18495, 45.37885, 45.57235, 45.76543, 45.95811, 46.15038, 46.34223, 
    46.53367, 46.72469, 46.9153, 47.1055, 47.29527, 47.48463, 47.67357, 
    47.86209, 48.05019, 48.23788, 48.42514, 48.61197, 48.79839, 48.98438, 
    49.16995, 49.35509, 49.53981, 49.72411, 49.90798, 50.09142, 50.27444, 
    50.45703, 50.63919, 50.82093, 51.00224, 51.18312, 51.36358, 51.54361, 
    51.7232, 51.90237, 52.08111, 52.25943, 52.43731, 52.61477, 52.79179, 
    52.96839, 53.14456, 53.3203,
  -31.94261, -31.80404, -31.6651, -31.5258, -31.38615, -31.24613, -31.10574, 
    -30.96499, -30.82388, -30.68239, -30.54054, -30.39832, -30.25572, 
    -30.11276, -29.96942, -29.82571, -29.68162, -29.53716, -29.39231, 
    -29.24709, -29.10149, -28.95551, -28.80915, -28.6624, -28.51527, 
    -28.36776, -28.21985, -28.07157, -27.92289, -27.77382, -27.62437, 
    -27.47452, -27.32428, -27.17365, -27.02262, -26.87119, -26.71937, 
    -26.56716, -26.41454, -26.26153, -26.10811, -25.9543, -25.80008, 
    -25.64546, -25.49044, -25.33501, -25.17917, -25.02293, -24.86628, 
    -24.70923, -24.55176, -24.39389, -24.2356, -24.0769, -23.91779, 
    -23.75827, -23.59834, -23.43798, -23.27722, -23.11603, -22.95444, 
    -22.79242, -22.62998, -22.46713, -22.30386, -22.14016, -21.97605, 
    -21.81151, -21.64655, -21.48117, -21.31537, -21.14914, -20.98249, 
    -20.81541, -20.64791, -20.47998, -20.31163, -20.14285, -19.97364, 
    -19.80401, -19.63394, -19.46345, -19.29253, -19.12118, -18.9494, 
    -18.77719, -18.60456, -18.43149, -18.25799, -18.08406, -17.9097, 
    -17.73491, -17.55968, -17.38403, -17.20794, -17.03143, -16.85448, 
    -16.6771, -16.49928, -16.32104, -16.14236, -15.96325, -15.78372, 
    -15.60375, -15.42334, -15.24251, -15.06125, -14.87955, -14.69743, 
    -14.51487, -14.33189, -14.14847, -13.96463, -13.78035, -13.59565, 
    -13.41052, -13.22496, -13.03898, -12.85256, -12.66573, -12.47846, 
    -12.29077, -12.10266, -11.91412, -11.72516, -11.53578, -11.34597, 
    -11.15575, -10.9651, -10.77404, -10.58255, -10.39065, -10.19833, 
    -10.0056, -9.812453, -9.618892, -9.424917, -9.230532, -9.035736, 
    -8.840531, -8.644918, -8.448899, -8.252474, -8.055645, -7.858413, 
    -7.66078, -7.462747, -7.264315, -7.065485, -6.866261, -6.666642, 
    -6.466631, -6.266229, -6.065437, -5.864258, -5.662694, -5.460745, 
    -5.258414, -5.055702, -4.852612, -4.649146, -4.445304, -4.24109, 
    -4.036505, -3.831552, -3.626231, -3.420547, -3.2145, -3.008093, 
    -2.801328, -2.594208, -2.386734, -2.17891, -1.970737, -1.762218, 
    -1.553355, -1.344151, -1.134609, -0.9247306, -0.7145187, -0.503976, 
    -0.2931053, -0.08190918, 0.1296096, 0.3414482, 0.5536037, 0.7660735, 
    0.9788544, 1.191944, 1.405338, 1.619035, 1.833031, 2.047324, 2.261909, 
    2.476785, 2.691947, 2.907393, 3.123118, 3.339122, 3.555398, 3.771945, 
    3.988759, 4.205837, 4.423174, 4.640769, 4.858616, 5.076713, 5.295055, 
    5.51364, 5.732464, 5.951523, 6.170813, 6.390331, 6.610073, 6.830034, 
    7.050212, 7.270602, 7.491201, 7.712004, 7.933008, 8.154209, 8.375602, 
    8.597184, 8.818951, 9.040898, 9.263022, 9.485319, 9.707784, 9.930412, 
    10.1532, 10.37615, 10.59924, 10.82249, 11.04587, 11.2694, 11.49306, 
    11.71685, 11.94076, 12.1648, 12.38896, 12.61322, 12.8376, 13.06208, 
    13.28666, 13.51133, 13.7361, 13.96095, 14.18588, 14.41089, 14.63597, 
    14.86113, 15.08634, 15.31161, 15.53694, 15.76232, 15.98774, 16.21321, 
    16.43871, 16.66424, 16.8898, 17.11538, 17.34098, 17.5666, 17.79222, 
    18.01785, 18.24347, 18.46909, 18.6947, 18.9203, 19.14588, 19.37144, 
    19.59696, 19.82246, 20.04792, 20.27333, 20.4987, 20.72402, 20.94929, 
    21.17449, 21.39963, 21.6247, 21.8497, 22.07462, 22.29946, 22.52421, 
    22.74887, 22.97344, 23.1979, 23.42226, 23.64651, 23.87064, 24.09466, 
    24.31856, 24.54233, 24.76597, 24.98947, 25.21284, 25.43606, 25.65913, 
    25.88205, 26.10481, 26.32742, 26.54986, 26.77213, 26.99422, 27.21614, 
    27.43788, 27.65943, 27.88079, 28.10196, 28.32294, 28.54371, 28.76427, 
    28.98463, 29.20477, 29.4247, 29.64441, 29.86389, 30.08314, 30.30217, 
    30.52095, 30.7395, 30.9578, 31.17586, 31.39367, 31.61122, 31.82852, 
    32.04556, 32.26233, 32.47883, 32.69506, 32.91103, 33.12671, 33.34211, 
    33.55722, 33.77205, 33.9866, 34.20084, 34.41479, 34.62844, 34.84179, 
    35.05482, 35.26756, 35.47998, 35.69208, 35.90387, 36.11534, 36.32648, 
    36.5373, 36.74779, 36.95795, 37.16778, 37.37727, 37.58642, 37.79523, 
    38.00369, 38.21181, 38.41958, 38.627, 38.83406, 39.04077, 39.24712, 
    39.45311, 39.65873, 39.86399, 40.06889, 40.27342, 40.47757, 40.68135, 
    40.88476, 41.08779, 41.29044, 41.49271, 41.6946, 41.89611, 42.09723, 
    42.29795, 42.49829, 42.69825, 42.8978, 43.09696, 43.29573, 43.4941, 
    43.69207, 43.88964, 44.08681, 44.28357, 44.47993, 44.67589, 44.87144, 
    45.06658, 45.26131, 45.45563, 45.64954, 45.84303, 46.03611, 46.22878, 
    46.42104, 46.61287, 46.80429, 46.99529, 47.18587, 47.37603, 47.56576, 
    47.75508, 47.94397, 48.13244, 48.32049, 48.50811, 48.69531, 48.88208, 
    49.06842, 49.25434, 49.43983, 49.6249, 49.80953, 49.99374, 50.17751, 
    50.36086, 50.54378, 50.72626, 50.90832, 51.08995, 51.27114, 51.45191, 
    51.63224, 51.81215, 51.99162, 52.17065, 52.34926, 52.52744, 52.70518, 
    52.8825, 53.05938, 53.23582, 53.41184,
  -32.04926, -31.91062, -31.77162, -31.63226, -31.49253, -31.35244, 
    -31.21198, -31.07116, -30.92997, -30.78841, -30.64647, -30.50417, 
    -30.3615, -30.21845, -30.07502, -29.93122, -29.78705, -29.64249, 
    -29.49756, -29.35224, -29.20654, -29.06046, -28.914, -28.76715, 
    -28.61992, -28.4723, -28.32429, -28.17589, -28.0271, -27.87792, 
    -27.72835, -27.57839, -27.42803, -27.27727, -27.12612, -26.97457, 
    -26.82262, -26.67028, -26.51753, -26.36438, -26.21083, -26.05688, 
    -25.90252, -25.74776, -25.59259, -25.43701, -25.28103, -25.12464, 
    -24.96783, -24.81062, -24.653, -24.49496, -24.33651, -24.17765, 
    -24.01837, -23.85868, -23.69857, -23.53804, -23.3771, -23.21573, 
    -23.05395, -22.89175, -22.72913, -22.56608, -22.40261, -22.23873, 
    -22.07441, -21.90968, -21.74451, -21.57893, -21.41292, -21.24648, 
    -21.07961, -20.91232, -20.7446, -20.57645, -20.40787, -20.23886, 
    -20.06942, -19.89955, -19.72925, -19.55852, -19.38736, -19.21577, 
    -19.04374, -18.87128, -18.69839, -18.52507, -18.35131, -18.17711, 
    -18.00249, -17.82743, -17.65194, -17.47601, -17.29964, -17.12285, 
    -16.94561, -16.76795, -16.58985, -16.41131, -16.23234, -16.05293, 
    -15.87309, -15.69281, -15.5121, -15.33096, -15.14938, -14.96737, 
    -14.78492, -14.60204, -14.41873, -14.23499, -14.05081, -13.8662, 
    -13.68115, -13.49568, -13.30977, -13.12344, -12.93667, -12.74948, 
    -12.56185, -12.3738, -12.18532, -11.99641, -11.80708, -11.61732, 
    -11.42713, -11.23652, -11.04549, -10.85403, -10.66215, -10.46986, 
    -10.27714, -10.084, -9.890444, -9.696471, -9.502083, -9.30728, -9.112062, 
    -8.916432, -8.720391, -8.52394, -8.32708, -8.129811, -7.932137, 
    -7.734059, -7.535576, -7.336692, -7.137407, -6.937723, -6.737641, 
    -6.537164, -6.336292, -6.135027, -5.933372, -5.731327, -5.528895, 
    -5.326077, -5.122875, -4.919291, -4.715328, -4.510986, -4.306268, 
    -4.101176, -3.895712, -3.689878, -3.483676, -3.277109, -3.070178, 
    -2.862886, -2.655236, -2.447228, -2.238867, -2.030154, -1.821091, 
    -1.611682, -1.401928, -1.191832, -0.9813973, -0.7706259, -0.5595206, 
    -0.3480841, -0.136319, 0.07577174, 0.2881854, 0.5009191, 0.71397, 
    0.9273351, 1.141012, 1.354996, 1.569286, 1.783879, 1.99877, 2.213957, 
    2.429437, 2.645207, 2.861263, 3.077602, 3.294221, 3.511116, 3.728284, 
    3.945722, 4.163426, 4.381393, 4.599619, 4.8181, 5.036834, 5.255816, 
    5.475043, 5.69451, 5.914216, 6.134155, 6.354324, 6.574719, 6.795336, 
    7.016172, 7.237222, 7.458483, 7.679951, 7.901621, 8.12349, 8.345553, 
    8.567808, 8.79025, 9.012873, 9.235675, 9.458652, 9.681797, 9.905109, 
    10.12858, 10.35221, 10.576, 10.79993, 11.02401, 11.24823, 11.47258, 
    11.69707, 11.92168, 12.14642, 12.37127, 12.59624, 12.82131, 13.0465, 
    13.27178, 13.49716, 13.72263, 13.94819, 14.17383, 14.39955, 14.62534, 
    14.8512, 15.07712, 15.30311, 15.52915, 15.75524, 15.98137, 16.20755, 
    16.43376, 16.66001, 16.88628, 17.11258, 17.3389, 17.56522, 17.79156, 
    18.0179, 18.24424, 18.47058, 18.69691, 18.92322, 19.14951, 19.37578, 
    19.60202, 19.82823, 20.0544, 20.28053, 20.50661, 20.73264, 20.95862, 
    21.18453, 21.41038, 21.63616, 21.86187, 22.0875, 22.31304, 22.5385, 
    22.76386, 22.98913, 23.2143, 23.43936, 23.66431, 23.88914, 24.11386, 
    24.33845, 24.56292, 24.78725, 25.01144, 25.2355, 25.45941, 25.68317, 
    25.90678, 26.13023, 26.35351, 26.57663, 26.79958, 27.02235, 27.24495, 
    27.46736, 27.68959, 27.91162, 28.13346, 28.35509, 28.57653, 28.79776, 
    29.01878, 29.23958, 29.46016, 29.68052, 29.90065, 30.12055, 30.34022, 
    30.55965, 30.77884, 30.99778, 31.21648, 31.43492, 31.6531, 31.87103, 
    32.08869, 32.30609, 32.52321, 32.74006, 32.95664, 33.17293, 33.38894, 
    33.60467, 33.8201, 34.03524, 34.25009, 34.46463, 34.67887, 34.89281, 
    35.10644, 35.31975, 35.53275, 35.74544, 35.9578, 36.16984, 36.38155, 
    36.59294, 36.80399, 37.01471, 37.22509, 37.43513, 37.64483, 37.85418, 
    38.06319, 38.27185, 38.48016, 38.68811, 38.8957, 39.10294, 39.30981, 
    39.51632, 39.72246, 39.92824, 40.13364, 40.33868, 40.54333, 40.74762, 
    40.95152, 41.15504, 41.35818, 41.56094, 41.76331, 41.9653, 42.16689, 
    42.36809, 42.5689, 42.76932, 42.96934, 43.16896, 43.36818, 43.567, 
    43.76542, 43.96343, 44.16105, 44.35825, 44.55504, 44.75143, 44.94741, 
    45.14297, 45.33812, 45.53286, 45.72718, 45.92109, 46.11458, 46.30765, 
    46.5003, 46.69254, 46.88435, 47.07573, 47.2667, 47.45724, 47.64736, 
    47.83706, 48.02632, 48.21516, 48.40358, 48.59156, 48.77912, 48.96624, 
    49.15294, 49.33921, 49.52505, 49.71045, 49.89543, 50.07997, 50.26408, 
    50.44776, 50.631, 50.81381, 50.99619, 51.17813, 51.35964, 51.54072, 
    51.72136, 51.90157, 52.08134, 52.26068, 52.43958, 52.61805, 52.79608, 
    52.97368, 53.15084, 53.32757, 53.50386,
  -32.15633, -32.01762, -31.87856, -31.73913, -31.59933, -31.45917, 
    -31.31864, -31.17775, -31.03648, -30.89484, -30.75284, -30.61045, 
    -30.4677, -30.32457, -30.18106, -30.03717, -29.89291, -29.74826, 
    -29.60323, -29.45782, -29.31203, -29.16586, -29.01929, -28.87234, 
    -28.72501, -28.57728, -28.42917, -28.28066, -28.13176, -27.98247, 
    -27.83278, -27.6827, -27.53222, -27.38135, -27.23007, -27.0784, 
    -26.92632, -26.77385, -26.62097, -26.46769, -26.314, -26.15991, 
    -26.00541, -25.85051, -25.6952, -25.53947, -25.38334, -25.2268, 
    -25.06984, -24.91248, -24.75469, -24.5965, -24.43789, -24.27886, 
    -24.11941, -23.95955, -23.79927, -23.63857, -23.47744, -23.3159, 
    -23.15394, -22.99155, -22.82874, -22.66551, -22.50185, -22.33776, 
    -22.17325, -22.00832, -21.84295, -21.67716, -21.51094, -21.34429, 
    -21.17721, -21.0097, -20.84176, -20.67339, -20.50459, -20.33535, 
    -20.16568, -19.99558, -19.82505, -19.65408, -19.48267, -19.31083, 
    -19.13856, -18.96585, -18.79271, -18.61913, -18.44511, -18.27065, 
    -18.09576, -17.92044, -17.74467, -17.56847, -17.39183, -17.21475, 
    -17.03724, -16.85928, -16.68089, -16.50206, -16.32279, -16.14309, 
    -15.96295, -15.78237, -15.60135, -15.41989, -15.238, -15.05567, -14.8729, 
    -14.6897, -14.50606, -14.32198, -14.13747, -13.95252, -13.76713, 
    -13.58132, -13.39506, -13.20838, -13.02126, -12.8337, -12.64572, 
    -12.4573, -12.26845, -12.07917, -11.88946, -11.69932, -11.50876, 
    -11.31776, -11.12634, -10.93449, -10.74222, -10.54952, -10.3564, 
    -10.16286, -9.968895, -9.77451, -9.579706, -9.384483, -9.188843, 
    -8.992786, -8.796316, -8.599431, -8.402134, -8.204426, -8.006309, 
    -7.807782, -7.608849, -7.409511, -7.209768, -7.009623, -6.809076, 
    -6.60813, -6.406787, -6.205048, -6.002913, -5.800387, -5.597469, 
    -5.394162, -5.190468, -4.986389, -4.781926, -4.577082, -4.371858, 
    -4.166256, -3.960279, -3.753929, -3.547208, -3.340117, -3.13266, 
    -2.924839, -2.716655, -2.508111, -2.29921, -2.089954, -1.880345, 
    -1.670386, -1.460079, -1.249427, -1.038433, -0.8270996, -0.6154286, 
    -0.4034232, -0.1910861, 0.02157977, 0.2345717, 0.4478867, 0.661522, 
    0.8754746, 1.089742, 1.30432, 1.519206, 1.734398, 1.949892, 2.165684, 
    2.381773, 2.598153, 2.814823, 3.031779, 3.249017, 3.466535, 3.684328, 
    3.902394, 4.120728, 4.339328, 4.558189, 4.777309, 4.996683, 5.216309, 
    5.436181, 5.656297, 5.876653, 6.097245, 6.318069, 6.539122, 6.760399, 
    6.981897, 7.203612, 7.425539, 7.647676, 7.870017, 8.092559, 8.315297, 
    8.538228, 8.761348, 8.984653, 9.208137, 9.431797, 9.65563, 9.87963, 
    10.10379, 10.32812, 10.55259, 10.77722, 11.00199, 11.22691, 11.45196, 
    11.67715, 11.90246, 12.1279, 12.35346, 12.57913, 12.80492, 13.0308, 
    13.2568, 13.48289, 13.70907, 13.93534, 14.16169, 14.38812, 14.61462, 
    14.8412, 15.06784, 15.29454, 15.5213, 15.7481, 15.97496, 16.20185, 
    16.42879, 16.65575, 16.88274, 17.10976, 17.33679, 17.56384, 17.7909, 
    18.01796, 18.24502, 18.47207, 18.69912, 18.92615, 19.15317, 19.38015, 
    19.60711, 19.83404, 20.06093, 20.28778, 20.51458, 20.74132, 20.96802, 
    21.19464, 21.42121, 21.6477, 21.87412, 22.10046, 22.32672, 22.55289, 
    22.77896, 23.00493, 23.23081, 23.45657, 23.68223, 23.90777, 24.13319, 
    24.35848, 24.58365, 24.80868, 25.03357, 25.25832, 25.48293, 25.70738, 
    25.93168, 26.15582, 26.37979, 26.60359, 26.82723, 27.05068, 27.27396, 
    27.49705, 27.71995, 27.94266, 28.16517, 28.38748, 28.60958, 28.83147, 
    29.05315, 29.27462, 29.49586, 29.71688, 29.93766, 30.15822, 30.37854, 
    30.59862, 30.81845, 31.03803, 31.25737, 31.47645, 31.69527, 31.91383, 
    32.13212, 32.35014, 32.56789, 32.78537, 33.00256, 33.21947, 33.43609, 
    33.65243, 33.86847, 34.08422, 34.29966, 34.5148, 34.72964, 34.94417, 
    35.15839, 35.37229, 35.58588, 35.79914, 36.01208, 36.2247, 36.43698, 
    36.64893, 36.86055, 37.07183, 37.28277, 37.49337, 37.70362, 37.91352, 
    38.12308, 38.33228, 38.54112, 38.74961, 38.95774, 39.1655, 39.3729, 
    39.57993, 39.78659, 39.99289, 40.1988, 40.40435, 40.60951, 40.81429, 
    41.0187, 41.22271, 41.42635, 41.62959, 41.83245, 42.03491, 42.23698, 
    42.43866, 42.63994, 42.84082, 43.04131, 43.24139, 43.44107, 43.64034, 
    43.83921, 44.03767, 44.23573, 44.43337, 44.6306, 44.82742, 45.02383, 
    45.21982, 45.41539, 45.61055, 45.80529, 45.99961, 46.1935, 46.38698, 
    46.58003, 46.77266, 46.96487, 47.15665, 47.348, 47.53893, 47.72943, 
    47.9195, 48.10914, 48.29835, 48.48713, 48.67548, 48.8634, 49.05088, 
    49.23793, 49.42455, 49.61074, 49.79649, 49.9818, 50.16668, 50.35113, 
    50.53513, 50.7187, 50.90184, 51.08454, 51.2668, 51.44862, 51.63001, 
    51.81096, 51.99147, 52.17154, 52.35118, 52.53038, 52.70914, 52.88746, 
    53.06535, 53.24279, 53.4198, 53.59637,
  -32.26381, -32.12504, -31.98591, -31.84641, -31.70655, -31.56632, 
    -31.42573, -31.28476, -31.14342, -31.00171, -30.85962, -30.71716, 
    -30.57433, -30.43111, -30.28752, -30.14355, -29.9992, -29.85446, 
    -29.70935, -29.56384, -29.41796, -29.27169, -29.12503, -28.97798, 
    -28.83054, -28.68271, -28.53449, -28.38587, -28.23687, -28.08746, 
    -27.93766, -27.78746, -27.63687, -27.48587, -27.33448, -27.18268, 
    -27.03048, -26.87788, -26.72487, -26.57146, -26.41763, -26.26341, 
    -26.10877, -25.95373, -25.79827, -25.6424, -25.48612, -25.32943, 
    -25.17232, -25.0148, -24.85686, -24.6985, -24.53973, -24.38054, 
    -24.22092, -24.06089, -23.90044, -23.73956, -23.57827, -23.41654, 
    -23.2544, -23.09183, -22.92883, -22.76541, -22.60156, -22.43728, 
    -22.27257, -22.10744, -21.94187, -21.77587, -21.60945, -21.44258, 
    -21.27529, -21.10757, -20.93941, -20.77082, -20.60179, -20.43233, 
    -20.26243, -20.09209, -19.92132, -19.75012, -19.57847, -19.40639, 
    -19.23387, -19.06091, -18.88751, -18.71367, -18.5394, -18.36468, 
    -18.18953, -18.01393, -17.8379, -17.66142, -17.4845, -17.30714, 
    -17.12934, -16.95111, -16.77242, -16.5933, -16.41374, -16.23374, 
    -16.05329, -15.8724, -15.69108, -15.50931, -15.3271, -15.14445, 
    -14.96136, -14.77783, -14.59386, -14.40946, -14.22461, -14.03932, 
    -13.8536, -13.66743, -13.48083, -13.29379, -13.10632, -12.91841, 
    -12.73006, -12.54128, -12.35206, -12.16241, -11.97232, -11.78181, 
    -11.59086, -11.39948, -11.20767, -11.01543, -10.82276, -10.62966, 
    -10.43614, -10.24219, -10.04781, -9.853013, -9.657791, -9.462148, 
    -9.266084, -9.069599, -8.872697, -8.675378, -8.477643, -8.279492, 
    -8.08093, -7.881955, -7.682569, -7.482775, -7.282573, -7.081964, 
    -6.880952, -6.679536, -6.477719, -6.275503, -6.072888, -5.869877, 
    -5.666472, -5.462675, -5.258486, -5.053908, -4.848944, -4.643595, 
    -4.437862, -4.231749, -4.025257, -3.818388, -3.611145, -3.403529, 
    -3.195543, -2.987189, -2.77847, -2.569387, -2.359943, -2.150141, 
    -1.939983, -1.729472, -1.51861, -1.307399, -1.095843, -0.8839434, 
    -0.6717038, -0.4591264, -0.2462143, -0.03297016, 0.1806032, 0.3945028, 
    0.6087258, 0.8232692, 1.03813, 1.253305, 1.468791, 1.684586, 1.900686, 
    2.117087, 2.333787, 2.550783, 2.76807, 2.985646, 3.203508, 3.421651, 
    3.640074, 3.858771, 4.077739, 4.296976, 4.516477, 4.736239, 4.956258, 
    5.17653, 5.397053, 5.617821, 5.838832, 6.060081, 6.281565, 6.503279, 
    6.725221, 6.947385, 7.169768, 7.392367, 7.615176, 7.838192, 8.061412, 
    8.284829, 8.508442, 8.732245, 8.956235, 9.180407, 9.404756, 9.629279, 
    9.853971, 10.07883, 10.30385, 10.52902, 10.75435, 10.97982, 11.20544, 
    11.4312, 11.65709, 11.88311, 12.10925, 12.33552, 12.5619, 12.7884, 
    13.015, 13.24171, 13.46851, 13.69541, 13.92239, 14.14946, 14.37661, 
    14.60384, 14.83113, 15.05849, 15.28591, 15.51339, 15.74092, 15.9685, 
    16.19612, 16.42377, 16.65146, 16.87918, 17.10692, 17.33467, 17.56245, 
    17.79023, 18.01802, 18.2458, 18.47358, 18.70135, 18.92911, 19.15685, 
    19.38456, 19.61224, 19.83989, 20.0675, 20.29507, 20.5226, 20.75006, 
    20.97748, 21.20483, 21.43211, 21.65932, 21.88646, 22.11352, 22.34049, 
    22.56737, 22.79416, 23.02085, 23.24744, 23.47391, 23.70028, 23.92653, 
    24.15265, 24.37865, 24.60452, 24.83026, 25.05585, 25.28131, 25.50661, 
    25.73176, 25.95675, 26.18158, 26.40625, 26.63074, 26.85507, 27.07921, 
    27.30317, 27.52694, 27.75052, 27.97391, 28.1971, 28.42008, 28.64286, 
    28.86542, 29.08777, 29.3099, 29.53181, 29.75349, 29.97493, 30.19614, 
    30.41712, 30.63785, 30.85833, 31.07856, 31.29854, 31.51826, 31.73772, 
    31.95692, 32.17584, 32.3945, 32.61287, 32.83097, 33.04879, 33.26632, 
    33.48356, 33.70051, 33.91716, 34.13352, 34.34957, 34.56532, 34.78075, 
    34.99588, 35.21069, 35.42518, 35.63935, 35.8532, 36.06672, 36.27991, 
    36.49277, 36.7053, 36.91748, 37.12933, 37.34083, 37.55199, 37.76279, 
    37.97325, 38.18335, 38.3931, 38.60249, 38.81151, 39.02017, 39.22847, 
    39.43639, 39.64395, 39.85114, 40.05795, 40.26438, 40.47043, 40.6761, 
    40.88139, 41.0863, 41.29081, 41.49494, 41.69867, 41.90202, 42.10497, 
    42.30752, 42.50967, 42.71142, 42.91278, 43.11372, 43.31427, 43.5144, 
    43.71413, 43.91346, 44.11237, 44.31086, 44.50895, 44.70662, 44.90387, 
    45.10071, 45.29713, 45.49312, 45.6887, 45.88385, 46.07859, 46.2729, 
    46.46678, 46.66023, 46.85326, 47.04586, 47.23804, 47.42978, 47.62109, 
    47.81197, 48.00242, 48.19244, 48.38202, 48.57117, 48.75988, 48.94816, 
    49.136, 49.32341, 49.51038, 49.69691, 49.883, 50.06866, 50.25388, 
    50.43866, 50.62299, 50.8069, 50.99035, 51.17337, 51.35595, 51.53809, 
    51.71979, 51.90105, 52.08186, 52.26224, 52.44217, 52.62167, 52.80072, 
    52.97933, 53.1575, 53.33523, 53.51252, 53.68937,
  -32.3717, -32.23287, -32.09368, -31.95412, -31.8142, -31.6739, -31.53323, 
    -31.39219, -31.25078, -31.109, -30.96684, -30.8243, -30.68139, -30.53809, 
    -30.39442, -30.25036, -30.10592, -29.9611, -29.8159, -29.6703, -29.52432, 
    -29.37796, -29.2312, -29.08405, -28.93651, -28.78858, -28.64026, 
    -28.49154, -28.34242, -28.19291, -28.04299, -27.89268, -27.74197, 
    -27.59085, -27.43934, -27.28742, -27.13509, -26.98236, -26.82923, 
    -26.67568, -26.52173, -26.36736, -26.21259, -26.05741, -25.90181, 
    -25.74579, -25.58937, -25.43252, -25.27526, -25.11759, -24.95949, 
    -24.80098, -24.64204, -24.48269, -24.32291, -24.16271, -24.00209, 
    -23.84104, -23.67956, -23.51766, -23.35534, -23.19258, -23.0294, 
    -22.86579, -22.70175, -22.53728, -22.37237, -22.20704, -22.04127, 
    -21.87507, -21.70844, -21.54136, -21.37386, -21.20592, -21.03754, 
    -20.86873, -20.69948, -20.52979, -20.35966, -20.1891, -20.01809, 
    -19.84665, -19.67476, -19.50243, -19.32967, -19.15646, -18.98281, 
    -18.80872, -18.63418, -18.4592, -18.28378, -18.10792, -17.93161, 
    -17.75486, -17.57767, -17.40003, -17.22195, -17.04342, -16.86445, 
    -16.68503, -16.50517, -16.32487, -16.14412, -15.96293, -15.7813, 
    -15.59922, -15.41669, -15.23373, -15.05031, -14.86646, -14.68216, 
    -14.49742, -14.31224, -14.12661, -13.94055, -13.75404, -13.56709, 
    -13.3797, -13.19187, -13.0036, -12.81489, -12.62574, -12.43615, 
    -12.24613, -12.05567, -11.86477, -11.67344, -11.48167, -11.28947, 
    -11.09683, -10.90377, -10.71027, -10.51634, -10.32198, -10.1272, 
    -9.931983, -9.736343, -9.540277, -9.343788, -9.146875, -8.94954, 
    -8.751784, -8.55361, -8.355017, -8.156006, -7.956581, -7.756741, 
    -7.556489, -7.355826, -7.154753, -6.953272, -6.751384, -6.549092, 
    -6.346396, -6.1433, -5.939803, -5.735909, -5.531618, -5.326932, 
    -5.121855, -4.916387, -4.71053, -4.504287, -4.29766, -4.09065, -3.88326, 
    -3.675492, -3.467348, -3.258831, -3.049942, -2.840684, -2.63106, 
    -2.421071, -2.210721, -2.000011, -1.788944, -1.577523, -1.365751, 
    -1.153629, -0.9411616, -0.7283502, -0.5151979, -0.3017075, -0.08788192, 
    0.1262761, 0.3407635, 0.5555775, 0.7707149, 0.9861729, 1.201948, 
    1.418038, 1.634439, 1.851148, 2.068162, 2.285478, 2.503091, 2.721, 
    2.9392, 3.157689, 3.376462, 3.595517, 3.814849, 4.034456, 4.254333, 
    4.474478, 4.694886, 4.915554, 5.136478, 5.357655, 5.579079, 5.800749, 
    6.022659, 6.244807, 6.467188, 6.689798, 6.912633, 7.135689, 7.358963, 
    7.58245, 7.806146, 8.030046, 8.254148, 8.478447, 8.702938, 8.927617, 
    9.152481, 9.377523, 9.602742, 9.828132, 10.05369, 10.27941, 10.50528, 
    10.73131, 10.95749, 11.18382, 11.41028, 11.63688, 11.86362, 12.09048, 
    12.31746, 12.54455, 12.77176, 12.99909, 13.22651, 13.45403, 13.68165, 
    13.90936, 14.13715, 14.36502, 14.59297, 14.82099, 15.04908, 15.27722, 
    15.50543, 15.73368, 15.96199, 16.19034, 16.41872, 16.64714, 16.87559, 
    17.10406, 17.33254, 17.56105, 17.78956, 18.01807, 18.24659, 18.4751, 
    18.7036, 18.93209, 19.16055, 19.389, 19.61741, 19.84579, 20.07413, 
    20.30243, 20.53067, 20.75887, 20.98701, 21.21508, 21.44309, 21.67103, 
    21.89889, 22.12667, 22.35436, 22.58197, 22.80947, 23.03688, 23.26418, 
    23.49138, 23.71846, 23.94542, 24.17226, 24.39897, 24.62555, 24.85199, 
    25.07829, 25.30445, 25.53046, 25.75631, 25.982, 26.20753, 26.4329, 
    26.65809, 26.8831, 27.10793, 27.33258, 27.55705, 27.78131, 28.00538, 
    28.22925, 28.45292, 28.67637, 28.89961, 29.12263, 29.34543, 29.568, 
    29.79035, 30.01246, 30.23433, 30.45596, 30.67735, 30.89849, 31.11937, 
    31.34, 31.56036, 31.78047, 32.0003, 32.21986, 32.43915, 32.65816, 
    32.87689, 33.09533, 33.31349, 33.53135, 33.74892, 33.96619, 34.18315, 
    34.39981, 34.61617, 34.8322, 35.04793, 35.26334, 35.47842, 35.69319, 
    35.90762, 36.12173, 36.3355, 36.54894, 36.76204, 36.97479, 37.18721, 
    37.39927, 37.61099, 37.82235, 38.03337, 38.24402, 38.45431, 38.66424, 
    38.87381, 39.08301, 39.29184, 39.5003, 39.70838, 39.91609, 40.12342, 
    40.33037, 40.53694, 40.74312, 40.94891, 41.15432, 41.35934, 41.56396, 
    41.76819, 41.97202, 42.17545, 42.37849, 42.58112, 42.78335, 42.98517, 
    43.18659, 43.3876, 43.58819, 43.78838, 43.98816, 44.18752, 44.38646, 
    44.58498, 44.78309, 44.98078, 45.17805, 45.3749, 45.57132, 45.76732, 
    45.96289, 46.15804, 46.35276, 46.54705, 46.74091, 46.93433, 47.12733, 
    47.3199, 47.51203, 47.70373, 47.89499, 48.08582, 48.27621, 48.46617, 
    48.65569, 48.84476, 49.03341, 49.22161, 49.40937, 49.59669, 49.78357, 
    49.97001, 50.15601, 50.34156, 50.52668, 50.71135, 50.89557, 51.07936, 
    51.2627, 51.44559, 51.62805, 51.81006, 51.99162, 52.17274, 52.35342, 
    52.53366, 52.71344, 52.89279, 53.07169, 53.25014, 53.42816, 53.60572, 
    53.78285,
  -32.48001, -32.34113, -32.20187, -32.06225, -31.92226, -31.7819, -31.64116, 
    -31.50006, -31.35858, -31.21672, -31.07448, -30.93187, -30.78888, 
    -30.6455, -30.50175, -30.35761, -30.21309, -30.06818, -29.92289, 
    -29.7772, -29.63113, -29.48467, -29.33782, -29.19057, -29.04294, 
    -28.8949, -28.74648, -28.59765, -28.44843, -28.2988, -28.14878, 
    -27.99835, -27.84752, -27.69629, -27.54466, -27.39262, -27.24017, 
    -27.08731, -26.93405, -26.78037, -26.62629, -26.47179, -26.31688, 
    -26.16155, -26.00581, -25.84966, -25.69308, -25.53609, -25.37868, 
    -25.22085, -25.0626, -24.90393, -24.74483, -24.58532, -24.42537, 
    -24.26501, -24.10421, -23.94299, -23.78134, -23.61927, -23.45676, 
    -23.29382, -23.13046, -22.96666, -22.80243, -22.63776, -22.47266, 
    -22.30713, -22.14116, -21.97475, -21.80791, -21.64063, -21.47292, 
    -21.30476, -21.13617, -20.96713, -20.79766, -20.62774, -20.45739, 
    -20.28659, -20.11535, -19.94367, -19.77154, -19.59897, -19.42596, 
    -19.2525, -19.0786, -18.90425, -18.72946, -18.55422, -18.37853, -18.2024, 
    -18.02582, -17.8488, -17.67133, -17.49341, -17.31504, -17.13623, 
    -16.95697, -16.77726, -16.59711, -16.4165, -16.23545, -16.05396, 
    -15.87201, -15.68962, -15.50678, -15.32349, -15.13976, -14.95558, 
    -14.77095, -14.58588, -14.40036, -14.2144, -14.02799, -13.84113, 
    -13.65383, -13.46609, -13.2779, -13.08927, -12.9002, -12.71068, 
    -12.52073, -12.33033, -12.13949, -11.94821, -11.7565, -11.56434, 
    -11.37175, -11.17872, -10.98526, -10.79136, -10.59702, -10.40226, 
    -10.20706, -10.01143, -9.815367, -9.618877, -9.421961, -9.224618, 
    -9.026849, -8.828655, -8.630039, -8.431001, -8.231543, -8.031665, 
    -7.831369, -7.630658, -7.429532, -7.227993, -7.026042, -6.82368, 
    -6.620911, -6.417734, -6.214153, -6.010168, -5.805782, -5.600996, 
    -5.395812, -5.190232, -4.984258, -4.777892, -4.571136, -4.363992, 
    -4.156463, -3.948549, -3.740254, -3.531579, -3.322528, -3.113102, 
    -2.903303, -2.693134, -2.482598, -2.271696, -2.060431, -1.848807, 
    -1.636824, -1.424487, -1.211797, -0.9987581, -0.7853718, -0.5716414, 
    -0.3575697, -0.1431594, 0.07158643, 0.286665, 0.5020732, 0.7178082, 
    0.9338668, 1.150246, 1.366943, 1.583954, 1.801276, 2.018906, 2.23684, 
    2.455076, 2.673609, 2.892438, 3.111557, 3.330964, 3.550655, 3.770627, 
    3.990876, 4.211398, 4.43219, 4.653249, 4.874569, 5.096149, 5.317983, 
    5.540069, 5.762402, 5.984978, 6.207793, 6.430845, 6.654128, 6.877638, 
    7.101372, 7.325325, 7.549494, 7.773874, 7.998462, 8.223252, 8.448241, 
    8.673425, 8.898798, 9.124358, 9.3501, 9.576018, 9.80211, 10.02837, 
    10.25479, 10.48138, 10.70812, 10.93501, 11.16204, 11.38922, 11.61654, 
    11.84399, 12.07156, 12.29926, 12.52708, 12.75501, 12.98306, 13.2112, 
    13.43945, 13.66779, 13.89623, 14.12475, 14.35335, 14.58203, 14.81077, 
    15.03959, 15.26847, 15.49741, 15.7264, 15.95543, 16.18451, 16.41363, 
    16.64279, 16.87197, 17.10117, 17.33039, 17.55963, 17.78888, 18.01813, 
    18.24738, 18.47663, 18.70587, 18.93509, 19.16429, 19.39346, 19.62261, 
    19.85172, 20.0808, 20.30983, 20.53881, 20.76774, 20.99661, 21.22541, 
    21.45415, 21.68282, 21.91141, 22.13991, 22.36833, 22.59666, 22.82489, 
    23.05302, 23.28105, 23.50896, 23.73676, 23.96445, 24.192, 24.41943, 
    24.64672, 24.87388, 25.10089, 25.32776, 25.55447, 25.78103, 26.00743, 
    26.23367, 26.45973, 26.68562, 26.91133, 27.13686, 27.36221, 27.58736, 
    27.81232, 28.03708, 28.26163, 28.48598, 28.71012, 28.93403, 29.15773, 
    29.38121, 29.60445, 29.82747, 30.05025, 30.27278, 30.49508, 30.71712, 
    30.93892, 31.16046, 31.38174, 31.60275, 31.8235, 32.04398, 32.26419, 
    32.48412, 32.70376, 32.92312, 33.1422, 33.36098, 33.57946, 33.79765, 
    34.01554, 34.23312, 34.45039, 34.66735, 34.884, 35.10033, 35.31634, 
    35.53202, 35.74738, 35.96241, 36.1771, 36.39146, 36.60547, 36.81915, 
    37.03248, 37.24546, 37.4581, 37.67038, 37.88231, 38.09387, 38.30508, 
    38.51593, 38.7264, 38.93652, 39.14626, 39.35562, 39.56461, 39.77323, 
    39.98146, 40.18932, 40.39679, 40.60387, 40.81056, 41.01686, 41.22278, 
    41.4283, 41.63342, 41.83814, 42.04246, 42.24638, 42.4499, 42.65301, 
    42.85572, 43.05801, 43.2599, 43.46138, 43.66243, 43.86308, 44.06331, 
    44.26312, 44.46251, 44.66148, 44.86003, 45.05816, 45.25586, 45.45314, 
    45.64999, 45.84641, 46.0424, 46.23796, 46.43309, 46.62779, 46.82206, 
    47.01589, 47.20928, 47.40224, 47.59476, 47.78685, 47.9785, 48.16971, 
    48.36047, 48.5508, 48.74069, 48.93014, 49.11914, 49.3077, 49.49582, 
    49.68349, 49.87072, 50.0575, 50.24384, 50.42974, 50.61518, 50.80019, 
    50.98475, 51.16885, 51.35252, 51.53573, 51.7185, 51.90082, 52.0827, 
    52.26412, 52.4451, 52.62563, 52.80572, 52.98536, 53.16455, 53.34329, 
    53.52158, 53.69943, 53.87683,
  -32.58875, -32.4498, -32.31049, -32.17081, -32.03075, -31.89033, -31.74953, 
    -31.60835, -31.4668, -31.32487, -31.18256, -31.03988, -30.89681, 
    -30.75336, -30.60952, -30.4653, -30.3207, -30.1757, -30.03032, -29.88455, 
    -29.73839, -29.59184, -29.44489, -29.29755, -29.14981, -29.00168, 
    -28.85315, -28.70421, -28.55488, -28.40515, -28.25502, -28.10448, 
    -27.95354, -27.80219, -27.65044, -27.49828, -27.34571, -27.19272, 
    -27.03933, -26.88553, -26.73131, -26.57668, -26.42163, -26.26617, 
    -26.11029, -25.95399, -25.79727, -25.64013, -25.48257, -25.32459, 
    -25.16619, -25.00736, -24.8481, -24.68843, -24.52832, -24.36778, 
    -24.20682, -24.04543, -23.88361, -23.72135, -23.55867, -23.39555, 
    -23.232, -23.06801, -22.90359, -22.73873, -22.57344, -22.40771, 
    -22.24154, -22.07493, -21.90788, -21.7404, -21.57247, -21.4041, 
    -21.23529, -21.06603, -20.89634, -20.7262, -20.55561, -20.38458, 
    -20.21311, -20.04119, -19.86882, -19.69601, -19.52275, -19.34904, 
    -19.17489, -19.00028, -18.82523, -18.64973, -18.47378, -18.29738, 
    -18.12053, -17.94324, -17.76549, -17.58729, -17.40864, -17.22954, 
    -17.04999, -16.86999, -16.68954, -16.50864, -16.32728, -16.14548, 
    -15.96323, -15.78052, -15.59737, -15.41376, -15.2297, -15.0452, 
    -14.86024, -14.67484, -14.48898, -14.30268, -14.11592, -13.92872, 
    -13.74107, -13.55297, -13.36443, -13.17544, -12.986, -12.79612, 
    -12.60579, -12.41502, -12.2238, -12.03214, -11.84004, -11.6475, 
    -11.45452, -11.26109, -11.06723, -10.87292, -10.67818, -10.48301, 
    -10.28739, -10.09135, -9.894866, -9.697952, -9.500607, -9.302832, 
    -9.104628, -8.905994, -8.706936, -8.507451, -8.307543, -8.107211, 
    -7.906459, -7.705286, -7.503695, -7.301688, -7.099265, -6.896428, 
    -6.693179, -6.48952, -6.285452, -6.080977, -5.876097, -5.670814, 
    -5.465129, -5.259045, -5.052563, -4.845685, -4.638414, -4.430751, 
    -4.222699, -4.014259, -3.805435, -3.596227, -3.386639, -3.176672, 
    -2.96633, -2.755614, -2.544527, -2.333071, -2.121249, -1.909063, 
    -1.696517, -1.483612, -1.270351, -1.056737, -0.8427727, -0.6284611, 
    -0.4138048, -0.1988066, 0.01653036, 0.2322033, 0.4482092, 0.664545, 
    0.8812077, 1.098194, 1.315501, 1.533126, 1.751064, 1.969314, 2.187871, 
    2.406732, 2.625895, 2.845355, 3.065109, 3.285153, 3.505485, 3.7261, 
    3.946995, 4.168166, 4.38961, 4.611322, 4.8333, 5.05554, 5.278036, 
    5.500786, 5.723787, 5.947033, 6.170521, 6.394247, 6.618207, 6.842397, 
    7.066813, 7.291451, 7.516306, 7.741375, 7.966654, 8.192137, 8.417821, 
    8.643702, 8.869775, 9.096036, 9.32248, 9.549104, 9.775903, 10.00287, 
    10.23001, 10.4573, 10.68476, 10.91236, 11.14011, 11.36801, 11.59605, 
    11.82421, 12.05251, 12.28094, 12.50948, 12.73814, 12.96691, 13.19579, 
    13.42476, 13.65384, 13.883, 14.11226, 14.34159, 14.571, 14.80049, 
    15.03004, 15.25966, 15.48933, 15.71906, 15.94883, 16.17865, 16.40851, 
    16.6384, 16.86832, 17.09827, 17.32823, 17.55821, 17.7882, 18.01819, 
    18.24818, 18.47817, 18.70815, 18.93811, 19.16805, 19.39796, 19.62785, 
    19.8577, 20.08752, 20.31729, 20.547, 20.77667, 21.00628, 21.23582, 
    21.46529, 21.69469, 21.92402, 22.15325, 22.3824, 22.61146, 22.84043, 
    23.06928, 23.29804, 23.52668, 23.7552, 23.98361, 24.21189, 24.44003, 
    24.66805, 24.89592, 25.12365, 25.35123, 25.57866, 25.80593, 26.03304, 
    26.25998, 26.48676, 26.71335, 26.93977, 27.166, 27.39204, 27.61789, 
    27.84354, 28.06899, 28.29424, 28.51928, 28.7441, 28.9687, 29.19308, 
    29.41723, 29.64116, 29.86485, 30.0883, 30.3115, 30.53447, 30.75718, 
    30.97963, 31.20183, 31.42377, 31.64544, 31.86684, 32.08797, 32.30882, 
    32.52939, 32.74967, 32.96967, 33.18938, 33.40879, 33.62791, 33.84672, 
    34.06523, 34.28343, 34.50132, 34.71889, 34.93615, 35.15309, 35.3697, 
    35.58598, 35.80193, 36.01756, 36.23284, 36.44778, 36.66238, 36.87664, 
    37.09055, 37.30411, 37.51731, 37.73016, 37.94265, 38.15478, 38.36654, 
    38.57794, 38.78897, 38.99963, 39.20991, 39.41982, 39.62934, 39.83849, 
    40.04726, 40.25563, 40.46363, 40.67123, 40.87844, 41.08525, 41.29167, 
    41.49769, 41.70331, 41.90853, 42.11335, 42.31776, 42.52176, 42.72536, 
    42.92854, 43.13131, 43.33367, 43.53561, 43.73714, 43.93824, 44.13893, 
    44.33919, 44.53904, 44.73845, 44.93744, 45.13601, 45.33414, 45.53185, 
    45.72913, 45.92598, 46.12239, 46.31837, 46.51391, 46.70902, 46.90369, 
    47.09792, 47.29172, 47.48507, 47.67799, 47.87046, 48.06249, 48.25408, 
    48.44523, 48.63593, 48.82619, 49.016, 49.20536, 49.39429, 49.58276, 
    49.77079, 49.95836, 50.14549, 50.33218, 50.51841, 50.70419, 50.88953, 
    51.07441, 51.25885, 51.44283, 51.62637, 51.80945, 51.99208, 52.17427, 
    52.356, 52.53728, 52.71811, 52.89849, 53.07842, 53.2579, 53.43693, 
    53.61551, 53.79364, 53.97131,
  -32.6979, -32.5589, -32.41953, -32.27979, -32.13968, -31.99919, -31.85832, 
    -31.71708, -31.57546, -31.43346, -31.29108, -31.14832, -31.00517, 
    -30.86165, -30.71773, -30.57343, -30.42875, -30.28367, -30.1382, 
    -29.99234, -29.84609, -29.69945, -29.55241, -29.40497, -29.25714, 
    -29.1089, -28.96027, -28.81124, -28.6618, -28.51196, -28.36172, 
    -28.21107, -28.06002, -27.90856, -27.75669, -27.6044, -27.45171, 
    -27.2986, -27.14509, -26.99116, -26.83681, -26.68204, -26.52686, 
    -26.37126, -26.21524, -26.0588, -25.90194, -25.74465, -25.58695, 
    -25.42881, -25.27025, -25.11127, -24.95186, -24.79202, -24.63175, 
    -24.47105, -24.30992, -24.14835, -23.98636, -23.82393, -23.66106, 
    -23.49776, -23.33403, -23.16986, -23.00525, -22.8402, -22.67471, 
    -22.50878, -22.34241, -22.1756, -22.00835, -21.84065, -21.67252, 
    -21.50393, -21.3349, -21.16543, -20.99551, -20.82515, -20.65434, 
    -20.48307, -20.31137, -20.13921, -19.9666, -19.79355, -19.62004, 
    -19.44608, -19.27168, -19.09682, -18.92151, -18.74575, -18.56953, 
    -18.39287, -18.21575, -18.03818, -17.86015, -17.68167, -17.50274, 
    -17.32336, -17.14352, -16.96322, -16.78247, -16.60127, -16.41962, 
    -16.23751, -16.05494, -15.87193, -15.68845, -15.50453, -15.32015, 
    -15.13532, -14.95003, -14.76429, -14.5781, -14.39146, -14.20436, 
    -14.01681, -13.82881, -13.64036, -13.45146, -13.26211, -13.0723, 
    -12.88205, -12.69135, -12.50021, -12.30861, -12.11657, -11.92408, 
    -11.73115, -11.53777, -11.34395, -11.14968, -10.95498, -10.75983, 
    -10.56424, -10.36821, -10.17175, -9.974845, -9.777506, -9.579731, 
    -9.381522, -9.18288, -8.983808, -8.784305, -8.584372, -8.384011, 
    -8.183225, -7.982013, -7.780378, -7.578321, -7.375843, -7.172946, 
    -6.969632, -6.765902, -6.561758, -6.357202, -6.152235, -5.946859, 
    -5.741076, -5.534888, -5.328297, -5.121305, -4.913913, -4.706124, 
    -4.49794, -4.289363, -4.080395, -3.871038, -3.661295, -3.451168, 
    -3.240659, -3.02977, -2.818504, -2.606863, -2.394851, -2.182468, 
    -1.969719, -1.756605, -1.543129, -1.329294, -1.115102, -0.900557, 
    -0.685661, -0.4704168, -0.2548276, -0.03889617, 0.1773745, 0.3939814, 
    0.6109215, 0.8281917, 1.045789, 1.26371, 1.481951, 1.70051, 1.919383, 
    2.138567, 2.358058, 2.577852, 2.797948, 3.01834, 3.239027, 3.460002, 
    3.681265, 3.90281, 4.124634, 4.346734, 4.569105, 4.791743, 5.014647, 
    5.23781, 5.461229, 5.684901, 5.908822, 6.132987, 6.357392, 6.582034, 
    6.806909, 7.032011, 7.257338, 7.482884, 7.708646, 7.93462, 8.160801, 
    8.387185, 8.613768, 8.840545, 9.067512, 9.294664, 9.521997, 9.749508, 
    9.97719, 10.20504, 10.43305, 10.66123, 10.88955, 11.11803, 11.34665, 
    11.57541, 11.8043, 12.03333, 12.26248, 12.49175, 12.72115, 12.95065, 
    13.18026, 13.40997, 13.63978, 13.86968, 14.09967, 14.32975, 14.5599, 
    14.79013, 15.02042, 15.25078, 15.48119, 15.71166, 15.94218, 16.17275, 
    16.40335, 16.63399, 16.86465, 17.09534, 17.32605, 17.55678, 17.78751, 
    18.01825, 18.24899, 18.47972, 18.71044, 18.94115, 19.17184, 19.4025, 
    19.63313, 19.86373, 20.09428, 20.32479, 20.55526, 20.78567, 21.01601, 
    21.2463, 21.47651, 21.70665, 21.93671, 22.16669, 22.39658, 22.62637, 
    22.85607, 23.08566, 23.31515, 23.54452, 23.77378, 24.00291, 24.23191, 
    24.46079, 24.68953, 24.91813, 25.14658, 25.37488, 25.60303, 25.83101, 
    26.05884, 26.28649, 26.51398, 26.74128, 26.9684, 27.19534, 27.42209, 
    27.64864, 27.87499, 28.10114, 28.32708, 28.55281, 28.77832, 29.00361, 
    29.22868, 29.45352, 29.67812, 29.90249, 30.12662, 30.3505, 30.57413, 
    30.79751, 31.02063, 31.24349, 31.46609, 31.68842, 31.91047, 32.13226, 
    32.35376, 32.57497, 32.7959, 33.01654, 33.23689, 33.45694, 33.67668, 
    33.89613, 34.11526, 34.33408, 34.55259, 34.77078, 34.98865, 35.2062, 
    35.42342, 35.6403, 35.85686, 36.07307, 36.28895, 36.50449, 36.71968, 
    36.93452, 37.14901, 37.36314, 37.57692, 37.79034, 38.0034, 38.21609, 
    38.42841, 38.64037, 38.85195, 39.06315, 39.27398, 39.48443, 39.6945, 
    39.90418, 40.11348, 40.32238, 40.5309, 40.73902, 40.94675, 41.15408, 
    41.361, 41.56753, 41.77365, 41.97937, 42.18468, 42.38959, 42.59408, 
    42.79816, 43.00182, 43.20507, 43.4079, 43.61031, 43.8123, 44.01387, 
    44.21502, 44.41573, 44.61603, 44.81589, 45.01533, 45.21433, 45.4129, 
    45.61105, 45.80875, 46.00602, 46.20285, 46.39925, 46.59521, 46.79073, 
    46.98581, 47.18044, 47.37464, 47.56839, 47.7617, 47.95456, 48.14698, 
    48.33895, 48.53047, 48.72155, 48.91218, 49.10236, 49.29209, 49.48137, 
    49.6702, 49.85858, 50.04651, 50.23399, 50.42101, 50.60758, 50.7937, 
    50.97937, 51.16459, 51.34935, 51.53365, 51.71751, 51.90091, 52.08385, 
    52.26635, 52.44838, 52.62997, 52.8111, 52.99177, 53.17199, 53.35176, 
    53.53107, 53.70994, 53.88834, 54.0663,
  -32.80749, -32.66843, -32.529, -32.3892, -32.24903, -32.10847, -31.96755, 
    -31.82624, -31.68455, -31.54249, -31.40004, -31.2572, -31.11399, 
    -30.97038, -30.82639, -30.68201, -30.53724, -30.39208, -30.24653, 
    -30.10059, -29.95425, -29.80751, -29.66038, -29.51285, -29.36492, 
    -29.21659, -29.06786, -28.91872, -28.76918, -28.61924, -28.46889, 
    -28.31813, -28.16696, -28.01539, -27.8634, -27.711, -27.55819, -27.40496, 
    -27.25131, -27.09726, -26.94278, -26.78788, -26.63257, -26.47683, 
    -26.32067, -26.16409, -26.00709, -25.84966, -25.6918, -25.53352, 
    -25.37481, -25.21567, -25.0561, -24.8961, -24.73566, -24.5748, -24.4135, 
    -24.25177, -24.0896, -23.92699, -23.76395, -23.60047, -23.43655, 
    -23.2722, -23.1074, -22.94216, -22.77648, -22.61035, -22.44378, 
    -22.27677, -22.10932, -21.94141, -21.77306, -21.60427, -21.43502, 
    -21.26533, -21.09519, -20.9246, -20.75356, -20.58207, -20.41013, 
    -20.23773, -20.06489, -19.89159, -19.71784, -19.54363, -19.36898, 
    -19.19386, -19.0183, -18.84227, -18.6658, -18.48886, -18.31147, 
    -18.13363, -17.95533, -17.77657, -17.59735, -17.41768, -17.23755, 
    -17.05696, -16.87592, -16.69442, -16.51246, -16.33004, -16.14717, 
    -15.96384, -15.78005, -15.59581, -15.4111, -15.22594, -15.04033, 
    -14.85425, -14.66773, -14.48074, -14.2933, -14.1054, -13.91705, 
    -13.72825, -13.53899, -13.34927, -13.15911, -12.96849, -12.77741, 
    -12.58589, -12.39392, -12.20149, -12.00862, -11.81529, -11.62152, 
    -11.4273, -11.23264, -11.03752, -10.84197, -10.64597, -10.44952, 
    -10.25264, -10.05531, -9.857543, -9.659337, -9.460693, -9.261614, 
    -9.062099, -8.862149, -8.661767, -8.460954, -8.25971, -8.058038, 
    -7.855938, -7.653413, -7.450463, -7.247091, -7.043297, -6.839084, 
    -6.634453, -6.429407, -6.223946, -6.018072, -5.811788, -5.605094, 
    -5.397994, -5.190489, -4.982581, -4.774272, -4.565564, -4.35646, 
    -4.146961, -3.93707, -3.726788, -3.516119, -3.305064, -3.093626, 
    -2.881808, -2.669611, -2.457039, -2.244093, -2.030777, -1.817093, 
    -1.603043, -1.388631, -1.173858, -0.9587288, -0.7432452, -0.5274101, 
    -0.3112264, -0.09469722, 0.1221746, 0.3393859, 0.5569338, 0.7748149, 
    0.9930263, 1.211565, 1.430427, 1.64961, 1.86911, 2.088923, 2.309048, 
    2.529479, 2.750214, 2.971249, 3.19258, 3.414204, 3.636118, 3.858317, 
    4.080798, 4.303557, 4.526591, 4.749896, 4.973467, 5.197301, 5.421394, 
    5.645742, 5.870342, 6.095188, 6.320277, 6.545605, 6.771168, 6.996962, 
    7.222982, 7.449224, 7.675685, 7.902359, 8.129242, 8.356331, 8.58362, 
    8.811106, 9.038784, 9.266649, 9.494698, 9.722924, 9.951324, 10.1799, 
    10.40863, 10.63753, 10.86658, 11.09578, 11.32513, 11.55462, 11.78424, 
    12.014, 12.24389, 12.4739, 12.70403, 12.93427, 13.16462, 13.39507, 
    13.62562, 13.85627, 14.087, 14.31782, 14.54872, 14.77969, 15.01073, 
    15.24183, 15.473, 15.70422, 15.93549, 16.1668, 16.39815, 16.62954, 
    16.86096, 17.0924, 17.32386, 17.55533, 17.78682, 18.01831, 18.2498, 
    18.48128, 18.71276, 18.94421, 19.17565, 19.40706, 19.63845, 19.86979, 
    20.1011, 20.33236, 20.56357, 20.79473, 21.02582, 21.25685, 21.48781, 
    21.7187, 21.9495, 22.18022, 22.41085, 22.64139, 22.87183, 23.10216, 
    23.33238, 23.56249, 23.79248, 24.02235, 24.25209, 24.48169, 24.71116, 
    24.94049, 25.16967, 25.39869, 25.62756, 25.85627, 26.08482, 26.31319, 
    26.54139, 26.76941, 26.99724, 27.22489, 27.45235, 27.6796, 27.90666, 
    28.13351, 28.36015, 28.58658, 28.81279, 29.03877, 29.26453, 29.49005, 
    29.71534, 29.9404, 30.1652, 30.38976, 30.61407, 30.83812, 31.06192, 
    31.28544, 31.50871, 31.7317, 31.95441, 32.17685, 32.39901, 32.62087, 
    32.84245, 33.06374, 33.28472, 33.50541, 33.72579, 33.94587, 34.16563, 
    34.38508, 34.60421, 34.82302, 35.04151, 35.25967, 35.4775, 35.695, 
    35.91216, 36.12897, 36.34545, 36.56157, 36.77736, 36.99278, 37.20786, 
    37.42257, 37.63692, 37.85092, 38.06454, 38.2778, 38.49069, 38.7032, 
    38.91534, 39.1271, 39.33847, 39.54947, 39.76008, 39.9703, 40.18013, 
    40.38956, 40.59861, 40.80725, 41.0155, 41.22334, 41.43078, 41.63782, 
    41.84444, 42.05067, 42.25647, 42.46187, 42.66685, 42.87141, 43.07556, 
    43.27929, 43.48259, 43.68548, 43.88794, 44.08997, 44.29157, 44.49275, 
    44.69349, 44.89381, 45.09369, 45.29313, 45.49215, 45.69072, 45.88885, 
    46.08655, 46.28381, 46.48063, 46.677, 46.87293, 47.06842, 47.26346, 
    47.45805, 47.6522, 47.8459, 48.03916, 48.23196, 48.42431, 48.61622, 
    48.80767, 48.99867, 49.18922, 49.37931, 49.56895, 49.75814, 49.94688, 
    50.13515, 50.32298, 50.51035, 50.69726, 50.88372, 51.06972, 51.25526, 
    51.44035, 51.62498, 51.80915, 51.99287, 52.17613, 52.35893, 52.54127, 
    52.72316, 52.90459, 53.08556, 53.26608, 53.44613, 53.62573, 53.80487, 
    53.98356, 54.16179,
  -32.9175, -32.77839, -32.63891, -32.49905, -32.35881, -32.2182, -32.07721, 
    -31.93584, -31.79409, -31.65195, -31.50943, -31.36653, -31.22324, 
    -31.07956, -30.93549, -30.79104, -30.64619, -30.50095, -30.35531, 
    -30.20928, -30.06286, -29.91603, -29.76881, -29.62119, -29.47316, 
    -29.32473, -29.1759, -29.02667, -28.87703, -28.72698, -28.57652, 
    -28.42565, -28.27438, -28.12268, -27.97058, -27.81807, -27.66513, 
    -27.51178, -27.35802, -27.20383, -27.04922, -26.8942, -26.73875, 
    -26.58288, -26.42658, -26.26986, -26.11272, -25.95514, -25.79714, 
    -25.63871, -25.47985, -25.32055, -25.16082, -25.00067, -24.84007, 
    -24.67904, -24.51758, -24.35567, -24.19334, -24.03056, -23.86734, 
    -23.70368, -23.53958, -23.37504, -23.21005, -23.04462, -22.87875, 
    -22.71243, -22.54566, -22.37844, -22.21078, -22.04268, -21.87412, 
    -21.70511, -21.53565, -21.36574, -21.19538, -21.02456, -20.85329, 
    -20.68157, -20.5094, -20.33677, -20.16368, -19.99014, -19.81615, 
    -19.6417, -19.46679, -19.29142, -19.11559, -18.93931, -18.76257, 
    -18.58537, -18.40771, -18.22959, -18.05101, -17.87197, -17.69247, 
    -17.51252, -17.3321, -17.15122, -16.96988, -16.78808, -16.60581, 
    -16.42309, -16.23991, -16.05626, -15.87216, -15.68759, -15.50257, 
    -15.31708, -15.13113, -14.94473, -14.75786, -14.57053, -14.38275, 
    -14.19451, -14.0058, -13.81664, -13.62702, -13.43695, -13.24641, 
    -13.05542, -12.86398, -12.67208, -12.47972, -12.28691, -12.09365, 
    -11.89994, -11.70577, -11.51115, -11.31608, -11.12056, -10.9246, 
    -10.72818, -10.53132, -10.33401, -10.13626, -9.938068, -9.73943, 
    -9.540351, -9.340831, -9.140872, -8.940475, -8.739642, -8.538374, 
    -8.336672, -8.134537, -7.931971, -7.728976, -7.525552, -7.321702, 
    -7.117428, -6.91273, -6.707611, -6.502071, -6.296114, -6.08974, 
    -5.882952, -5.675751, -5.46814, -5.26012, -5.051693, -4.842862, 
    -4.633628, -4.423994, -4.213962, -4.003533, -3.792711, -3.581497, 
    -3.369894, -3.157905, -2.945531, -2.732775, -2.51964, -2.306128, 
    -2.092242, -1.877985, -1.663358, -1.448365, -1.233009, -1.017292, 
    -0.8012179, -0.5847886, -0.3680072, -0.1508769, 0.06659938, 0.2844186, 
    0.5025776, 0.7210733, 0.9399025, 1.159062, 1.378549, 1.598359, 1.81849, 
    2.038937, 2.259699, 2.48077, 2.702148, 2.92383, 3.14581, 3.368087, 
    3.590656, 3.813513, 4.036655, 4.260079, 4.48378, 4.707754, 4.931998, 
    5.156507, 5.381278, 5.606307, 5.831589, 6.057121, 6.282898, 6.508918, 
    6.735174, 6.961663, 7.188381, 7.415324, 7.642488, 7.869866, 8.097457, 
    8.325255, 8.553256, 8.781456, 9.00985, 9.238432, 9.4672, 9.696149, 
    9.925273, 10.15457, 10.38403, 10.61366, 10.84344, 11.07337, 11.30345, 
    11.53368, 11.76404, 11.99454, 12.22517, 12.45592, 12.68679, 12.91777, 
    13.14886, 13.38006, 13.61136, 13.84275, 14.07424, 14.3058, 14.53745, 
    14.76917, 15.00097, 15.23283, 15.46474, 15.69672, 15.92874, 16.16081, 
    16.39292, 16.62506, 16.85723, 17.08943, 17.32165, 17.55388, 17.78612, 
    18.01837, 18.25062, 18.48286, 18.71509, 18.9473, 19.1795, 19.41166, 
    19.6438, 19.8759, 20.10797, 20.33998, 20.57195, 20.80385, 21.0357, 
    21.26748, 21.4992, 21.73083, 21.96239, 22.19386, 22.42523, 22.65652, 
    22.8877, 23.11877, 23.34974, 23.58059, 23.81132, 24.04193, 24.27241, 
    24.50275, 24.73295, 24.96301, 25.19292, 25.42268, 25.65228, 25.88171, 
    26.11098, 26.34008, 26.569, 26.79774, 27.02629, 27.25465, 27.48282, 
    27.71079, 27.93856, 28.16611, 28.39346, 28.62059, 28.8475, 29.07418, 
    29.30063, 29.52685, 29.75283, 29.97857, 30.20406, 30.42931, 30.65429, 
    30.87902, 31.10349, 31.32769, 31.55162, 31.77528, 31.99866, 32.22176, 
    32.44457, 32.66709, 32.88932, 33.11126, 33.33289, 33.55422, 33.77524, 
    33.99596, 34.21635, 34.43643, 34.65619, 34.87563, 35.09473, 35.31351, 
    35.53196, 35.75006, 35.96782, 36.18525, 36.40232, 36.61905, 36.83542, 
    37.05144, 37.2671, 37.4824, 37.69733, 37.9119, 38.1261, 38.33993, 
    38.55338, 38.76646, 38.97915, 39.19146, 39.40339, 39.61493, 39.82608, 
    40.03685, 40.24721, 40.45718, 40.66675, 40.87592, 41.08469, 41.29305, 
    41.50101, 41.70855, 41.91569, 42.12241, 42.32872, 42.53461, 42.74009, 
    42.94514, 43.14977, 43.35398, 43.55776, 43.76112, 43.96404, 44.16654, 
    44.36861, 44.57024, 44.77144, 44.9722, 45.17253, 45.37242, 45.57187, 
    45.77088, 45.96945, 46.16758, 46.36526, 46.56249, 46.75928, 46.95563, 
    47.15152, 47.34697, 47.54197, 47.73652, 47.93061, 48.12425, 48.31744, 
    48.51018, 48.70247, 48.89429, 49.08567, 49.27658, 49.46704, 49.65705, 
    49.8466, 50.03568, 50.22431, 50.41248, 50.6002, 50.78745, 50.97424, 
    51.16058, 51.34645, 51.53186, 51.71682, 51.90131, 52.08534, 52.26892, 
    52.45203, 52.63467, 52.81686, 52.99859, 53.17986, 53.36067, 53.54101, 
    53.7209, 53.90033, 54.07929, 54.2578,
  -33.02795, -32.88878, -32.74924, -32.60933, -32.46904, -32.32837, 
    -32.18731, -32.04588, -31.90406, -31.76186, -31.61928, -31.4763, 
    -31.33294, -31.18919, -31.04505, -30.90051, -30.75559, -30.61027, 
    -30.46455, -30.31844, -30.17192, -30.02501, -29.8777, -29.72998, 
    -29.58187, -29.43334, -29.28441, -29.13508, -28.98534, -28.83518, 
    -28.68462, -28.53365, -28.38226, -28.23046, -28.07824, -27.92561, 
    -27.77256, -27.61909, -27.4652, -27.31089, -27.15615, -27.001, -26.84542, 
    -26.68941, -26.53298, -26.37612, -26.21883, -26.06112, -25.90297, 
    -25.74439, -25.58537, -25.42593, -25.26605, -25.10573, -24.94497, 
    -24.78378, -24.62215, -24.46008, -24.29757, -24.13462, -23.97122, 
    -23.80739, -23.6431, -23.47838, -23.3132, -23.14758, -22.98152, -22.815, 
    -22.64804, -22.48063, -22.31276, -22.14445, -21.97568, -21.80646, 
    -21.63678, -21.46666, -21.29607, -21.12504, -20.95354, -20.78159, 
    -20.60918, -20.43632, -20.263, -20.08921, -19.91497, -19.74027, 
    -19.56511, -19.38949, -19.21341, -19.03687, -18.85986, -18.68239, 
    -18.50446, -18.32607, -18.14721, -17.9679, -17.78811, -17.60787, 
    -17.42716, -17.24599, -17.06435, -16.88225, -16.69969, -16.51666, 
    -16.33316, -16.14921, -15.96478, -15.7799, -15.59455, -15.40873, 
    -15.22246, -15.03572, -14.84851, -14.66084, -14.47271, -14.28412, 
    -14.09507, -13.90555, -13.71557, -13.52513, -13.33423, -13.14287, 
    -12.95105, -12.75877, -12.56604, -12.37284, -12.17919, -11.98509, 
    -11.79052, -11.5955, -11.40003, -11.20411, -11.00773, -10.8109, 
    -10.61362, -10.41589, -10.21771, -10.01909, -9.820015, -9.620499, 
    -9.420537, -9.220134, -9.019288, -8.818002, -8.616277, -8.414115, 
    -8.211515, -8.008482, -7.805015, -7.601116, -7.396787, -7.192029, 
    -6.986845, -6.781234, -6.5752, -6.368744, -6.161869, -5.954575, 
    -5.746864, -5.53874, -5.330203, -5.121255, -4.911899, -4.702137, 
    -4.49197, -4.281402, -4.070433, -3.859068, -3.647307, -3.435153, 
    -3.222609, -3.009677, -2.79636, -2.582659, -2.368578, -2.154119, 
    -1.939285, -1.724079, -1.508502, -1.292559, -1.076252, -0.8595835, 
    -0.6425565, -0.4251742, -0.2074394, 0.01064482, 0.2290754, 0.4478491, 
    0.6669629, 0.8864136, 1.106198, 1.326312, 1.546754, 1.767519, 1.988605, 
    2.210007, 2.431723, 2.653748, 2.876079, 3.098714, 3.321647, 3.544875, 
    3.768395, 3.992203, 4.216294, 4.440666, 4.665314, 4.890235, 5.115424, 
    5.340877, 5.566591, 5.792561, 6.018783, 6.245254, 6.471968, 6.698922, 
    6.926112, 7.153533, 7.381181, 7.609052, 7.837141, 8.065444, 8.293956, 
    8.522674, 8.751592, 8.980706, 9.210011, 9.439505, 9.669179, 9.899032, 
    10.12906, 10.35925, 10.58961, 10.82013, 11.0508, 11.28162, 11.51259, 
    11.74369, 11.97493, 12.2063, 12.4378, 12.66942, 12.90115, 13.13299, 
    13.36494, 13.59699, 13.82914, 14.06138, 14.2937, 14.5261, 14.75858, 
    14.99113, 15.22375, 15.45643, 15.68916, 15.92194, 16.15477, 16.38764, 
    16.62055, 16.85348, 17.08644, 17.31942, 17.55242, 17.78542, 18.01843, 
    18.25144, 18.48444, 18.71743, 18.95041, 19.18337, 19.4163, 19.6492, 
    19.88206, 20.11488, 20.34766, 20.58038, 20.81305, 21.04566, 21.2782, 
    21.51066, 21.74306, 21.97536, 22.20759, 22.43972, 22.67175, 22.90369, 
    23.13551, 23.36723, 23.59883, 23.8303, 24.06166, 24.29287, 24.52396, 
    24.7549, 24.9857, 25.21635, 25.44684, 25.67717, 25.90734, 26.13734, 
    26.36716, 26.59681, 26.82627, 27.05555, 27.28463, 27.51352, 27.7422, 
    27.97068, 28.19895, 28.42701, 28.65484, 28.88246, 29.10984, 29.33699, 
    29.56391, 29.79059, 30.01702, 30.2432, 30.46913, 30.6948, 30.92022, 
    31.14536, 31.37024, 31.59484, 31.81917, 32.04322, 32.26698, 32.49046, 
    32.71364, 32.93652, 33.15911, 33.38139, 33.60337, 33.82504, 34.04639, 
    34.26742, 34.48814, 34.70853, 34.92859, 35.14832, 35.36772, 35.58678, 
    35.8055, 36.02388, 36.24191, 36.45958, 36.67691, 36.89388, 37.11049, 
    37.32674, 37.54263, 37.75814, 37.97329, 38.18807, 38.40247, 38.61649, 
    38.83013, 39.04338, 39.25626, 39.46874, 39.68083, 39.89253, 40.10383, 
    40.31474, 40.52524, 40.73534, 40.94504, 41.15434, 41.36322, 41.57169, 
    41.77975, 41.98739, 42.19462, 42.40143, 42.60782, 42.81379, 43.01933, 
    43.22445, 43.42914, 43.6334, 43.83723, 44.04063, 44.24359, 44.44612, 
    44.64822, 44.84987, 45.05109, 45.25186, 45.4522, 45.65209, 45.85154, 
    46.05054, 46.24909, 46.4472, 46.64486, 46.84206, 47.03882, 47.23513, 
    47.43098, 47.62638, 47.82133, 48.01582, 48.20985, 48.40343, 48.59656, 
    48.78922, 48.98143, 49.17317, 49.36446, 49.55529, 49.74565, 49.93556, 
    50.125, 50.31398, 50.5025, 50.69056, 50.87815, 51.06528, 51.25195, 
    51.43816, 51.6239, 51.80917, 51.99399, 52.17834, 52.36222, 52.54564, 
    52.7286, 52.91109, 53.09311, 53.27468, 53.45578, 53.63641, 53.81659, 
    53.99629, 54.17554, 54.35432,
  -33.13883, -32.99961, -32.86002, -32.72005, -32.5797, -32.43897, -32.29786, 
    -32.15636, -32.01448, -31.87222, -31.72956, -31.58652, -31.44309, 
    -31.29927, -31.15505, -31.01044, -30.86544, -30.72004, -30.57424, 
    -30.42805, -30.28145, -30.13445, -29.98705, -29.83924, -29.69104, 
    -29.54242, -29.39339, -29.24396, -29.09412, -28.94386, -28.7932, 
    -28.64211, -28.49062, -28.33871, -28.18638, -28.03363, -27.88046, 
    -27.72687, -27.57286, -27.41843, -27.26357, -27.10828, -26.95257, 
    -26.79643, -26.63987, -26.48287, -26.32544, -26.16758, -26.00929, 
    -25.85056, -25.6914, -25.5318, -25.37176, -25.21129, -25.05037, 
    -24.88902, -24.72723, -24.56499, -24.40231, -24.23918, -24.07561, 
    -23.9116, -23.74714, -23.58223, -23.41687, -23.25106, -23.0848, 
    -22.91809, -22.75093, -22.58332, -22.41525, -22.24673, -22.07775, 
    -21.90832, -21.73843, -21.56809, -21.39729, -21.22602, -21.0543, 
    -20.88213, -20.70949, -20.53639, -20.36283, -20.1888, -20.01432, 
    -19.83937, -19.66396, -19.48808, -19.31174, -19.13494, -18.95767, 
    -18.77994, -18.60174, -18.42307, -18.24394, -18.06434, -17.88428, 
    -17.70375, -17.52275, -17.34128, -17.15935, -16.97695, -16.79408, 
    -16.61074, -16.42694, -16.24267, -16.05793, -15.87272, -15.68705, 
    -15.50091, -15.3143, -15.12722, -14.93968, -14.75167, -14.5632, 
    -14.37425, -14.18484, -13.99497, -13.80463, -13.61383, -13.42256, 
    -13.23083, -13.03864, -12.84598, -12.65286, -12.45928, -12.26524, 
    -12.07074, -11.87578, -11.68036, -11.48449, -11.28815, -11.09136, 
    -10.89412, -10.69642, -10.49827, -10.29966, -10.1006, -9.901096, 
    -9.70114, -9.500737, -9.299887, -9.098591, -8.896851, -8.694668, 
    -8.492043, -8.288979, -8.085476, -7.881535, -7.677159, -7.472349, 
    -7.267106, -7.061432, -6.855329, -6.648798, -6.441843, -6.234462, 
    -6.02666, -5.818438, -5.609797, -5.400741, -5.19127, -4.981387, 
    -4.771093, -4.560392, -4.349285, -4.137774, -3.925863, -3.713552, 
    -3.500845, -3.287744, -3.074251, -2.860368, -2.6461, -2.431447, 
    -2.216412, -2.000999, -1.785209, -1.569046, -1.352513, -1.135612, 
    -0.9183462, -0.7007183, -0.4827316, -0.2643889, -0.04569335, 0.173352, 
    0.392744, 0.6124794, 0.8325552, 1.052968, 1.273714, 1.494791, 1.716195, 
    1.937922, 2.159969, 2.382332, 2.605009, 2.827995, 3.051286, 3.27488, 
    3.498772, 3.722959, 3.947436, 4.1722, 4.397247, 4.622574, 4.848176, 
    5.074049, 5.300189, 5.526592, 5.753254, 5.980171, 6.207339, 6.434753, 
    6.66241, 6.890306, 7.118434, 7.346792, 7.575375, 7.804179, 8.033198, 
    8.26243, 8.491869, 8.721511, 8.951351, 9.181384, 9.411607, 9.642014, 
    9.8726, 10.10336, 10.33429, 10.56539, 10.79665, 11.02806, 11.25963, 
    11.49134, 11.72319, 11.95518, 12.1873, 12.41955, 12.65192, 12.88441, 
    13.11701, 13.34971, 13.58252, 13.81543, 14.04842, 14.28151, 14.51467, 
    14.74791, 14.98123, 15.21461, 15.44805, 15.68155, 15.9151, 16.14869, 
    16.38233, 16.616, 16.8497, 17.08343, 17.31718, 17.55094, 17.78471, 
    18.01849, 18.25227, 18.48604, 18.7198, 18.95354, 19.18727, 19.42097, 
    19.65463, 19.88826, 20.12185, 20.35539, 20.58888, 20.82231, 21.05568, 
    21.28898, 21.52221, 21.75537, 21.98844, 22.22142, 22.45431, 22.6871, 
    22.91979, 23.15237, 23.38484, 23.61719, 23.84942, 24.08152, 24.31349, 
    24.54532, 24.77701, 25.00855, 25.23994, 25.47118, 25.70225, 25.93315, 
    26.16389, 26.39445, 26.62482, 26.85502, 27.08502, 27.31483, 27.54444, 
    27.77384, 28.00304, 28.23203, 28.4608, 28.68935, 28.91767, 29.14576, 
    29.37362, 29.60124, 29.82861, 30.05574, 30.28262, 30.50924, 30.7356, 
    30.9617, 31.18753, 31.41309, 31.63837, 31.86337, 32.08809, 32.31252, 
    32.53666, 32.76051, 32.98405, 33.2073, 33.43024, 33.65286, 33.87518, 
    34.09717, 34.31885, 34.5402, 34.76123, 34.98192, 35.20228, 35.4223, 
    35.64198, 35.86132, 36.08031, 36.29895, 36.51724, 36.73517, 36.95274, 
    37.16994, 37.38679, 37.60326, 37.81937, 38.0351, 38.25045, 38.46543, 
    38.68002, 38.89423, 39.10805, 39.32148, 39.53452, 39.74716, 39.95941, 
    40.17126, 40.38271, 40.59375, 40.80439, 41.01461, 41.22443, 41.43384, 
    41.64283, 41.8514, 42.05956, 42.2673, 42.47461, 42.6815, 42.88796, 
    43.09399, 43.2996, 43.50478, 43.70952, 43.91383, 44.11769, 44.32113, 
    44.52412, 44.72668, 44.92879, 45.13046, 45.33169, 45.53247, 45.7328, 
    45.93269, 46.13212, 46.3311, 46.52964, 46.72772, 46.92535, 47.12252, 
    47.31924, 47.5155, 47.71131, 47.90665, 48.10154, 48.29597, 48.48994, 
    48.68344, 48.87649, 49.06907, 49.26119, 49.45285, 49.64404, 49.83477, 
    50.02504, 50.21484, 50.40417, 50.59304, 50.78144, 50.96938, 51.15685, 
    51.34385, 51.53038, 51.71645, 51.90205, 52.08718, 52.27185, 52.45605, 
    52.63977, 52.82304, 53.00583, 53.18816, 53.37002, 53.55141, 53.73233, 
    53.91279, 54.09278, 54.27231, 54.45136,
  -33.25014, -33.11088, -32.97123, -32.83121, -32.6908, -32.55002, -32.40885, 
    -32.26729, -32.12535, -31.98302, -31.84031, -31.6972, -31.5537, -31.4098, 
    -31.26552, -31.12083, -30.97575, -30.83028, -30.6844, -30.53812, 
    -30.39144, -30.24436, -30.09687, -29.94897, -29.80067, -29.65196, 
    -29.50284, -29.35331, -29.20337, -29.05302, -28.90225, -28.75106, 
    -28.59945, -28.44743, -28.29499, -28.14213, -27.98885, -27.83514, 
    -27.68101, -27.52645, -27.37147, -27.21606, -27.06022, -26.90395, 
    -26.74724, -26.59011, -26.43254, -26.27454, -26.11611, -25.95723, 
    -25.79792, -25.63817, -25.47798, -25.31735, -25.15628, -24.99476, 
    -24.8328, -24.6704, -24.50755, -24.34425, -24.18051, -24.01632, 
    -23.85168, -23.68658, -23.52104, -23.35504, -23.18859, -23.02169, 
    -22.85434, -22.68652, -22.51825, -22.34953, -22.18034, -22.0107, 
    -21.8406, -21.67004, -21.49902, -21.32753, -21.15559, -20.98318, 
    -20.81031, -20.63697, -20.46317, -20.28891, -20.11418, -19.93899, 
    -19.76332, -19.5872, -19.4106, -19.23354, -19.05601, -18.87801, 
    -18.69954, -18.5206, -18.34119, -18.16131, -17.98096, -17.80015, 
    -17.61886, -17.4371, -17.25487, -17.07217, -16.889, -16.70536, -16.52124, 
    -16.33666, -16.1516, -15.96607, -15.78008, -15.59361, -15.40666, 
    -15.21925, -15.03137, -14.84302, -14.6542, -14.46491, -14.27515, 
    -14.08492, -13.89422, -13.70305, -13.51142, -13.31931, -13.12675, 
    -12.93371, -12.74021, -12.54624, -12.35181, -12.15691, -11.96156, 
    -11.76574, -11.56945, -11.37271, -11.17551, -10.97784, -10.77972, 
    -10.58115, -10.38211, -10.18262, -9.982679, -9.782284, -9.581436, 
    -9.380137, -9.17839, -8.976193, -8.773551, -8.570463, -8.366931, 
    -8.162956, -7.95854, -7.753685, -7.548392, -7.342662, -7.136497, -6.9299, 
    -6.722871, -6.515412, -6.307526, -6.099214, -5.890477, -5.681319, 
    -5.47174, -5.261744, -5.051331, -4.840504, -4.629265, -4.417617, 
    -4.205562, -3.993102, -3.780239, -3.566975, -3.353314, -3.139257, 
    -2.924807, -2.709967, -2.494739, -2.279125, -2.06313, -1.846754, 
    -1.630002, -1.412875, -1.195377, -0.9775104, -0.7592784, -0.5406838, 
    -0.3217298, -0.1024194, 0.1172443, 0.3372582, 0.5576189, 0.7783234, 
    0.9993681, 1.22075, 1.442466, 1.664511, 1.886884, 2.10958, 2.332595, 
    2.555927, 2.779571, 3.003525, 3.227783, 3.452343, 3.6772, 3.902351, 
    4.127792, 4.353519, 4.579529, 4.805816, 5.032377, 5.259209, 5.486306, 
    5.713665, 5.941282, 6.169152, 6.397271, 6.625636, 6.85424, 7.083081, 
    7.312154, 7.541454, 7.770978, 8.00072, 8.230676, 8.460841, 8.691212, 
    8.921782, 9.152549, 9.383506, 9.61465, 9.845975, 10.07748, 10.30915, 
    10.54099, 10.773, 11.00516, 11.23747, 11.46994, 11.70254, 11.93529, 
    12.16816, 12.40117, 12.6343, 12.86755, 13.1009, 13.33437, 13.56794, 
    13.80161, 14.03537, 14.26922, 14.50316, 14.73717, 14.97125, 15.2054, 
    15.43961, 15.67388, 15.9082, 16.14257, 16.37697, 16.61142, 16.84589, 
    17.08039, 17.31492, 17.54945, 17.784, 18.01855, 18.2531, 18.48765, 
    18.72218, 18.9567, 19.1912, 19.42567, 19.66011, 19.89451, 20.12887, 
    20.36318, 20.59744, 20.83164, 21.06578, 21.29985, 21.53385, 21.76777, 
    22.00161, 22.23536, 22.46901, 22.70257, 22.93602, 23.16936, 23.40259, 
    23.6357, 23.86868, 24.10154, 24.33426, 24.56684, 24.79928, 25.03157, 
    25.26371, 25.49569, 25.72751, 25.95915, 26.19063, 26.42193, 26.65304, 
    26.88397, 27.1147, 27.34524, 27.57558, 27.80571, 28.03564, 28.26534, 
    28.49483, 28.7241, 28.95313, 29.18194, 29.4105, 29.63883, 29.86691, 
    30.09474, 30.32232, 30.54963, 30.77669, 31.00348, 31.23, 31.45624, 
    31.68221, 31.90789, 32.13328, 32.35839, 32.5832, 32.80771, 33.03192, 
    33.25583, 33.47942, 33.7027, 33.92567, 34.14831, 34.37064, 34.59263, 
    34.81429, 35.03562, 35.25661, 35.47726, 35.69757, 35.91753, 36.13713, 
    36.35639, 36.57529, 36.79382, 37.012, 37.2298, 37.44725, 37.66431, 
    37.88101, 38.09732, 38.31326, 38.52881, 38.74398, 38.95876, 39.17315, 
    39.38714, 39.60073, 39.81394, 40.02674, 40.23913, 40.45112, 40.66271, 
    40.87388, 41.08464, 41.29499, 41.50492, 41.71443, 41.92352, 42.13219, 
    42.34044, 42.54826, 42.75565, 42.96261, 43.16914, 43.37523, 43.58089, 
    43.78612, 43.99091, 44.19525, 44.39915, 44.60262, 44.80564, 45.00821, 
    45.21033, 45.41201, 45.61324, 45.81401, 46.01434, 46.21421, 46.41363, 
    46.61259, 46.81109, 47.00914, 47.20673, 47.40386, 47.60053, 47.79674, 
    47.99249, 48.18777, 48.3826, 48.57695, 48.77085, 48.96428, 49.15724, 
    49.34973, 49.54176, 49.73332, 49.92442, 50.11504, 50.30519, 50.49488, 
    50.6841, 50.87285, 51.06112, 51.24893, 51.43627, 51.62313, 51.80953, 
    51.99545, 52.1809, 52.36589, 52.5504, 52.73444, 52.918, 53.1011, 
    53.28373, 53.46589, 53.64757, 53.82878, 54.00953, 54.1898, 54.3696, 
    54.54893,
  -33.3619, -33.22258, -33.08289, -32.94281, -32.80235, -32.66151, -32.52029, 
    -32.37867, -32.23667, -32.09428, -31.9515, -31.80832, -31.66476, 
    -31.52079, -31.37644, -31.23168, -31.08653, -30.94097, -30.79502, 
    -30.64866, -30.5019, -30.35473, -30.20716, -30.05917, -29.91078, 
    -29.76198, -29.61277, -29.46314, -29.3131, -29.16265, -29.01177, 
    -28.86048, -28.70877, -28.55664, -28.40409, -28.25112, -28.09772, 
    -27.9439, -27.78964, -27.63497, -27.47986, -27.32432, -27.16835, 
    -27.01195, -26.85512, -26.69785, -26.54014, -26.382, -26.22342, -26.0644, 
    -25.90495, -25.74504, -25.5847, -25.42392, -25.26269, -25.10101, 
    -24.93889, -24.77632, -24.6133, -24.44983, -24.28592, -24.12155, 
    -23.95673, -23.79145, -23.62573, -23.45954, -23.29291, -23.12581, 
    -22.95826, -22.79025, -22.62178, -22.45285, -22.28345, -22.1136, 
    -21.94329, -21.77251, -21.60127, -21.42957, -21.25739, -21.08476, 
    -20.91166, -20.73809, -20.56405, -20.38955, -20.21458, -20.03913, 
    -19.86322, -19.68684, -19.50999, -19.33267, -19.15487, -18.9766, 
    -18.79787, -18.61866, -18.43897, -18.25881, -18.07818, -17.89708, 
    -17.7155, -17.53345, -17.35093, -17.16792, -16.98445, -16.8005, 
    -16.61608, -16.43118, -16.2458, -16.05995, -15.87363, -15.68683, 
    -15.49956, -15.31182, -15.12359, -14.9349, -14.74573, -14.55609, 
    -14.36598, -14.17539, -13.98433, -13.7928, -13.60079, -13.40832, 
    -13.21537, -13.02196, -12.82807, -12.63372, -12.4389, -12.2436, 
    -12.04785, -11.85162, -11.65493, -11.45778, -11.26016, -11.06208, 
    -10.86354, -10.66454, -10.46507, -10.26515, -10.06477, -9.863932, 
    -9.662638, -9.46089, -9.258689, -9.056036, -8.852932, -8.649379, 
    -8.445377, -8.24093, -8.036036, -7.8307, -7.624922, -7.418704, -7.212047, 
    -7.004952, -6.797422, -6.589459, -6.381064, -6.17224, -5.962987, 
    -5.753308, -5.543205, -5.33268, -5.121736, -4.910373, -4.698595, 
    -4.486403, -4.2738, -4.060789, -3.84737, -3.633548, -3.419323, -3.2047, 
    -2.98968, -2.774265, -2.558459, -2.342264, -2.125683, -1.908718, 
    -1.691373, -1.473649, -1.255551, -1.037081, -0.8182409, -0.5990351, 
    -0.3794664, -0.1595376, 0.06074801, 0.2813873, 0.502377, 0.7237138, 
    0.9453945, 1.167416, 1.389774, 1.612466, 1.835488, 2.058836, 2.282508, 
    2.506499, 2.730806, 2.955425, 3.180352, 3.405584, 3.631116, 3.856946, 
    4.083068, 4.309479, 4.536176, 4.763153, 4.990407, 5.217935, 5.445731, 
    5.673791, 5.902112, 6.130689, 6.359518, 6.588594, 6.817914, 7.047472, 
    7.277265, 7.507287, 7.737535, 7.968004, 8.198689, 8.429586, 8.66069, 
    8.891996, 9.123501, 9.355199, 9.587085, 9.819154, 10.0514, 10.28382, 
    10.51642, 10.74917, 10.98209, 11.21516, 11.44838, 11.68174, 11.91524, 
    12.14888, 12.38265, 12.61654, 12.85055, 13.08468, 13.31892, 13.55326, 
    13.78769, 14.02223, 14.25685, 14.49156, 14.72634, 14.9612, 15.19612, 
    15.43111, 15.66615, 15.90125, 16.13639, 16.37158, 16.6068, 16.84206, 
    17.07734, 17.31264, 17.54795, 17.78328, 18.01861, 18.25394, 18.48927, 
    18.72458, 18.95988, 19.19516, 19.43041, 19.66562, 19.9008, 20.13594, 
    20.37103, 20.60607, 20.84105, 21.07596, 21.3108, 21.54558, 21.78027, 
    22.01488, 22.2494, 22.48382, 22.71814, 22.95236, 23.18647, 23.42046, 
    23.65434, 23.88808, 24.1217, 24.35518, 24.58852, 24.82172, 25.05477, 
    25.28766, 25.52039, 25.75295, 25.98535, 26.21757, 26.44961, 26.68147, 
    26.91313, 27.14461, 27.37588, 27.60695, 27.83782, 28.06847, 28.2989, 
    28.52911, 28.7591, 28.98886, 29.21838, 29.44766, 29.67669, 29.90549, 
    30.13402, 30.3623, 30.59032, 30.81808, 31.04556, 31.27277, 31.4997, 
    31.72635, 31.95272, 32.17879, 32.40458, 32.63007, 32.85525, 33.08013, 
    33.3047, 33.52895, 33.7529, 33.97652, 34.19981, 34.42278, 34.64542, 
    34.86773, 35.08969, 35.31132, 35.5326, 35.75354, 35.97412, 36.19435, 
    36.41422, 36.63374, 36.85288, 37.07166, 37.29008, 37.50811, 37.72578, 
    37.94307, 38.15997, 38.37649, 38.59262, 38.80836, 39.02372, 39.23868, 
    39.45324, 39.6674, 39.88116, 40.09451, 40.30746, 40.52, 40.73212, 
    40.94384, 41.15513, 41.36601, 41.57647, 41.7865, 41.99612, 42.2053, 
    42.41406, 42.62238, 42.83028, 43.03774, 43.24477, 43.45135, 43.6575, 
    43.86321, 44.06848, 44.2733, 44.47768, 44.68161, 44.88509, 45.08812, 
    45.2907, 45.49283, 45.69451, 45.89573, 46.0965, 46.29681, 46.49665, 
    46.69604, 46.89498, 47.09345, 47.29145, 47.489, 47.68608, 47.88269, 
    48.07885, 48.27453, 48.46975, 48.66449, 48.85877, 49.05259, 49.24593, 
    49.4388, 49.6312, 49.82312, 50.01458, 50.20557, 50.39608, 50.58612, 
    50.77569, 50.96478, 51.1534, 51.34155, 51.52922, 51.71641, 51.90314, 
    52.08938, 52.27516, 52.46046, 52.64528, 52.82963, 53.0135, 53.1969, 
    53.37983, 53.56228, 53.74426, 53.92576, 54.10679, 54.28735, 54.46743, 
    54.64703,
  -33.47409, -33.33473, -33.19499, -33.05486, -32.91435, -32.77346, 
    -32.63217, -32.4905, -32.34844, -32.20599, -32.06314, -31.91991, 
    -31.77627, -31.63224, -31.48782, -31.34299, -31.19776, -31.05213, 
    -30.9061, -30.75966, -30.61282, -30.46557, -30.31791, -30.16985, 
    -30.02137, -29.87247, -29.72317, -29.57345, -29.42331, -29.27276, 
    -29.12178, -28.97039, -28.81858, -28.66634, -28.51368, -28.36059, 
    -28.20708, -28.05314, -27.89877, -27.74397, -27.58874, -27.43308, 
    -27.27699, -27.12045, -26.96349, -26.80609, -26.64824, -26.48996, 
    -26.33124, -26.17208, -26.01247, -25.85242, -25.69193, -25.53099, 
    -25.3696, -25.20777, -25.04549, -24.88275, -24.71957, -24.55593, 
    -24.39184, -24.2273, -24.0623, -23.89684, -23.73093, -23.56456, 
    -23.39774, -23.23045, -23.0627, -22.89449, -22.72582, -22.55669, 
    -22.38709, -22.21703, -22.0465, -21.87551, -21.70405, -21.53213, 
    -21.35973, -21.18687, -21.01354, -20.83973, -20.66546, -20.49072, 
    -20.3155, -20.13981, -19.96365, -19.78702, -19.60991, -19.43233, 
    -19.25427, -19.07574, -18.89673, -18.71725, -18.53729, -18.35685, 
    -18.17594, -17.99455, -17.81268, -17.63034, -17.44751, -17.26421, 
    -17.08043, -16.89618, -16.71144, -16.52623, -16.34054, -16.15437, 
    -15.96772, -15.7806, -15.59299, -15.40491, -15.21635, -15.02731, 
    -14.8378, -14.64781, -14.45734, -14.26639, -14.07497, -13.88307, 
    -13.6907, -13.49785, -13.30453, -13.11073, -12.91646, -12.72172, 
    -12.52651, -12.33082, -12.13466, -11.93804, -11.74094, -11.54337, 
    -11.34534, -11.14684, -10.94787, -10.74844, -10.54855, -10.34819, 
    -10.14737, -9.946089, -9.744349, -9.54215, -9.339494, -9.136382, 
    -8.932815, -8.728795, -8.524323, -8.3194, -8.114029, -7.90821, -7.701945, 
    -7.495235, -7.288083, -7.08049, -6.872458, -6.663988, -6.455082, 
    -6.245743, -6.035972, -5.82577, -5.615141, -5.404086, -5.192606, 
    -4.980706, -4.768385, -4.555647, -4.342494, -4.128928, -3.914952, 
    -3.700568, -3.485778, -3.270585, -3.054991, -2.839, -2.622612, -2.405833, 
    -2.188663, -1.971106, -1.753164, -1.534841, -1.316139, -1.097061, 
    -0.8776105, -0.6577901, -0.4376031, -0.2170524, 0.003858696, 0.225127, 
    0.4467493, 0.6687223, 0.8910426, 1.113707, 1.336712, 1.560053, 1.783729, 
    2.007734, 2.232066, 2.45672, 2.681694, 2.906982, 3.132583, 3.358491, 
    3.584703, 3.811215, 4.038023, 4.265122, 4.492511, 4.720183, 4.948134, 
    5.176363, 5.404861, 5.633628, 5.862658, 6.091947, 6.32149, 6.551283, 
    6.781322, 7.011603, 7.24212, 7.47287, 7.703847, 7.935049, 8.166468, 
    8.398102, 8.629945, 8.861992, 9.09424, 9.326683, 9.559316, 9.792135, 
    10.02514, 10.25831, 10.49166, 10.72517, 10.95884, 11.19267, 11.42666, 
    11.66078, 11.89505, 12.12946, 12.36399, 12.59865, 12.83344, 13.06834, 
    13.30335, 13.53846, 13.77367, 14.00898, 14.24438, 14.47987, 14.71543, 
    14.95107, 15.18677, 15.42254, 15.65837, 15.89425, 16.13018, 16.36615, 
    16.60216, 16.83819, 17.07426, 17.31034, 17.54645, 17.78256, 18.01867, 
    18.25479, 18.4909, 18.727, 18.96309, 19.19915, 19.43518, 19.67118, 
    19.90714, 20.14307, 20.37894, 20.61476, 20.85052, 21.08621, 21.32184, 
    21.55739, 21.79286, 22.02824, 22.26354, 22.49874, 22.73384, 22.96883, 
    23.20371, 23.43847, 23.67311, 23.90763, 24.14202, 24.37626, 24.61037, 
    24.84432, 25.07813, 25.31178, 25.54527, 25.77859, 26.01173, 26.24471, 
    26.4775, 26.7101, 26.94251, 27.17473, 27.40674, 27.63855, 27.87015, 
    28.10154, 28.3327, 28.56365, 28.79436, 29.02484, 29.25508, 29.48508, 
    29.71484, 29.94434, 30.17359, 30.40258, 30.6313, 30.85976, 31.08794, 
    31.31585, 31.54348, 31.77082, 31.99787, 32.22464, 32.4511, 32.67727, 
    32.90313, 33.12867, 33.35392, 33.57884, 33.80344, 34.02772, 34.25167, 
    34.4753, 34.69859, 34.92154, 35.14415, 35.36641, 35.58833, 35.8099, 
    36.03111, 36.25196, 36.47246, 36.69258, 36.91235, 37.13174, 37.35076, 
    37.5694, 37.78766, 38.00555, 38.22304, 38.44015, 38.65687, 38.87319, 
    39.08912, 39.30465, 39.51978, 39.73451, 39.94883, 40.16274, 40.37624, 
    40.58932, 40.802, 41.01425, 41.22609, 41.4375, 41.64849, 41.85905, 
    42.06918, 42.27888, 42.48816, 42.69699, 42.9054, 43.11336, 43.32088, 
    43.52796, 43.7346, 43.9408, 44.14655, 44.35184, 44.5567, 44.7611, 
    44.96505, 45.16854, 45.37158, 45.57417, 45.77629, 45.97796, 46.17917, 
    46.37991, 46.5802, 46.78002, 46.97938, 47.17827, 47.3767, 47.57466, 
    47.77215, 47.96917, 48.16572, 48.3618, 48.55742, 48.75256, 48.94722, 
    49.14142, 49.33514, 49.52839, 49.72116, 49.91346, 50.10528, 50.29663, 
    50.4875, 50.67789, 50.86781, 51.05725, 51.24621, 51.43469, 51.6227, 
    51.81023, 51.99728, 52.18385, 52.36995, 52.55556, 52.7407, 52.92536, 
    53.10954, 53.29324, 53.47646, 53.65921, 53.84148, 54.02327, 54.20459, 
    54.38543, 54.56578, 54.74567,
  -33.58673, -33.44733, -33.30753, -33.16736, -33.0268, -32.88585, -32.74451, 
    -32.60279, -32.46067, -32.31816, -32.17525, -32.03195, -31.88825, 
    -31.74416, -31.59966, -31.45477, -31.30947, -31.16376, -31.01766, 
    -30.87114, -30.72422, -30.57689, -30.42915, -30.28099, -30.13243, 
    -29.98345, -29.83405, -29.68424, -29.534, -29.38335, -29.23228, 
    -29.08079, -28.92887, -28.77653, -28.62376, -28.47056, -28.31693, 
    -28.16288, -28.0084, -27.85348, -27.69813, -27.54234, -27.38612, 
    -27.22946, -27.07236, -26.91483, -26.75685, -26.59843, -26.43957, 
    -26.28026, -26.12051, -25.96032, -25.79967, -25.63858, -25.47704, 
    -25.31504, -25.1526, -24.9897, -24.82635, -24.66254, -24.49828, 
    -24.33356, -24.16839, -24.00276, -23.83666, -23.67011, -23.50309, 
    -23.33561, -23.16767, -22.99927, -22.8304, -22.66106, -22.49126, 
    -22.32099, -22.15025, -21.97904, -21.80737, -21.63522, -21.4626, 
    -21.28951, -21.11595, -20.94191, -20.7674, -20.59242, -20.41696, 
    -20.24103, -20.06462, -19.88773, -19.71037, -19.53253, -19.35421, 
    -19.17541, -18.99613, -18.81638, -18.63614, -18.45543, -18.27423, 
    -18.09256, -17.9104, -17.72776, -17.54464, -17.36104, -17.17696, 
    -16.9924, -16.80735, -16.62182, -16.43582, -16.24932, -16.06235, 
    -15.8749, -15.68696, -15.49854, -15.30964, -15.12026, -14.9304, 
    -14.74006, -14.54923, -14.35793, -14.16615, -13.97388, -13.78114, 
    -13.58792, -13.39422, -13.20004, -13.00539, -12.81025, -12.61465, 
    -12.41856, -12.222, -12.02497, -11.82747, -11.62949, -11.43104, 
    -11.23212, -11.03273, -10.83287, -10.63254, -10.43175, -10.23049, 
    -10.02876, -9.826573, -9.623922, -9.42081, -9.217237, -9.013206, 
    -8.808717, -8.603772, -8.398374, -8.192521, -7.986217, -7.779464, 
    -7.572262, -7.364613, -7.156519, -6.947982, -6.739003, -6.529585, 
    -6.319729, -6.109437, -5.89871, -5.687552, -5.475964, -5.263948, 
    -5.051506, -4.838641, -4.625354, -4.411648, -4.197526, -3.982989, 
    -3.76804, -3.552682, -3.336916, -3.120746, -2.904175, -2.687203, 
    -2.469836, -2.252074, -2.033921, -1.81538, -1.596454, -1.377145, 
    -1.157457, -0.9373917, -0.7169532, -0.4961444, -0.2749682, -0.05342805, 
    0.168473, 0.3907316, 0.6133445, 0.8363082, 1.059619, 1.283275, 1.50727, 
    1.731603, 1.956269, 2.181265, 2.406587, 2.632231, 2.858194, 3.084472, 
    3.31106, 3.537956, 3.765155, 3.992653, 4.220446, 4.448531, 4.676902, 
    4.905556, 5.134489, 5.363696, 5.593174, 5.822917, 6.052922, 6.283185, 
    6.5137, 6.744463, 6.975471, 7.206718, 7.4382, 7.669912, 7.90185, 
    8.134009, 8.366385, 8.598972, 8.831766, 9.064762, 9.297956, 9.531342, 
    9.764915, 9.998672, 10.23261, 10.46671, 10.70099, 10.93543, 11.17002, 
    11.40477, 11.63967, 11.87471, 12.10989, 12.3452, 12.58063, 12.81619, 
    13.05187, 13.28766, 13.52355, 13.75955, 13.99564, 14.23182, 14.46809, 
    14.70444, 14.94086, 15.17735, 15.41391, 15.65053, 15.8872, 16.12391, 
    16.36067, 16.59747, 16.8343, 17.07116, 17.30803, 17.54493, 17.78183, 
    18.01874, 18.25565, 18.49255, 18.72944, 18.96631, 19.20317, 19.43999, 
    19.67678, 19.91353, 20.15024, 20.38691, 20.62351, 20.86006, 21.09654, 
    21.33295, 21.56929, 21.80554, 22.04171, 22.27779, 22.51377, 22.74965, 
    22.98542, 23.22108, 23.45662, 23.69203, 23.92732, 24.16248, 24.3975, 
    24.63237, 24.8671, 25.10167, 25.33608, 25.57033, 25.80441, 26.03832, 
    26.27205, 26.50559, 26.73895, 26.97211, 27.20507, 27.43783, 27.67039, 
    27.90273, 28.13485, 28.36676, 28.59843, 28.82988, 29.06109, 29.29206, 
    29.52278, 29.75326, 29.98348, 30.21344, 30.44314, 30.67258, 30.90174, 
    31.13063, 31.35924, 31.58757, 31.81561, 32.04335, 32.27081, 32.49796, 
    32.7248, 32.95134, 33.17757, 33.40348, 33.62908, 33.85435, 34.07929, 
    34.30391, 34.52818, 34.75212, 34.97573, 35.19899, 35.42189, 35.64445, 
    35.86665, 36.0885, 36.30998, 36.5311, 36.75185, 36.97223, 37.19223, 
    37.41186, 37.63111, 37.84998, 38.06845, 38.28654, 38.50425, 38.72155, 
    38.93846, 39.15497, 39.37107, 39.58678, 39.80207, 40.01695, 40.23142, 
    40.44548, 40.65912, 40.87234, 41.08514, 41.29751, 41.50946, 41.72098, 
    41.93207, 42.14273, 42.35295, 42.56274, 42.77209, 42.981, 43.18946, 
    43.39749, 43.60507, 43.8122, 44.01888, 44.22511, 44.43089, 44.63622, 
    44.84109, 45.04551, 45.24947, 45.45297, 45.65601, 45.85859, 46.0607, 
    46.26236, 46.46354, 46.66426, 46.86451, 47.0643, 47.26362, 47.46246, 
    47.66084, 47.85874, 48.05617, 48.25313, 48.44961, 48.64562, 48.84115, 
    49.03621, 49.23079, 49.42489, 49.61852, 49.81166, 50.00433, 50.19651, 
    50.38822, 50.57945, 50.7702, 50.96046, 51.15025, 51.33956, 51.52838, 
    51.71672, 51.90458, 52.09196, 52.27886, 52.46527, 52.6512, 52.83665, 
    53.02163, 53.20611, 53.39012, 53.57364, 53.75668, 53.93925, 54.12133, 
    54.30293, 54.48405, 54.66468, 54.84484,
  -33.69982, -33.56037, -33.42053, -33.28031, -33.1397, -32.9987, -32.85731, 
    -32.71553, -32.57335, -32.43078, -32.28782, -32.14445, -32.00069, 
    -31.85653, -31.71197, -31.56701, -31.42164, -31.27586, -31.12968, 
    -30.98309, -30.83609, -30.68868, -30.54086, -30.39262, -30.24397, 
    -30.0949, -29.94541, -29.79551, -29.64518, -29.49444, -29.34327, 
    -29.19167, -29.03965, -28.8872, -28.73433, -28.58102, -28.42729, 
    -28.27312, -28.11852, -27.96348, -27.80801, -27.6521, -27.49575, 
    -27.33897, -27.18174, -27.02407, -26.86596, -26.70741, -26.54841, 
    -26.38896, -26.22906, -26.06872, -25.90793, -25.74668, -25.58498, 
    -25.42283, -25.26023, -25.09717, -24.93365, -24.76968, -24.60525, 
    -24.44036, -24.27501, -24.10919, -23.94292, -23.77618, -23.60897, 
    -23.44131, -23.27317, -23.10457, -22.9355, -22.76596, -22.59596, 
    -22.42548, -22.25453, -22.08311, -21.91122, -21.73885, -21.56601, 
    -21.39269, -21.2189, -21.04463, -20.86989, -20.69466, -20.51896, 
    -20.34278, -20.16613, -19.98899, -19.81137, -19.63327, -19.45469, 
    -19.27563, -19.09608, -18.91605, -18.73554, -18.55455, -18.37307, 
    -18.19111, -18.00866, -17.82573, -17.64232, -17.45842, -17.27403, 
    -17.08916, -16.9038, -16.71796, -16.53164, -16.34482, -16.15753, 
    -15.96974, -15.78147, -15.59272, -15.40348, -15.21375, -15.02355, 
    -14.83285, -14.64167, -14.45001, -14.25786, -14.06523, -13.87212, 
    -13.67852, -13.48445, -13.28989, -13.09484, -12.89932, -12.70332, 
    -12.50684, -12.30988, -12.11244, -11.91453, -11.71614, -11.51727, 
    -11.31793, -11.11811, -10.91782, -10.71706, -10.51583, -10.31413, 
    -10.11196, -9.909317, -9.706211, -9.502641, -9.298606, -9.094109, 
    -8.889151, -8.683731, -8.477854, -8.27152, -8.06473, -7.857485, 
    -7.649788, -7.441641, -7.233045, -7.024001, -6.814511, -6.604578, 
    -6.394202, -6.183387, -5.972134, -5.760444, -5.548321, -5.335765, 
    -5.12278, -4.909368, -4.695529, -4.481268, -4.266586, -4.051486, 
    -3.83597, -3.62004, -3.403699, -3.18695, -2.969795, -2.752237, -2.534278, 
    -2.315922, -2.09717, -1.878026, -1.658494, -1.438574, -1.218272, 
    -0.9975891, -0.776529, -0.5550948, -0.3332897, -0.1111167, 0.1114208, 
    0.3343194, 0.557576, 0.781187, 1.005149, 1.229459, 1.454112, 1.679106, 
    1.904437, 2.130101, 2.356095, 2.582414, 2.809056, 3.036015, 3.263289, 
    3.490873, 3.718763, 3.946955, 4.175447, 4.404232, 4.633307, 4.862668, 
    5.09231, 5.32223, 5.552423, 5.782886, 6.013612, 6.244598, 6.475841, 
    6.707334, 6.939074, 7.171055, 7.403275, 7.635726, 7.868407, 8.101311, 
    8.334434, 8.56777, 8.801315, 9.035066, 9.269015, 9.50316, 9.737494, 
    9.972013, 10.20671, 10.44158, 10.67663, 10.91184, 11.1472, 11.38273, 
    11.6184, 11.85421, 12.09017, 12.32626, 12.56248, 12.79882, 13.03528, 
    13.27185, 13.50853, 13.74531, 13.98219, 14.21917, 14.45623, 14.69337, 
    14.93058, 15.16786, 15.40522, 15.64263, 15.88009, 16.1176, 16.35516, 
    16.59275, 16.83038, 17.06803, 17.3057, 17.54339, 17.7811, 18.0188, 
    18.25651, 18.49421, 18.73189, 18.96956, 19.20721, 19.44483, 19.68242, 
    19.91997, 20.15748, 20.39493, 20.63233, 20.86967, 21.10695, 21.34415, 
    21.58128, 21.81832, 22.05528, 22.29215, 22.52891, 22.76558, 23.00213, 
    23.23857, 23.4749, 23.7111, 23.94716, 24.1831, 24.41889, 24.65454, 
    24.89004, 25.12538, 25.36056, 25.59558, 25.83043, 26.0651, 26.29959, 
    26.53389, 26.76801, 27.00192, 27.23564, 27.46915, 27.70246, 27.93554, 
    28.16842, 28.40106, 28.63347, 28.86566, 29.0976, 29.3293, 29.56075, 
    29.79196, 30.0229, 30.25359, 30.48401, 30.71416, 30.94403, 31.17363, 
    31.40295, 31.63198, 31.86072, 32.08916, 32.31731, 32.54515, 32.77268, 
    32.99991, 33.22682, 33.45341, 33.67968, 33.90562, 34.13123, 34.35651, 
    34.58145, 34.80605, 35.0303, 35.25421, 35.47776, 35.70096, 35.92381, 
    36.14629, 36.3684, 36.59015, 36.81152, 37.03252, 37.25315, 37.47339, 
    37.69324, 37.91272, 38.1318, 38.35049, 38.56878, 38.78668, 39.00417, 
    39.22126, 39.43795, 39.65422, 39.87009, 40.08554, 40.30058, 40.51519, 
    40.72938, 40.94315, 41.1565, 41.36942, 41.58191, 41.79396, 42.00558, 
    42.21676, 42.42751, 42.63781, 42.84768, 43.0571, 43.26607, 43.4746, 
    43.68267, 43.8903, 44.09747, 44.30419, 44.51045, 44.71626, 44.9216, 
    45.12649, 45.33091, 45.53487, 45.73837, 45.9414, 46.14397, 46.34606, 
    46.54769, 46.74885, 46.94954, 47.14975, 47.34949, 47.54876, 47.74755, 
    47.94587, 48.14371, 48.34107, 48.53795, 48.73436, 48.93028, 49.12573, 
    49.32069, 49.51518, 49.70918, 49.9027, 50.09574, 50.28829, 50.48036, 
    50.67195, 50.86305, 51.05367, 51.2438, 51.43344, 51.62261, 51.81129, 
    51.99948, 52.18719, 52.37441, 52.56114, 52.74739, 52.93316, 53.11843, 
    53.30323, 53.48754, 53.67136, 53.8547, 54.03756, 54.21992, 54.40181, 
    54.58321, 54.76413, 54.94456,
  -33.81335, -33.67386, -33.53398, -33.39371, -33.25305, -33.112, -32.97056, 
    -32.82873, -32.6865, -32.54387, -32.40085, -32.25743, -32.11361, 
    -31.96938, -31.82475, -31.67972, -31.53428, -31.38844, -31.24218, 
    -31.09552, -30.94844, -30.80095, -30.65305, -30.50473, -30.35599, 
    -30.20684, -30.05726, -29.90727, -29.75685, -29.60601, -29.45474, 
    -29.30305, -29.15093, -28.99837, -28.84539, -28.69198, -28.53814, 
    -28.38386, -28.22914, -28.07399, -27.9184, -27.76237, -27.6059, 
    -27.44899, -27.29163, -27.13383, -26.97559, -26.8169, -26.65776, 
    -26.49817, -26.33813, -26.17764, -26.0167, -25.8553, -25.69345, 
    -25.53115, -25.36838, -25.20516, -25.04148, -24.87734, -24.71274, 
    -24.54768, -24.38215, -24.21616, -24.0497, -23.88278, -23.71539, 
    -23.54753, -23.37921, -23.21041, -23.04114, -22.8714, -22.70119, 
    -22.53051, -22.35935, -22.18772, -22.01561, -21.84302, -21.66996, 
    -21.49641, -21.32239, -21.14789, -20.97291, -20.79745, -20.62151, 
    -20.44509, -20.26818, -20.09079, -19.91292, -19.73456, -19.55572, 
    -19.37639, -19.19658, -19.01628, -18.83549, -18.65422, -18.47246, 
    -18.29021, -18.10748, -17.92425, -17.74054, -17.55634, -17.37165, 
    -17.18647, -17.00081, -16.81465, -16.62801, -16.44087, -16.25325, 
    -16.06514, -15.87654, -15.68744, -15.49786, -15.3078, -15.11724, 
    -14.92619, -14.73466, -14.54264, -14.35013, -14.15713, -13.96364, 
    -13.76967, -13.57522, -13.38027, -13.18485, -12.98893, -12.79254, 
    -12.59566, -12.3983, -12.20045, -12.00212, -11.80332, -11.60403, 
    -11.40427, -11.20402, -11.0033, -10.80211, -10.60044, -10.39829, 
    -10.19567, -9.992584, -9.789023, -9.584993, -9.380495, -9.17553, 
    -8.970099, -8.764205, -8.557847, -8.351028, -8.14375, -7.936014, 
    -7.72782, -7.519172, -7.310071, -7.100518, -6.890515, -6.680065, 
    -6.469168, -6.257828, -6.046045, -5.833822, -5.621161, -5.408063, 
    -5.194532, -4.98057, -4.766178, -4.551358, -4.336114, -4.120448, 
    -3.904361, -3.687857, -3.470938, -3.253607, -3.035866, -2.817717, 
    -2.599164, -2.38021, -2.160856, -1.941107, -1.720964, -1.500432, 
    -1.279512, -1.058207, -0.8365222, -0.6144591, -0.3920212, -0.1692118, 
    0.05396578, 0.2775083, 0.5014123, 0.7256745, 0.9502914, 1.175259, 
    1.400575, 1.626235, 1.852234, 2.078571, 2.305241, 2.532239, 2.759563, 
    2.987209, 3.215172, 3.443448, 3.672034, 3.900926, 4.130119, 4.35961, 
    4.589393, 4.819466, 5.049823, 5.28046, 5.511374, 5.742559, 5.974012, 
    6.205728, 6.437702, 6.66993, 6.902407, 7.135128, 7.36809, 7.601287, 
    7.834715, 8.068369, 8.302243, 8.536335, 8.770638, 9.005147, 9.239859, 
    9.474766, 9.709866, 9.945152, 10.18062, 10.41627, 10.65208, 10.88807, 
    11.12421, 11.36051, 11.59697, 11.83356, 12.0703, 12.30718, 12.54418, 
    12.78131, 13.01856, 13.25593, 13.4934, 13.73097, 13.96865, 14.20642, 
    14.44427, 14.68221, 14.92022, 15.1583, 15.39645, 15.63466, 15.87293, 
    16.11124, 16.3496, 16.588, 16.82642, 17.06488, 17.30336, 17.54185, 
    17.78036, 18.01886, 18.25737, 18.49588, 18.73437, 18.97284, 19.21129, 
    19.44972, 19.68811, 19.92646, 20.16476, 20.40302, 20.64122, 20.87936, 
    21.11744, 21.35544, 21.59336, 21.8312, 22.06895, 22.30661, 22.54417, 
    22.78163, 23.01897, 23.25621, 23.49332, 23.7303, 23.96715, 24.20387, 
    24.44045, 24.67688, 24.91315, 25.14927, 25.38523, 25.62102, 25.85664, 
    26.09208, 26.32734, 26.5624, 26.79728, 27.03196, 27.26644, 27.50071, 
    27.73477, 27.96861, 28.20222, 28.43562, 28.66878, 28.9017, 29.13438, 
    29.36682, 29.59901, 29.83094, 30.06262, 30.29403, 30.52517, 30.75604, 
    30.98664, 31.21695, 31.44697, 31.67671, 31.90615, 32.1353, 32.36414, 
    32.59268, 32.82091, 33.04882, 33.27642, 33.50369, 33.73064, 33.95725, 
    34.18354, 34.40948, 34.63509, 34.86035, 35.08526, 35.30982, 35.53403, 
    35.75788, 35.98136, 36.20448, 36.42723, 36.64961, 36.87161, 37.09324, 
    37.31448, 37.53534, 37.75581, 37.97589, 38.19558, 38.41487, 38.63376, 
    38.85225, 39.07034, 39.28801, 39.50528, 39.72213, 39.93857, 40.15459, 
    40.37019, 40.58537, 40.80012, 41.01444, 41.22834, 41.4418, 41.65483, 
    41.86742, 42.07957, 42.29129, 42.50256, 42.71338, 42.92376, 43.1337, 
    43.34318, 43.55221, 43.76078, 43.96891, 44.17657, 44.38377, 44.59052, 
    44.79681, 45.00262, 45.20798, 45.41288, 45.6173, 45.82125, 46.02474, 
    46.22776, 46.4303, 46.63237, 46.83397, 47.03509, 47.23573, 47.4359, 
    47.63559, 47.8348, 48.03353, 48.23178, 48.42955, 48.62683, 48.82364, 
    49.01995, 49.21579, 49.41114, 49.60601, 49.80039, 49.99428, 50.18769, 
    50.38061, 50.57304, 50.76499, 50.95644, 51.14742, 51.33789, 51.52789, 
    51.71739, 51.9064, 52.09492, 52.28296, 52.47051, 52.65756, 52.84413, 
    53.03021, 53.2158, 53.4009, 53.58551, 53.76963, 53.95327, 54.13641, 
    54.31907, 54.50124, 54.68292, 54.86412, 55.04483,
  -33.92735, -33.78781, -33.64788, -33.50757, -33.36686, -33.22577, 
    -33.08427, -32.94239, -32.80011, -32.65743, -32.51435, -32.37087, 
    -32.22699, -32.0827, -31.93801, -31.79291, -31.6474, -31.50149, 
    -31.35516, -31.20843, -31.06127, -30.91371, -30.76573, -30.61732, 
    -30.46851, -30.31927, -30.1696, -30.01952, -29.86901, -29.71807, 
    -29.56671, -29.41492, -29.2627, -29.11005, -28.95696, -28.80344, 
    -28.64949, -28.4951, -28.34027, -28.185, -28.02929, -27.87314, -27.71655, 
    -27.55951, -27.40203, -27.2441, -27.08573, -26.9269, -26.76763, -26.6079, 
    -26.44772, -26.28708, -26.12599, -25.96445, -25.80245, -25.63998, 
    -25.47706, -25.31368, -25.14984, -24.98553, -24.82076, -24.65553, 
    -24.48983, -24.32366, -24.15702, -23.98992, -23.82234, -23.6543, 
    -23.48578, -23.31679, -23.14732, -22.97738, -22.80697, -22.63608, 
    -22.46471, -22.29286, -22.12054, -21.94773, -21.77445, -21.60068, 
    -21.42643, -21.2517, -21.07649, -20.90079, -20.72461, -20.54794, 
    -20.37078, -20.19314, -20.01501, -19.8364, -19.6573, -19.4777, -19.29762, 
    -19.11705, -18.93599, -18.75444, -18.5724, -18.38987, -18.20684, 
    -18.02333, -17.83932, -17.65482, -17.46983, -17.28434, -17.09837, 
    -16.9119, -16.72493, -16.53748, -16.34953, -16.16109, -15.97215, 
    -15.78272, -15.5928, -15.40239, -15.21148, -15.02009, -14.82819, 
    -14.63581, -14.44294, -14.24957, -14.05572, -13.86137, -13.66653, 
    -13.47121, -13.27539, -13.07909, -12.8823, -12.68502, -12.48725, -12.289, 
    -12.09026, -11.89104, -11.69133, -11.49115, -11.29047, -11.08932, 
    -10.88769, -10.68558, -10.48299, -10.27992, -10.07638, -9.872363, 
    -9.667872, -9.462909, -9.257474, -9.05157, -8.845198, -8.638359, 
    -8.431054, -8.223286, -8.015055, -7.806363, -7.597212, -7.387604, 
    -7.17754, -6.967022, -6.756052, -6.544632, -6.332764, -6.120449, 
    -5.90769, -5.694489, -5.480847, -5.266768, -5.052253, -4.837304, 
    -4.621924, -4.406115, -4.18988, -3.97322, -3.756139, -3.538639, 
    -3.320722, -3.102392, -2.88365, -2.6645, -2.444944, -2.224986, -2.004627, 
    -1.783871, -1.562721, -1.34118, -1.119251, -0.8969374, -0.6742418, 
    -0.4511676, -0.2277181, -0.003896533, 0.2202936, 0.4448491, 0.6697663, 
    0.8950419, 1.120672, 1.346654, 1.572983, 1.799656, 2.026669, 2.254019, 
    2.481701, 2.709712, 2.938048, 3.166705, 3.395679, 3.624965, 3.85456, 
    4.08446, 4.314661, 4.545158, 4.775947, 5.007023, 5.238383, 5.470022, 
    5.701936, 5.93412, 6.16657, 6.399281, 6.632248, 6.865468, 7.098934, 
    7.332644, 7.566591, 7.800772, 8.035181, 8.269814, 8.504664, 8.73973, 
    8.975004, 9.210483, 9.446159, 9.682031, 9.918091, 10.15433, 10.39076, 
    10.62735, 10.86412, 11.10105, 11.33813, 11.57537, 11.81276, 12.05029, 
    12.28795, 12.52575, 12.76367, 13.00172, 13.23988, 13.47815, 13.71652, 
    13.955, 14.19357, 14.43222, 14.67096, 14.90978, 15.14867, 15.38762, 
    15.62664, 15.86571, 16.10483, 16.344, 16.5832, 16.82244, 17.06171, 
    17.30099, 17.5403, 17.77961, 18.01893, 18.25825, 18.49756, 18.73686, 
    18.97614, 19.2154, 19.45464, 19.69383, 19.93299, 20.17211, 20.41117, 
    20.65018, 20.88912, 21.128, 21.36681, 21.60553, 21.84418, 22.08273, 
    22.32119, 22.55955, 22.7978, 23.03594, 23.27397, 23.51188, 23.74965, 
    23.9873, 24.2248, 24.46217, 24.69938, 24.93644, 25.17335, 25.41008, 
    25.64665, 25.88305, 26.11926, 26.35529, 26.59113, 26.82678, 27.06223, 
    27.29747, 27.5325, 27.76732, 28.00191, 28.23629, 28.47043, 28.70434, 
    28.93801, 29.17144, 29.40462, 29.63755, 29.87022, 30.10262, 30.33477, 
    30.56664, 30.79823, 31.02955, 31.26058, 31.49132, 31.72177, 31.95193, 
    32.18178, 32.41132, 32.64056, 32.86949, 33.09809, 33.32638, 33.55434, 
    33.78197, 34.00926, 34.23622, 34.46284, 34.68912, 34.91504, 35.14062, 
    35.36584, 35.59069, 35.81519, 36.03933, 36.26309, 36.48648, 36.7095, 
    36.93213, 37.15438, 37.37625, 37.59773, 37.81882, 38.03951, 38.25981, 
    38.4797, 38.69919, 38.91828, 39.13696, 39.35522, 39.57307, 39.7905, 
    40.00752, 40.22411, 40.44028, 40.65602, 40.87133, 41.08622, 41.30066, 
    41.51467, 41.72824, 41.94138, 42.15406, 42.36631, 42.57811, 42.78946, 
    43.00035, 43.2108, 43.42079, 43.63033, 43.83941, 44.04802, 44.25618, 
    44.46388, 44.67111, 44.87787, 45.08417, 45.29, 45.49536, 45.70025, 
    45.90467, 46.10861, 46.31208, 46.51507, 46.71758, 46.91962, 47.12117, 
    47.32225, 47.52285, 47.72296, 47.92259, 48.12173, 48.32039, 48.51857, 
    48.71626, 48.91346, 49.11017, 49.3064, 49.50214, 49.69739, 49.89215, 
    50.08641, 50.28019, 50.47348, 50.66628, 50.85858, 51.05039, 51.24171, 
    51.43254, 51.62288, 51.81272, 52.00207, 52.19093, 52.37929, 52.56716, 
    52.75454, 52.94143, 53.12782, 53.31372, 53.49912, 53.68404, 53.86846, 
    54.05239, 54.23582, 54.41877, 54.60123, 54.78319, 54.96466, 55.14565,
  -34.04179, -33.90221, -33.76225, -33.62189, -33.48114, -33.33999, 
    -33.19846, -33.05652, -32.91418, -32.77145, -32.62831, -32.48478, 
    -32.34084, -32.19649, -32.05173, -31.90657, -31.761, -31.61502, 
    -31.46862, -31.32182, -31.17459, -31.02695, -30.87889, -30.73041, 
    -30.58151, -30.43218, -30.28244, -30.13226, -29.98166, -29.83064, 
    -29.67918, -29.52729, -29.37498, -29.22222, -29.06903, -28.91541, 
    -28.76135, -28.60685, -28.45191, -28.29653, -28.1407, -27.98443, 
    -27.82772, -27.67056, -27.51295, -27.35489, -27.19639, -27.03743, 
    -26.87802, -26.71815, -26.55783, -26.39705, -26.23582, -26.07412, 
    -25.91197, -25.74935, -25.58628, -25.42273, -25.25873, -25.09426, 
    -24.92932, -24.76391, -24.59804, -24.4317, -24.26488, -24.0976, 
    -23.92984, -23.7616, -23.59289, -23.42371, -23.25405, -23.08391, 
    -22.91329, -22.7422, -22.57062, -22.39856, -22.22602, -22.053, -21.87949, 
    -21.7055, -21.53103, -21.35606, -21.18062, -21.00468, -20.82826, 
    -20.65134, -20.47394, -20.29605, -20.11767, -19.9388, -19.75943, 
    -19.57958, -19.39923, -19.21839, -19.03705, -18.85522, -18.6729, 
    -18.49008, -18.30677, -18.12296, -17.93866, -17.75386, -17.56856, 
    -17.38277, -17.19648, -17.0097, -16.82242, -16.63464, -16.44636, 
    -16.25759, -16.06833, -15.87856, -15.6883, -15.49754, -15.30629, 
    -15.11454, -14.92229, -14.72955, -14.53631, -14.34257, -14.14835, 
    -13.95362, -13.75841, -13.5627, -13.36649, -13.1698, -12.97261, 
    -12.77493, -12.57676, -12.3781, -12.17895, -11.97931, -11.77918, 
    -11.57857, -11.37747, -11.17588, -10.97381, -10.77126, -10.56822, 
    -10.36471, -10.16071, -9.956236, -9.751283, -9.545853, -9.339947, 
    -9.133568, -8.926716, -8.719394, -8.511601, -8.303341, -8.094613, 
    -7.885421, -7.675766, -7.465649, -7.255072, -7.044037, -6.832545, 
    -6.620599, -6.408201, -6.195352, -5.982055, -5.768311, -5.554123, 
    -5.339492, -5.124422, -4.908914, -4.692971, -4.476594, -4.259787, 
    -4.042552, -3.82489, -3.606806, -3.388301, -3.169378, -2.95004, -2.73029, 
    -2.510129, -2.289562, -2.068591, -1.847219, -1.625448, -1.403283, 
    -1.180726, -0.9577795, -0.7344477, -0.5107334, -0.28664, -0.06217084, 
    0.1626708, 0.3878815, 0.6134578, 0.8393961, 1.065693, 1.292345, 1.519347, 
    1.746698, 1.974392, 2.202426, 2.430796, 2.659499, 2.88853, 3.117885, 
    3.34756, 3.577551, 3.807855, 4.038466, 4.269382, 4.500597, 4.732107, 
    4.963908, 5.195995, 5.428364, 5.661012, 5.893932, 6.12712, 6.360573, 
    6.594286, 6.828253, 7.06247, 7.296932, 7.531635, 7.766574, 8.001744, 
    8.23714, 8.472756, 8.70859, 8.944634, 9.180885, 9.417336, 9.653985, 
    9.890824, 10.12785, 10.36505, 10.60244, 10.83999, 11.0777, 11.31558, 
    11.55361, 11.79179, 12.03012, 12.26858, 12.50718, 12.7459, 12.98475, 
    13.22371, 13.46278, 13.70196, 13.94124, 14.18062, 14.42008, 14.65963, 
    14.89926, 15.13896, 15.37873, 15.61856, 15.85844, 16.09838, 16.33836, 
    16.57837, 16.81843, 17.05851, 17.29861, 17.53873, 17.77886, 18.01899, 
    18.25913, 18.49925, 18.73937, 18.97947, 19.21955, 19.45959, 19.69961, 
    19.93958, 20.17951, 20.41938, 20.6592, 20.89896, 21.13865, 21.37826, 
    21.6178, 21.85725, 22.09661, 22.33588, 22.57504, 22.8141, 23.05304, 
    23.29187, 23.53057, 23.76915, 24.00759, 24.24589, 24.48405, 24.72206, 
    24.95991, 25.1976, 25.43513, 25.67248, 25.90966, 26.14665, 26.38346, 
    26.62008, 26.8565, 27.09272, 27.32873, 27.56453, 27.80011, 28.03547, 
    28.27061, 28.50551, 28.74017, 28.9746, 29.20877, 29.4427, 29.67637, 
    29.90978, 30.14293, 30.37581, 30.60841, 30.84074, 31.07278, 31.30453, 
    31.536, 31.76716, 31.99803, 32.2286, 32.45885, 32.68879, 32.91842, 
    33.14772, 33.3767, 33.60535, 33.83367, 34.06165, 34.28929, 34.51658, 
    34.74353, 34.97013, 35.19637, 35.42225, 35.64777, 35.87292, 36.0977, 
    36.32211, 36.54615, 36.7698, 36.99307, 37.21596, 37.43845, 37.66056, 
    37.88226, 38.10357, 38.32448, 38.54498, 38.76508, 38.98476, 39.20404, 
    39.42289, 39.64133, 39.85935, 40.07694, 40.29411, 40.51085, 40.72716, 
    40.94303, 41.15847, 41.37347, 41.58803, 41.80215, 42.01582, 42.22905, 
    42.44183, 42.65416, 42.86603, 43.07745, 43.28841, 43.49892, 43.70896, 
    43.91854, 44.12766, 44.33632, 44.5445, 44.75222, 44.95947, 45.16624, 
    45.37255, 45.57838, 45.78373, 45.98861, 46.19301, 46.39693, 46.60037, 
    46.80333, 47.00581, 47.2078, 47.40931, 47.61033, 47.81087, 48.01092, 
    48.21048, 48.40955, 48.60814, 48.80623, 49.00383, 49.20094, 49.39756, 
    49.59369, 49.78932, 49.98446, 50.1791, 50.37325, 50.56691, 50.76007, 
    50.95273, 51.1449, 51.33657, 51.52775, 51.71843, 51.90861, 52.0983, 
    52.28749, 52.47618, 52.66438, 52.85207, 53.03928, 53.22598, 53.41219, 
    53.5979, 53.78312, 53.96784, 54.15207, 54.3358, 54.51903, 54.70177, 
    54.88402, 55.06577, 55.24702,
  -34.15669, -34.01707, -33.87707, -33.73667, -33.59587, -33.45469, -33.3131, 
    -33.17112, -33.02873, -32.88594, -32.74276, -32.59916, -32.45517, 
    -32.31076, -32.16594, -32.02072, -31.87508, -31.72903, -31.58257, 
    -31.43569, -31.28839, -31.14068, -30.99254, -30.84398, -30.695, -30.5456, 
    -30.39577, -30.24551, -30.09482, -29.9437, -29.79215, -29.64017, 
    -29.48775, -29.3349, -29.18161, -29.02788, -28.87372, -28.71911, 
    -28.56406, -28.40856, -28.25262, -28.09624, -27.93941, -27.78212, 
    -27.62439, -27.46621, -27.30757, -27.14848, -26.98893, -26.82893, 
    -26.66847, -26.50755, -26.34617, -26.18432, -26.02202, -25.85925, 
    -25.69602, -25.53232, -25.36815, -25.20352, -25.03842, -24.87284, 
    -24.70679, -24.54028, -24.37328, -24.20582, -24.03787, -23.86945, 
    -23.70056, -23.53118, -23.36132, -23.19098, -23.02017, -22.84887, 
    -22.67708, -22.50481, -22.33206, -22.15882, -21.98509, -21.81088, 
    -21.63617, -21.46098, -21.2853, -21.10913, -20.93246, -20.75531, 
    -20.57766, -20.39952, -20.22088, -20.04176, -19.86213, -19.68201, 
    -19.50139, -19.32028, -19.13867, -18.95657, -18.77396, -18.59086, 
    -18.40726, -18.22316, -18.03856, -17.85346, -17.66786, -17.48176, 
    -17.29516, -17.10806, -16.92047, -16.73236, -16.54376, -16.35466, 
    -16.16506, -15.97496, -15.78436, -15.59325, -15.40165, -15.20955, 
    -15.01694, -14.82384, -14.63024, -14.43614, -14.24153, -14.04644, 
    -13.85084, -13.65474, -13.45815, -13.26106, -13.06347, -12.86539, 
    -12.66682, -12.46775, -12.26818, -12.06813, -11.86758, -11.66654, 
    -11.46501, -11.26299, -11.06048, -10.85748, -10.654, -10.45004, 
    -10.24558, -10.04065, -9.83523, -9.629332, -9.422954, -9.216098, 
    -9.008765, -8.800957, -8.592675, -8.383921, -8.174695, -7.965001, 
    -7.754839, -7.544211, -7.333119, -7.121564, -6.909549, -6.697075, 
    -6.484145, -6.270759, -6.056921, -5.842632, -5.627895, -5.412711, 
    -5.197083, -4.981013, -4.764503, -4.547556, -4.330174, -4.11236, 
    -3.894116, -3.675445, -3.456348, -3.23683, -3.016893, -2.796538, 
    -2.57577, -2.354591, -2.133004, -1.911012, -1.688618, -1.465825, 
    -1.242635, -1.019053, -0.7950816, -0.5707237, -0.3459826, -0.1208619, 
    0.1046352, 0.3305051, 0.5567443, 0.7833494, 1.010317, 1.237643, 1.465323, 
    1.693355, 1.921735, 2.150458, 2.37952, 2.608918, 2.838649, 3.068707, 
    3.299088, 3.529789, 3.760806, 3.992134, 4.223769, 4.455706, 4.687942, 
    4.920472, 5.153292, 5.386397, 5.619782, 5.853444, 6.087377, 6.321577, 
    6.556039, 6.790759, 7.025732, 7.260952, 7.496417, 7.732119, 7.968055, 
    8.204219, 8.440607, 8.677214, 8.914034, 9.151063, 9.388295, 9.625726, 
    9.86335, 10.10116, 10.33916, 10.57733, 10.81567, 11.05418, 11.29286, 
    11.53169, 11.77067, 12.00979, 12.24906, 12.48846, 12.72799, 12.96764, 
    13.20742, 13.4473, 13.68729, 13.92738, 14.16757, 14.40785, 14.64822, 
    14.88866, 15.12918, 15.36976, 15.61041, 15.85112, 16.09187, 16.33267, 
    16.57351, 16.81438, 17.05528, 17.29621, 17.53715, 17.7781, 18.01906, 
    18.26001, 18.50097, 18.7419, 18.98282, 19.22372, 19.46459, 19.70542, 
    19.94622, 20.18696, 20.42766, 20.6683, 20.90887, 21.14938, 21.38981, 
    21.63016, 21.87043, 22.1106, 22.35068, 22.59065, 22.83052, 23.07027, 
    23.30991, 23.54942, 23.7888, 24.02804, 24.26715, 24.5061, 24.74491, 
    24.98355, 25.22204, 25.46036, 25.6985, 25.93647, 26.17425, 26.41184, 
    26.64924, 26.88644, 27.12344, 27.36023, 27.5968, 27.83315, 28.06928, 
    28.30518, 28.54085, 28.77627, 29.01145, 29.24639, 29.48107, 29.71549, 
    29.94965, 30.18354, 30.41715, 30.6505, 30.88356, 31.11633, 31.34881, 
    31.581, 31.81289, 32.04448, 32.27576, 32.50673, 32.73738, 32.9677, 
    33.19771, 33.42739, 33.65673, 33.88575, 34.11441, 34.34274, 34.57072, 
    34.79834, 35.02561, 35.25252, 35.47907, 35.70525, 35.93106, 36.1565, 
    36.38156, 36.60624, 36.83054, 37.05445, 37.27797, 37.50109, 37.72382, 
    37.94616, 38.16808, 38.38961, 38.61072, 38.83142, 39.05171, 39.27158, 
    39.49104, 39.71006, 39.92867, 40.14684, 40.36459, 40.5819, 40.79878, 
    41.01522, 41.23122, 41.44678, 41.66189, 41.87656, 42.09078, 42.30454, 
    42.51786, 42.73072, 42.94312, 43.15506, 43.36654, 43.57756, 43.78811, 
    43.9982, 44.20782, 44.41697, 44.62565, 44.83386, 45.04159, 45.24885, 
    45.45563, 45.66193, 45.86776, 46.0731, 46.27795, 46.48233, 46.68622, 
    46.88963, 47.09255, 47.29498, 47.49692, 47.69837, 47.89933, 48.09981, 
    48.29979, 48.49927, 48.69826, 48.89676, 49.09476, 49.29227, 49.48928, 
    49.68579, 49.88181, 50.07733, 50.27235, 50.46687, 50.6609, 50.85442, 
    51.04744, 51.23997, 51.43199, 51.62352, 51.81454, 52.00507, 52.19509, 
    52.38461, 52.57363, 52.76215, 52.95017, 53.13769, 53.32471, 53.51123, 
    53.69725, 53.88277, 54.06779, 54.25231, 54.43633, 54.61985, 54.80288, 
    54.9854, 55.16743, 55.34896,
  -34.27205, -34.1324, -33.99235, -33.85191, -33.71107, -33.56984, -33.42821, 
    -33.28618, -33.14375, -33.00091, -32.85767, -32.71402, -32.56997, 
    -32.42551, -32.28063, -32.13535, -31.98965, -31.84353, -31.697, 
    -31.55005, -31.40269, -31.2549, -31.10669, -30.95805, -30.80899, 
    -30.65951, -30.50959, -30.35925, -30.20847, -30.05727, -29.90563, 
    -29.75355, -29.60104, -29.44809, -29.2947, -29.14087, -28.9866, 
    -28.83188, -28.67672, -28.52112, -28.36506, -28.20856, -28.05161, 
    -27.89421, -27.73635, -27.57804, -27.41928, -27.26005, -27.10037, 
    -26.94024, -26.77964, -26.61857, -26.45705, -26.29506, -26.13261, 
    -25.96969, -25.8063, -25.64245, -25.47812, -25.31332, -25.14805, 
    -24.98231, -24.81609, -24.6494, -24.48223, -24.31458, -24.14646, 
    -23.97785, -23.80877, -23.6392, -23.46915, -23.29861, -23.12759, 
    -22.95609, -22.7841, -22.61162, -22.43865, -22.2652, -22.09125, 
    -21.91681, -21.74188, -21.56646, -21.39055, -21.21414, -21.03724, 
    -20.85984, -20.68194, -20.50355, -20.32467, -20.14528, -19.96539, 
    -19.78501, -19.60413, -19.42275, -19.24086, -19.05848, -18.87559, 
    -18.69221, -18.50832, -18.32392, -18.13903, -17.95363, -17.76773, 
    -17.58132, -17.39441, -17.207, -17.01908, -16.83066, -16.64174, -16.4523, 
    -16.26237, -16.07193, -15.88099, -15.68954, -15.49758, -15.30513, 
    -15.11217, -14.9187, -14.72473, -14.53026, -14.33529, -14.13981, 
    -13.94383, -13.74735, -13.55037, -13.35289, -13.1549, -12.95642, 
    -12.75744, -12.55796, -12.35798, -12.1575, -11.95653, -11.75506, 
    -11.5531, -11.35065, -11.1477, -10.94426, -10.74033, -10.53591, -10.331, 
    -10.1256, -9.91972, -9.713351, -9.506499, -9.299165, -9.09135, -8.883055, 
    -8.674281, -8.465032, -8.255306, -8.045107, -7.834436, -7.623296, 
    -7.411686, -7.19961, -6.987069, -6.774065, -6.5606, -6.346675, -6.132294, 
    -5.917458, -5.702168, -5.486428, -5.27024, -5.053606, -4.836527, 
    -4.619007, -4.401048, -4.182652, -3.963822, -3.74456, -3.52487, 
    -3.304753, -3.084213, -2.863251, -2.641872, -2.420078, -2.197872, 
    -1.975257, -1.752235, -1.52881, -1.304985, -1.080764, -0.8561485, 
    -0.631143, -0.4057505, -0.1799744, 0.04618191, 0.272715, 0.4996212, 
    0.7268971, 0.9545391, 1.182543, 1.410906, 1.639624, 1.868693, 2.098109, 
    2.327868, 2.557967, 2.788401, 3.019166, 3.250259, 3.481674, 3.713408, 
    3.945457, 4.177817, 4.410482, 4.643449, 4.876713, 5.11027, 5.344115, 
    5.578244, 5.812652, 6.047335, 6.282288, 6.517505, 6.752983, 6.988717, 
    7.224701, 7.460932, 7.697403, 7.934111, 8.171049, 8.408214, 8.645599, 
    8.883202, 9.121015, 9.359033, 9.597252, 9.835667, 10.07427, 10.31306, 
    10.55203, 10.79117, 11.03048, 11.26996, 11.50959, 11.74938, 11.98931, 
    12.22939, 12.4696, 12.70994, 12.95041, 13.191, 13.4317, 13.67251, 
    13.91342, 14.15443, 14.39553, 14.63671, 14.87798, 15.11932, 15.36073, 
    15.6022, 15.84373, 16.08531, 16.32694, 16.56861, 16.81031, 17.05204, 
    17.29379, 17.53556, 17.77734, 18.01912, 18.26091, 18.50269, 18.74445, 
    18.9862, 19.22793, 19.46962, 19.71128, 19.9529, 20.19448, 20.436, 
    20.67746, 20.91886, 21.16019, 21.40144, 21.64262, 21.8837, 22.1247, 
    22.36559, 22.60639, 22.84707, 23.08764, 23.32808, 23.56841, 23.8086, 
    24.04865, 24.28856, 24.52832, 24.76793, 25.00738, 25.24667, 25.48578, 
    25.72472, 25.96348, 26.20206, 26.44044, 26.67863, 26.91662, 27.1544, 
    27.39197, 27.62932, 27.86645, 28.10335, 28.34002, 28.57645, 28.81264, 
    29.04859, 29.28428, 29.51972, 29.7549, 29.98981, 30.22445, 30.45881, 
    30.69289, 30.92669, 31.16021, 31.39342, 31.62634, 31.85896, 32.09127, 
    32.32327, 32.55495, 32.78632, 33.01736, 33.24807, 33.47845, 33.7085, 
    33.9382, 34.16756, 34.39658, 34.62524, 34.85355, 35.08149, 35.30908, 
    35.5363, 35.76315, 35.98962, 36.21571, 36.44143, 36.66676, 36.8917, 
    37.11626, 37.34042, 37.56418, 37.78754, 38.0105, 38.23305, 38.45519, 
    38.67692, 38.89823, 39.11913, 39.3396, 39.55965, 39.77927, 39.99847, 
    40.21723, 40.43555, 40.65344, 40.8709, 41.0879, 41.30447, 41.52058, 
    41.73625, 41.95147, 42.16624, 42.38055, 42.5944, 42.80779, 43.02072, 
    43.23319, 43.44519, 43.65673, 43.86779, 44.07839, 44.28851, 44.49816, 
    44.70734, 44.91603, 45.12426, 45.33199, 45.53925, 45.74603, 45.95232, 
    46.15813, 46.36345, 46.56828, 46.77262, 46.97647, 47.17984, 47.38271, 
    47.58508, 47.78697, 47.98835, 48.18925, 48.38964, 48.58955, 48.78895, 
    48.98785, 49.18625, 49.38416, 49.58156, 49.77847, 49.97486, 50.17076, 
    50.36616, 50.56106, 50.75545, 50.94934, 51.14272, 51.33561, 51.52798, 
    51.71985, 51.91122, 52.10209, 52.29245, 52.4823, 52.67165, 52.8605, 
    53.04884, 53.23668, 53.42401, 53.61084, 53.79717, 53.98299, 54.16831, 
    54.35312, 54.53744, 54.72125, 54.90456, 55.08736, 55.26967, 55.45147,
  -34.38787, -34.24818, -34.1081, -33.96762, -33.82675, -33.68547, -33.5438, 
    -33.40172, -33.25924, -33.11636, -32.97306, -32.82936, -32.68526, 
    -32.54074, -32.39581, -32.25046, -32.1047, -31.95852, -31.81193, 
    -31.66491, -31.51747, -31.36961, -31.22133, -31.07262, -30.92348, 
    -30.77392, -30.62392, -30.4735, -30.32264, -30.17134, -30.01961, 
    -29.86744, -29.71484, -29.56179, -29.4083, -29.25437, -29.1, -28.94518, 
    -28.78991, -28.63419, -28.47803, -28.32141, -28.16434, -28.00682, 
    -27.84884, -27.69041, -27.53151, -27.37216, -27.21235, -27.05208, 
    -26.89134, -26.73014, -26.56847, -26.40634, -26.24374, -26.08067, 
    -25.91713, -25.75312, -25.58863, -25.42367, -25.25824, -25.09233, 
    -24.92594, -24.75908, -24.59173, -24.42391, -24.2556, -24.08681, 
    -23.91753, -23.74778, -23.57753, -23.4068, -23.23558, -23.06387, 
    -22.89167, -22.71899, -22.54581, -22.37214, -22.19797, -22.02331, 
    -21.84816, -21.67251, -21.49636, -21.31972, -21.14257, -20.96494, 
    -20.78679, -20.60816, -20.42902, -20.24937, -20.06923, -19.88858, 
    -19.70744, -19.52578, -19.34362, -19.16096, -18.9778, -18.79412, 
    -18.60995, -18.42526, -18.24007, -18.05437, -17.86817, -17.68146, 
    -17.49424, -17.30651, -17.11827, -16.92953, -16.74028, -16.55052, 
    -16.36025, -16.16947, -15.97819, -15.78639, -15.59409, -15.40128, 
    -15.20796, -15.01413, -14.8198, -14.62496, -14.42961, -14.23376, 
    -14.0374, -13.84053, -13.64316, -13.44528, -13.2469, -13.04801, 
    -12.84862, -12.64873, -12.44834, -12.24744, -12.04605, -11.84415, 
    -11.64176, -11.43886, -11.23547, -11.03159, -10.82721, -10.62233, 
    -10.41697, -10.21111, -10.00476, -9.797917, -9.59059, -9.382775, 
    -9.174476, -8.965692, -8.756426, -8.546678, -8.336451, -8.125746, 
    -7.914565, -7.702909, -7.490779, -7.27818, -7.065111, -6.851574, 
    -6.637572, -6.423106, -6.208179, -5.992793, -5.776949, -5.560651, 
    -5.343899, -5.126698, -4.909047, -4.690951, -4.472412, -4.253431, 
    -4.034012, -3.814158, -3.59387, -3.373152, -3.152005, -2.930434, 
    -2.708441, -2.486028, -2.263199, -2.039957, -1.816304, -1.592245, 
    -1.367781, -1.142916, -0.9176533, -0.6919966, -0.4659488, -0.2395134, 
    -0.0126938, 0.2145064, 0.4420837, 0.6700346, 0.8983553, 1.127042, 
    1.356091, 1.5855, 1.815262, 2.045376, 2.275836, 2.50664, 2.737782, 
    2.96926, 3.201068, 3.433202, 3.665659, 3.898434, 4.131523, 4.364921, 
    4.598623, 4.832626, 5.066926, 5.301517, 5.536394, 5.771554, 6.006991, 
    6.242702, 6.47868, 6.714921, 6.951421, 7.188175, 7.425177, 7.662423, 
    7.899908, 8.137627, 8.375573, 8.613744, 8.852134, 9.090735, 9.329546, 
    9.56856, 9.807771, 10.04717, 10.28676, 10.52654, 10.76648, 11.0066, 
    11.24689, 11.48733, 11.72793, 11.96868, 12.20957, 12.45059, 12.69175, 
    12.93304, 13.17445, 13.41597, 13.65761, 13.89934, 14.14118, 14.38311, 
    14.62512, 14.86721, 15.10939, 15.35163, 15.59393, 15.83629, 16.0787, 
    16.32116, 16.56367, 16.8062, 17.04876, 17.29135, 17.53395, 17.77657, 
    18.01919, 18.26181, 18.50442, 18.74702, 18.98961, 19.23217, 19.4747, 
    19.71719, 19.95964, 20.20205, 20.4444, 20.6867, 20.92893, 21.17109, 
    21.41317, 21.65517, 21.89708, 22.1389, 22.38062, 22.62224, 22.86374, 
    23.10513, 23.3464, 23.58754, 23.82855, 24.06942, 24.31014, 24.55071, 
    24.79113, 25.03139, 25.27148, 25.5114, 25.75115, 25.99071, 26.23008, 
    26.46926, 26.70824, 26.94702, 27.18559, 27.42394, 27.66208, 27.89999, 
    28.13767, 28.37512, 28.61233, 28.84929, 29.08601, 29.32247, 29.55867, 
    29.7946, 30.03027, 30.26566, 30.50078, 30.73561, 30.97016, 31.20441, 
    31.43836, 31.67202, 31.90537, 32.13841, 32.37113, 32.60354, 32.83562, 
    33.06738, 33.2988, 33.52989, 33.76064, 33.99105, 34.22111, 34.45081, 
    34.68016, 34.90916, 35.13779, 35.36605, 35.59394, 35.82146, 36.0486, 
    36.27536, 36.50173, 36.72772, 36.95331, 37.17851, 37.40331, 37.62771, 
    37.85171, 38.0753, 38.29847, 38.52124, 38.74358, 38.96551, 39.18702, 
    39.40809, 39.62875, 39.84896, 40.06875, 40.2881, 40.50701, 40.72548, 
    40.9435, 41.16108, 41.37822, 41.59489, 41.81112, 42.02689, 42.24221, 
    42.45706, 42.67146, 42.88538, 43.09885, 43.31184, 43.52436, 43.73642, 
    43.948, 44.15911, 44.36974, 44.57989, 44.78956, 44.99875, 45.20746, 
    45.41568, 45.62342, 45.83067, 46.03743, 46.2437, 46.44949, 46.65477, 
    46.85957, 47.06387, 47.26768, 47.47099, 47.67381, 47.87612, 48.07794, 
    48.27925, 48.48007, 48.68038, 48.8802, 49.07951, 49.27831, 49.47661, 
    49.67441, 49.8717, 50.06849, 50.26477, 50.46054, 50.65582, 50.85057, 
    51.04483, 51.23857, 51.43181, 51.62454, 51.81676, 52.00848, 52.19968, 
    52.39038, 52.58057, 52.77025, 52.95942, 53.14808, 53.33624, 53.52389, 
    53.71103, 53.89766, 54.08378, 54.2694, 54.45451, 54.63911, 54.82321, 
    55.00681, 55.18989, 55.37247, 55.55455,
  -34.50416, -34.36444, -34.22432, -34.08381, -33.94289, -33.80157, 
    -33.65986, -33.51774, -33.37521, -33.23228, -33.08894, -32.94519, 
    -32.80103, -32.65646, -32.51147, -32.36606, -32.22024, -32.074, 
    -31.92734, -31.78026, -31.63276, -31.48483, -31.33647, -31.18769, 
    -31.03848, -30.88883, -30.73876, -30.58825, -30.4373, -30.28592, 
    -30.13411, -29.98185, -29.82915, -29.67601, -29.52242, -29.36839, 
    -29.21392, -29.05899, -28.90362, -28.74779, -28.59152, -28.43479, 
    -28.2776, -28.11996, -27.96186, -27.8033, -27.64429, -27.48481, 
    -27.32486, -27.16446, -27.00358, -26.84224, -26.68044, -26.51816, 
    -26.35541, -26.19219, -26.0285, -25.86433, -25.69969, -25.53457, 
    -25.36897, -25.2029, -25.03634, -24.86931, -24.70179, -24.53378, 
    -24.3653, -24.19632, -24.02686, -23.85691, -23.68647, -23.51555, 
    -23.34413, -23.17222, -22.99982, -22.82692, -22.65353, -22.47964, 
    -22.30526, -22.13038, -21.955, -21.77912, -21.60275, -21.42587, 
    -21.24849, -21.0706, -20.89222, -20.71333, -20.53394, -20.35404, 
    -20.17364, -19.99273, -19.81132, -19.62939, -19.44696, -19.26403, 
    -19.08058, -18.89662, -18.71216, -18.52718, -18.3417, -18.1557, 
    -17.96919, -17.78217, -17.59464, -17.4066, -17.21805, -17.02898, 
    -16.8394, -16.64931, -16.45871, -16.26759, -16.07597, -15.88383, 
    -15.69117, -15.49801, -15.30433, -15.11015, -14.91545, -14.72023, 
    -14.52451, -14.32828, -14.13153, -13.93428, -13.73652, -13.53824, 
    -13.33946, -13.14017, -12.94038, -12.74007, -12.53926, -12.33795, 
    -12.13613, -11.9338, -11.73097, -11.52764, -11.32381, -11.11948, 
    -10.91465, -10.70932, -10.50349, -10.29717, -10.09035, -9.883036, 
    -9.675231, -9.466935, -9.258149, -9.048875, -8.839113, -8.628866, 
    -8.418136, -8.206923, -7.995228, -7.783055, -7.570405, -7.357279, 
    -7.143679, -6.929608, -6.715066, -6.500058, -6.284583, -6.068644, 
    -5.852243, -5.635384, -5.418067, -5.200294, -4.982069, -4.763395, 
    -4.544272, -4.324704, -4.104693, -3.884243, -3.663354, -3.442031, 
    -3.220276, -2.998091, -2.775481, -2.552446, -2.328991, -2.105119, 
    -1.880831, -1.656133, -1.431026, -1.205515, -0.9796011, -0.7532892, 
    -0.5265822, -0.2994836, -0.07199687, 0.1558746, 0.384127, 0.612757, 
    0.8417607, 1.071134, 1.300874, 1.530977, 1.761438, 1.992254, 2.22342, 
    2.454933, 2.686789, 2.918983, 3.151511, 3.384369, 3.617553, 3.851059, 
    4.084882, 4.319017, 4.553461, 4.788208, 5.023255, 5.258596, 5.494228, 
    5.730145, 5.966342, 6.202815, 6.439559, 6.67657, 6.913842, 7.15137, 
    7.38915, 7.627176, 7.865444, 8.103948, 8.342683, 8.581644, 8.820827, 
    9.060225, 9.299832, 9.539646, 9.779659, 10.01987, 10.26026, 10.50084, 
    10.7416, 10.98253, 11.22363, 11.46489, 11.70631, 11.94788, 12.18959, 
    12.43144, 12.67343, 12.91554, 13.15777, 13.40013, 13.64259, 13.88516, 
    14.12782, 14.37059, 14.61343, 14.85637, 15.09937, 15.34245, 15.58559, 
    15.82879, 16.07204, 16.31534, 16.55868, 16.80206, 17.04546, 17.28889, 
    17.53234, 17.77579, 18.01926, 18.26272, 18.50617, 18.74961, 18.99304, 
    19.23644, 19.47981, 19.72314, 19.96644, 20.20968, 20.45287, 20.69601, 
    20.93907, 21.18207, 21.42499, 21.66782, 21.91057, 22.15322, 22.39577, 
    22.63822, 22.88055, 23.12277, 23.36486, 23.60682, 23.84866, 24.09035, 
    24.33189, 24.57328, 24.81452, 25.05559, 25.29649, 25.53722, 25.77777, 
    26.01814, 26.25832, 26.4983, 26.73808, 26.97766, 27.21702, 27.45617, 
    27.6951, 27.9338, 28.17226, 28.41049, 28.64848, 28.88622, 29.12371, 
    29.36094, 29.59791, 29.83461, 30.07104, 30.30719, 30.54306, 30.77865, 
    31.01394, 31.24895, 31.48364, 31.71804, 31.95213, 32.1859, 32.41935, 
    32.65249, 32.88529, 33.11777, 33.34991, 33.58171, 33.81317, 34.04428, 
    34.27504, 34.50544, 34.73549, 34.96517, 35.19449, 35.42344, 35.652, 
    35.8802, 36.10801, 36.33543, 36.56247, 36.78912, 37.01536, 37.24121, 
    37.46666, 37.6917, 37.91634, 38.14056, 38.36436, 38.58775, 38.81072, 
    39.03326, 39.25538, 39.47707, 39.69833, 39.91914, 40.13953, 40.35947, 
    40.57896, 40.79802, 41.01662, 41.23477, 41.45247, 41.66972, 41.88651, 
    42.10283, 42.3187, 42.5341, 42.74903, 42.9635, 43.1775, 43.39102, 
    43.60407, 43.81665, 44.02875, 44.24036, 44.4515, 44.66216, 44.87233, 
    45.08201, 45.29121, 45.49992, 45.70813, 45.91586, 46.1231, 46.32984, 
    46.53608, 46.74183, 46.94708, 47.15183, 47.35609, 47.55984, 47.76309, 
    47.96584, 48.16808, 48.36982, 48.57106, 48.77179, 48.97202, 49.17173, 
    49.37094, 49.56964, 49.76783, 49.96552, 50.16269, 50.35935, 50.5555, 
    50.75115, 50.94628, 51.1409, 51.335, 51.5286, 51.72168, 51.91425, 
    52.10631, 52.29786, 52.4889, 52.67942, 52.86942, 53.05892, 53.24791, 
    53.43638, 53.62434, 53.81179, 53.99873, 54.18515, 54.37107, 54.55648, 
    54.74137, 54.92575, 55.10963, 55.293, 55.47586, 55.65821,
  -34.62092, -34.48116, -34.34101, -34.20046, -34.05951, -33.91816, -33.7764, 
    -33.63424, -33.49166, -33.34869, -33.2053, -33.0615, -32.91729, 
    -32.77266, -32.62762, -32.48216, -32.33628, -32.18998, -32.04325, 
    -31.89611, -31.74854, -31.60054, -31.45212, -31.30326, -31.15397, 
    -31.00426, -30.8541, -30.70351, -30.55248, -30.40102, -30.24911, 
    -30.09677, -29.94398, -29.79074, -29.63706, -29.48293, -29.32836, 
    -29.17333, -29.01785, -28.86192, -28.70554, -28.54869, -28.39139, 
    -28.23363, -28.07542, -27.91674, -27.7576, -27.59799, -27.43792, 
    -27.27738, -27.11637, -26.95489, -26.79295, -26.63053, -26.46763, 
    -26.30427, -26.14042, -25.9761, -25.8113, -25.64602, -25.48027, 
    -25.31403, -25.1473, -24.98009, -24.8124, -24.64422, -24.47555, -24.3064, 
    -24.13675, -23.96661, -23.79598, -23.62486, -23.45325, -23.28114, 
    -23.10853, -22.93542, -22.76182, -22.58772, -22.41312, -22.23802, 
    -22.06242, -21.88631, -21.7097, -21.53259, -21.35497, -21.17685, 
    -20.99822, -20.81909, -20.63944, -20.45929, -20.27863, -20.09746, 
    -19.91578, -19.73359, -19.55089, -19.36767, -19.18394, -18.9997, 
    -18.81495, -18.62968, -18.4439, -18.25761, -18.0708, -17.88347, 
    -17.69563, -17.50728, -17.3184, -17.12901, -16.93911, -16.74869, 
    -16.55775, -16.3663, -16.17433, -15.98184, -15.78884, -15.59532, 
    -15.40129, -15.20674, -15.01167, -14.81609, -14.61999, -14.42338, 
    -14.22625, -14.02861, -13.83046, -13.63179, -13.43261, -13.23291, 
    -13.03271, -12.83199, -12.63076, -12.42902, -12.22678, -12.02402, 
    -11.82076, -11.61699, -11.41272, -11.20794, -11.00265, -10.79687, 
    -10.59058, -10.38379, -10.1765, -9.968712, -9.760428, -9.551649, 
    -9.342375, -9.132608, -8.92235, -8.711602, -8.500365, -8.288642, 
    -8.076433, -7.863741, -7.650567, -7.436913, -7.222781, -7.008173, 
    -6.79309, -6.577535, -6.361509, -6.145015, -5.928056, -5.710632, 
    -5.492746, -5.274402, -5.0556, -4.836343, -4.616635, -4.396476, 
    -4.175871, -3.954821, -3.733329, -3.511398, -3.28903, -3.066229, 
    -2.842997, -2.619337, -2.395253, -2.170747, -1.945821, -1.720481, 
    -1.494727, -1.268565, -1.041997, -0.815026, -0.587656, -0.3598903, 
    -0.1317323, 0.09681441, 0.3257462, 0.5550594, 0.7847503, 1.014815, 
    1.24525, 1.476052, 1.707215, 1.938738, 2.170614, 2.402841, 2.635415, 
    2.86833, 3.101583, 3.335171, 3.569087, 3.803328, 4.03789, 4.272768, 
    4.507958, 4.743454, 4.979254, 5.215351, 5.451742, 5.688421, 5.925384, 
    6.162625, 6.400141, 6.637926, 6.875975, 7.114284, 7.352847, 7.591659, 
    7.830715, 8.07001, 8.309539, 8.549297, 8.789278, 9.029477, 9.26989, 
    9.510509, 9.75133, 9.992349, 10.23356, 10.47495, 10.71653, 10.95828, 
    11.2002, 11.44228, 11.68452, 11.92692, 12.16946, 12.41214, 12.65495, 
    12.8979, 13.14097, 13.38416, 13.62745, 13.87086, 14.11437, 14.35797, 
    14.60166, 14.84543, 15.08928, 15.3332, 15.57719, 15.82123, 16.06533, 
    16.30948, 16.55367, 16.79789, 17.04214, 17.28642, 17.53071, 17.77501, 
    18.01932, 18.26363, 18.50794, 18.75223, 18.9965, 19.24075, 19.48496, 
    19.72915, 19.97328, 20.21737, 20.46141, 20.70539, 20.9493, 21.19313, 
    21.4369, 21.68057, 21.92416, 22.16765, 22.41104, 22.65432, 22.89749, 
    23.14054, 23.38346, 23.62626, 23.86892, 24.11144, 24.35381, 24.59602, 
    24.83808, 25.07997, 25.3217, 25.56324, 25.80461, 26.04579, 26.28678, 
    26.52757, 26.76815, 27.00853, 27.2487, 27.48864, 27.72836, 27.96786, 
    28.20712, 28.44613, 28.68491, 28.92343, 29.1617, 29.39971, 29.63745, 
    29.87492, 30.11212, 30.34904, 30.58567, 30.82202, 31.05807, 31.29382, 
    31.52927, 31.76441, 31.99924, 32.23375, 32.46794, 32.7018, 32.93534, 
    33.16854, 33.4014, 33.63391, 33.86609, 34.09791, 34.32938, 34.56048, 
    34.79123, 35.0216, 35.25161, 35.48124, 35.71049, 35.93937, 36.16785, 
    36.39595, 36.62365, 36.85096, 37.07786, 37.30437, 37.53046, 37.75615, 
    37.98143, 38.20629, 38.43073, 38.65474, 38.87834, 39.1015, 39.32423, 
    39.54653, 39.76839, 39.98982, 40.2108, 40.43133, 40.65142, 40.87106, 
    41.09024, 41.30897, 41.52724, 41.74506, 41.96241, 42.17929, 42.39571, 
    42.61166, 42.82714, 43.04215, 43.25668, 43.47074, 43.68432, 43.89742, 
    44.11003, 44.32217, 44.53381, 44.74497, 44.95564, 45.16582, 45.37551, 
    45.58471, 45.79341, 46.00161, 46.20932, 46.41653, 46.62324, 46.82945, 
    47.03516, 47.24036, 47.44506, 47.64926, 47.85295, 48.05613, 48.2588, 
    48.46097, 48.66263, 48.86377, 49.06441, 49.26453, 49.46415, 49.66325, 
    49.86184, 50.05991, 50.25747, 50.45451, 50.65105, 50.84706, 51.04256, 
    51.23755, 51.43202, 51.62597, 51.81941, 52.01233, 52.20473, 52.39662, 
    52.58799, 52.77885, 52.96918, 53.15901, 53.34832, 53.53711, 53.72538, 
    53.91314, 54.10038, 54.28711, 54.47332, 54.65903, 54.84421, 55.02888, 
    55.21304, 55.39669, 55.57982, 55.76244,
  -34.73815, -34.59836, -34.45818, -34.31759, -34.17661, -34.03521, 
    -33.89342, -33.75121, -33.6086, -33.46558, -33.32215, -33.1783, 
    -33.03404, -32.88936, -32.74426, -32.59875, -32.45281, -32.30645, 
    -32.15967, -32.01246, -31.86483, -31.71676, -31.56827, -31.41934, 
    -31.26998, -31.12019, -30.96996, -30.81929, -30.66818, -30.51663, 
    -30.36464, -30.21221, -30.05933, -29.906, -29.75223, -29.598, -29.44333, 
    -29.2882, -29.13262, -28.97658, -28.82009, -28.66313, -28.50572, 
    -28.34785, -28.18951, -28.03071, -27.87144, -27.71171, -27.55151, 
    -27.39084, -27.2297, -27.06809, -26.906, -26.74344, -26.58041, -26.41689, 
    -26.2529, -26.08843, -25.92347, -25.75804, -25.59212, -25.42571, 
    -25.25882, -25.09144, -24.92358, -24.75522, -24.58638, -24.41704, 
    -24.24721, -24.07688, -23.90606, -23.73475, -23.56293, -23.39062, 
    -23.21781, -23.0445, -22.87069, -22.69638, -22.52156, -22.34624, 
    -22.17041, -21.99408, -21.81725, -21.6399, -21.46205, -21.28368, 
    -21.10481, -20.92543, -20.74553, -20.56513, -20.38421, -20.20278, 
    -20.02083, -19.83837, -19.6554, -19.47191, -19.2879, -19.10338, 
    -18.91833, -18.73278, -18.5467, -18.36011, -18.17299, -17.98536, 
    -17.79721, -17.60854, -17.41935, -17.22964, -17.03941, -16.84866, 
    -16.65739, -16.4656, -16.27328, -16.08045, -15.8871, -15.69323, 
    -15.49883, -15.30392, -15.10849, -14.91253, -14.71606, -14.51907, 
    -14.32156, -14.12353, -13.92498, -13.72592, -13.52633, -13.32623, 
    -13.12562, -12.92449, -12.72284, -12.52068, -12.31801, -12.11482, 
    -11.91112, -11.70691, -11.50219, -11.29696, -11.09123, -10.88498, 
    -10.67823, -10.47097, -10.26322, -10.05495, -9.846188, -9.636923, 
    -9.42716, -9.216899, -9.006143, -8.794891, -8.583147, -8.370912, 
    -8.158186, -7.944973, -7.731273, -7.517088, -7.302422, -7.087274, 
    -6.871647, -6.655543, -6.438965, -6.221914, -6.004392, -5.786402, 
    -5.567945, -5.349025, -5.129643, -4.909802, -4.689505, -4.468753, 
    -4.24755, -4.025897, -3.803798, -3.581256, -3.358273, -3.134852, 
    -2.910996, -2.686707, -2.46199, -2.236846, -2.01128, -1.785293, -1.55889, 
    -1.332073, -1.104846, -0.8772123, -0.6491752, -0.4207383, -0.1919051, 
    0.03732099, 0.2669362, 0.4969369, 0.7273193, 0.9580797, 1.189214, 
    1.420719, 1.65259, 1.884823, 2.117415, 2.350361, 2.583657, 2.817298, 
    3.051281, 3.285602, 3.520255, 3.755237, 3.990543, 4.226169, 4.46211, 
    4.698361, 4.934918, 5.171777, 5.408932, 5.646379, 5.884112, 6.122128, 
    6.36042, 6.598985, 6.837818, 7.076912, 7.316264, 7.555867, 7.795718, 
    8.03581, 8.276139, 8.516699, 8.757485, 8.998491, 9.239714, 9.481145, 
    9.722781, 9.964616, 10.20665, 10.44886, 10.69126, 10.93384, 11.17658, 
    11.41949, 11.66257, 11.90579, 12.14917, 12.39268, 12.63634, 12.88012, 
    13.12403, 13.36806, 13.6122, 13.85645, 14.1008, 14.34525, 14.58979, 
    14.83441, 15.07911, 15.32388, 15.56872, 15.81361, 16.05857, 16.30356, 
    16.5486, 16.79368, 17.03879, 17.28392, 17.52907, 17.77423, 18.01939, 
    18.26455, 18.50971, 18.75486, 18.99998, 19.24509, 19.49016, 19.73519, 
    19.98018, 20.22513, 20.47001, 20.71484, 20.9596, 21.20429, 21.4489, 
    21.69342, 21.93785, 22.18219, 22.42642, 22.67055, 22.91456, 23.15845, 
    23.40221, 23.64585, 23.88934, 24.13269, 24.37589, 24.61894, 24.86183, 
    25.10455, 25.3471, 25.58947, 25.83165, 26.07365, 26.31545, 26.55706, 
    26.79846, 27.03965, 27.28062, 27.52137, 27.76189, 28.00218, 28.24224, 
    28.48205, 28.72161, 28.96093, 29.19998, 29.43877, 29.67729, 29.91554, 
    30.15351, 30.3912, 30.6286, 30.86571, 31.10252, 31.33903, 31.57523, 
    31.81112, 32.0467, 32.28196, 32.51688, 32.75149, 32.98575, 33.21968, 
    33.45327, 33.68651, 33.9194, 34.15194, 34.38411, 34.61592, 34.84737, 
    35.07845, 35.30915, 35.53947, 35.76941, 35.99897, 36.22813, 36.4569, 
    36.68527, 36.91325, 37.14082, 37.36798, 37.59473, 37.82107, 38.04699, 
    38.27249, 38.49757, 38.72221, 38.94643, 39.17022, 39.39357, 39.61649, 
    39.83896, 40.06099, 40.28257, 40.5037, 40.72438, 40.94461, 41.16438, 
    41.38369, 41.60253, 41.82092, 42.03883, 42.25628, 42.47326, 42.68976, 
    42.90579, 43.12134, 43.33641, 43.551, 43.76511, 43.97873, 44.19187, 
    44.40451, 44.61667, 44.82834, 45.03951, 45.25019, 45.46037, 45.67006, 
    45.87925, 46.08793, 46.29611, 46.50379, 46.71097, 46.91764, 47.12381, 
    47.32946, 47.53461, 47.73925, 47.94338, 48.147, 48.3501, 48.55269, 
    48.75477, 48.95634, 49.15739, 49.35792, 49.55794, 49.75744, 49.95642, 
    50.15489, 50.35284, 50.55026, 50.74717, 50.94357, 51.13943, 51.33479, 
    51.52962, 51.72393, 51.91772, 52.11099, 52.30374, 52.49597, 52.68768, 
    52.87887, 53.06953, 53.25969, 53.44931, 53.63842, 53.82701, 54.01508, 
    54.20263, 54.38966, 54.57617, 54.76217, 54.94764, 55.1326, 55.31704, 
    55.50097, 55.68438, 55.86727,
  -34.85585, -34.71603, -34.57582, -34.4352, -34.29418, -34.15275, -34.01092, 
    -33.86868, -33.72602, -33.58296, -33.43948, -33.29559, -33.15128, 
    -33.00655, -32.8614, -32.71584, -32.56984, -32.42343, -32.27658, 
    -32.12932, -31.98162, -31.83349, -31.68493, -31.53593, -31.3865, 
    -31.23664, -31.08633, -30.93558, -30.7844, -30.63277, -30.48069, 
    -30.32817, -30.1752, -30.02179, -29.86792, -29.7136, -29.55883, -29.4036, 
    -29.24792, -29.09177, -28.93517, -28.77811, -28.62059, -28.4626, 
    -28.30415, -28.14523, -27.98584, -27.82598, -27.66566, -27.50486, 
    -27.34358, -27.18184, -27.01962, -26.85691, -26.69373, -26.53008, 
    -26.36593, -26.20131, -26.0362, -25.87061, -25.70453, -25.53796, 
    -25.37091, -25.20336, -25.03532, -24.86679, -24.69777, -24.52825, 
    -24.35824, -24.18773, -24.01672, -23.84521, -23.6732, -23.50069, 
    -23.32768, -23.15416, -22.98014, -22.80561, -22.63058, -22.45504, 
    -22.27899, -22.10244, -21.92537, -21.74779, -21.5697, -21.3911, 
    -21.21199, -21.03236, -20.85221, -20.67155, -20.49038, -20.30869, 
    -20.12647, -19.94375, -19.7605, -19.57673, -19.39245, -19.20764, 
    -19.02231, -18.83646, -18.65009, -18.4632, -18.27579, -18.08785, 
    -17.89939, -17.7104, -17.52089, -17.33086, -17.1403, -16.94922, 
    -16.75762, -16.56549, -16.37284, -16.17966, -15.98595, -15.79172, 
    -15.59697, -15.4017, -15.20589, -15.00957, -14.81272, -14.61535, 
    -14.41745, -14.21904, -14.0201, -13.82063, -13.62065, -13.42014, 
    -13.21912, -13.01757, -12.81551, -12.61292, -12.40982, -12.2062, 
    -12.00207, -11.79742, -11.59225, -11.38657, -11.18038, -10.97367, 
    -10.76646, -10.55873, -10.3505, -10.14176, -9.932514, -9.722763, 
    -9.512508, -9.301752, -9.090495, -8.878739, -8.666485, -8.453735, 
    -8.240492, -8.026754, -7.812527, -7.59781, -7.382607, -7.166917, 
    -6.950744, -6.734089, -6.516956, -6.299345, -6.081258, -5.862699, 
    -5.643669, -5.42417, -5.204206, -4.983778, -4.762888, -4.54154, 
    -4.319736, -4.097478, -3.874769, -3.651613, -3.428011, -3.203966, 
    -2.979482, -2.754562, -2.529208, -2.303423, -2.077211, -1.850575, 
    -1.623518, -1.396043, -1.168154, -0.9398531, -0.7111451, -0.482033, 
    -0.2525204, -0.02261083, 0.207692, 0.4383845, 0.6694627, 0.900923, 
    1.132761, 1.364974, 1.597557, 1.830506, 2.063817, 2.297486, 2.531509, 
    2.765882, 3.0006, 3.235659, 3.471054, 3.706782, 3.942837, 4.179216, 
    4.415913, 4.652924, 4.890244, 5.127869, 5.365794, 5.604014, 5.842524, 
    6.081318, 6.320394, 6.559744, 6.799366, 7.039252, 7.279397, 7.519799, 
    7.760449, 8.001345, 8.242479, 8.483848, 8.725445, 8.967264, 9.209302, 
    9.451552, 9.694009, 9.936666, 10.17952, 10.42256, 10.66579, 10.9092, 
    11.15278, 11.39653, 11.64044, 11.8845, 12.12871, 12.37307, 12.61757, 
    12.8622, 13.10696, 13.35184, 13.59683, 13.84193, 14.08713, 14.33243, 
    14.57783, 14.8233, 15.06886, 15.31449, 15.56018, 15.80594, 16.05175, 
    16.29761, 16.54351, 16.78944, 17.03541, 17.2814, 17.52741, 17.77343, 
    18.01946, 18.26549, 18.51151, 18.75751, 19.0035, 19.24946, 19.49539, 
    19.74129, 19.98714, 20.23294, 20.47869, 20.72437, 20.96999, 21.21553, 
    21.461, 21.70638, 21.95166, 22.19685, 22.44193, 22.68691, 22.93177, 
    23.1765, 23.42111, 23.66559, 23.90993, 24.15412, 24.39816, 24.64204, 
    24.88576, 25.12932, 25.37269, 25.61589, 25.85891, 26.10173, 26.34436, 
    26.58678, 26.829, 27.071, 27.31279, 27.55435, 27.79568, 28.03678, 
    28.27763, 28.51825, 28.75861, 28.99871, 29.23856, 29.47813, 29.71744, 
    29.95647, 30.19522, 30.43369, 30.67186, 30.90974, 31.14732, 31.38459, 
    31.62155, 31.8582, 32.09452, 32.33053, 32.5662, 32.80155, 33.03655, 
    33.27121, 33.50553, 33.7395, 33.97311, 34.20637, 34.43926, 34.67178, 
    34.90394, 35.13572, 35.36712, 35.59813, 35.82877, 36.05901, 36.28885, 
    36.5183, 36.74735, 36.97599, 37.20423, 37.43205, 37.65946, 37.88645, 
    38.11302, 38.33917, 38.56488, 38.79017, 39.01502, 39.23944, 39.46341, 
    39.68694, 39.91003, 40.13266, 40.35485, 40.57658, 40.79786, 41.01868, 
    41.23903, 41.45892, 41.67835, 41.8973, 42.11579, 42.3338, 42.55133, 
    42.76839, 42.98497, 43.20107, 43.41668, 43.63181, 43.84645, 44.0606, 
    44.27426, 44.48742, 44.70009, 44.91227, 45.12395, 45.33512, 45.5458, 
    45.75598, 45.96565, 46.17481, 46.38347, 46.59163, 46.79927, 47.0064, 
    47.21303, 47.41914, 47.62474, 47.82982, 48.03439, 48.23845, 48.44198, 
    48.645, 48.8475, 49.04949, 49.25095, 49.45189, 49.65232, 49.85222, 
    50.0516, 50.25046, 50.44879, 50.64661, 50.84389, 51.04066, 51.2369, 
    51.43262, 51.62782, 51.82248, 52.01663, 52.21025, 52.40334, 52.59592, 
    52.78796, 52.97948, 53.17048, 53.36095, 53.5509, 53.74033, 53.92923, 
    54.11761, 54.30547, 54.4928, 54.67961, 54.8659, 55.05166, 55.23691, 
    55.42163, 55.60583, 55.78952, 55.97269,
  -34.97403, -34.83418, -34.69394, -34.55329, -34.41224, -34.27078, 
    -34.12891, -33.98663, -33.84394, -33.70083, -33.55731, -33.41337, 
    -33.26902, -33.12424, -32.97905, -32.83342, -32.68738, -32.54091, 
    -32.39401, -32.24668, -32.09892, -31.95073, -31.8021, -31.65304, 
    -31.50354, -31.3536, -31.20322, -31.0524, -30.90113, -30.74942, 
    -30.59727, -30.44466, -30.29161, -30.1381, -29.98414, -29.82973, 
    -29.67486, -29.51954, -29.36375, -29.20751, -29.0508, -28.89363, -28.736, 
    -28.5779, -28.41933, -28.26029, -28.10078, -27.94081, -27.78035, 
    -27.61943, -27.45802, -27.29614, -27.13378, -26.97094, -26.80762, 
    -26.64382, -26.47953, -26.31476, -26.1495, -25.98375, -25.81751, 
    -25.65078, -25.48356, -25.31585, -25.14764, -24.97894, -24.80974, 
    -24.64004, -24.46984, -24.29915, -24.12795, -23.95625, -23.78405, 
    -23.61134, -23.43812, -23.2644, -23.09017, -22.91544, -22.74019, 
    -22.56443, -22.38816, -22.21138, -22.03409, -21.85628, -21.67795, 
    -21.49911, -21.31975, -21.13988, -20.95949, -20.77857, -20.59714, 
    -20.41519, -20.23271, -20.04972, -19.8662, -19.68216, -19.49759, 
    -19.3125, -19.12689, -18.94075, -18.75409, -18.56689, -18.37918, 
    -18.19093, -18.00216, -17.81286, -17.62304, -17.43268, -17.2418, 
    -17.05039, -16.85845, -16.66598, -16.47298, -16.27946, -16.08541, 
    -15.89082, -15.69571, -15.50007, -15.3039, -15.10721, -14.90998, 
    -14.71223, -14.51395, -14.31514, -14.11581, -13.91595, -13.71556, 
    -13.51465, -13.31321, -13.11125, -12.90876, -12.70575, -12.50222, 
    -12.29817, -12.0936, -11.8885, -11.68289, -11.47676, -11.27011, 
    -11.06295, -10.85527, -10.64707, -10.43836, -10.22915, -10.01941, 
    -9.809175, -9.598428, -9.387174, -9.175415, -8.963152, -8.750386, 
    -8.537121, -8.323356, -8.109094, -7.894336, -7.679085, -7.463341, 
    -7.247108, -7.030386, -6.813179, -6.595487, -6.377314, -6.15866, 
    -5.939529, -5.719923, -5.499843, -5.279293, -5.058274, -4.83679, 
    -4.614842, -4.392434, -4.169568, -3.946246, -3.722472, -3.498248, 
    -3.273577, -3.048462, -2.822906, -2.596912, -2.370483, -2.143622, 
    -1.916333, -1.688618, -1.460481, -1.231925, -1.002954, -0.773571, 
    -0.5437796, -0.3135835, -0.08298621, 0.1480085, 0.379397, 0.6111754, 
    0.84334, 1.075887, 1.308812, 1.542111, 1.77578, 2.009816, 2.244213, 
    2.478968, 2.714077, 2.949534, 3.185337, 3.421479, 3.657958, 3.894768, 
    4.131904, 4.369363, 4.607139, 4.845228, 5.083624, 5.322324, 5.561323, 
    5.800614, 6.040195, 6.280058, 6.5202, 6.760615, 7.001299, 7.242245, 
    7.483449, 7.724906, 7.96661, 8.208556, 8.450739, 8.693153, 8.935793, 
    9.178652, 9.421726, 9.66501, 9.908497, 10.15218, 10.39606, 10.64012, 
    10.88437, 11.12879, 11.37338, 11.61813, 11.86304, 12.1081, 12.35331, 
    12.59866, 12.84414, 13.08975, 13.33548, 13.58133, 13.82729, 14.07335, 
    14.31951, 14.56577, 14.81211, 15.05852, 15.30502, 15.55158, 15.7982, 
    16.04487, 16.2916, 16.53837, 16.78517, 17.03201, 17.27887, 17.52574, 
    17.77263, 18.01953, 18.26642, 18.51331, 18.76019, 19.00704, 19.25387, 
    19.50067, 19.74743, 19.99415, 20.24082, 20.48743, 20.73398, 20.98046, 
    21.22687, 21.47319, 21.71943, 21.96558, 22.21162, 22.45757, 22.7034, 
    22.94911, 23.1947, 23.44016, 23.68549, 23.93067, 24.17571, 24.4206, 
    24.66532, 24.90989, 25.15428, 25.39849, 25.64253, 25.88638, 26.13003, 
    26.37349, 26.61674, 26.85978, 27.1026, 27.34521, 27.58759, 27.82973, 
    28.07164, 28.3133, 28.55472, 28.79589, 29.03679, 29.27743, 29.51781, 
    29.7579, 29.99772, 30.23726, 30.4765, 30.71545, 30.95411, 31.19246, 
    31.43049, 31.66822, 31.90563, 32.14272, 32.37947, 32.6159, 32.85199, 
    33.08773, 33.32314, 33.55819, 33.79289, 34.02723, 34.26121, 34.49482, 
    34.72806, 34.96092, 35.19341, 35.42551, 35.65723, 35.88856, 36.11949, 
    36.35003, 36.58015, 36.80988, 37.0392, 37.26811, 37.4966, 37.72467, 
    37.95232, 38.17953, 38.40633, 38.63269, 38.85862, 39.0841, 39.30915, 
    39.53374, 39.7579, 39.9816, 40.20485, 40.42765, 40.64998, 40.87186, 
    41.09327, 41.31421, 41.53469, 41.75469, 41.97422, 42.19328, 42.41186, 
    42.62996, 42.84757, 43.0647, 43.28135, 43.4975, 43.71317, 43.92834, 
    44.14302, 44.3572, 44.57089, 44.78408, 44.99676, 45.20895, 45.42062, 
    45.6318, 45.84246, 46.05262, 46.26228, 46.47141, 46.68004, 46.88815, 
    47.09575, 47.30283, 47.5094, 47.71545, 47.92098, 48.12599, 48.33048, 
    48.53445, 48.7379, 48.94083, 49.14323, 49.34511, 49.54646, 49.74729, 
    49.94759, 50.14737, 50.34662, 50.54535, 50.74355, 50.94121, 51.13836, 
    51.33497, 51.53105, 51.72661, 51.92164, 52.11613, 52.31011, 52.50355, 
    52.69646, 52.88885, 53.0807, 53.27203, 53.46283, 53.6531, 53.84284, 
    54.03206, 54.22075, 54.40891, 54.59654, 54.78365, 54.97023, 55.15628, 
    55.34182, 55.52682, 55.7113, 55.89526, 56.0787,
  -35.09268, -34.95282, -34.81255, -34.67187, -34.53078, -34.38929, 
    -34.24739, -34.10507, -33.96234, -33.81919, -33.67564, -33.53165, 
    -33.38725, -33.24243, -33.09719, -32.95152, -32.80542, -32.65889, 
    -32.51194, -32.36455, -32.21673, -32.06848, -31.91979, -31.77066, 
    -31.62109, -31.47108, -31.32063, -31.16974, -31.0184, -30.86661, 
    -30.71437, -30.56168, -30.40854, -30.25495, -30.1009, -29.9464, 
    -29.79144, -29.63601, -29.48013, -29.32378, -29.16697, -29.0097, 
    -28.85195, -28.69374, -28.53506, -28.37591, -28.21628, -28.05618, 
    -27.89561, -27.73455, -27.57302, -27.41101, -27.24851, -27.08554, 
    -26.92208, -26.75813, -26.59369, -26.42877, -26.26336, -26.09746, 
    -25.93106, -25.76418, -25.59679, -25.42891, -25.26054, -25.09166, 
    -24.92229, -24.75241, -24.58203, -24.41115, -24.23977, -24.06788, 
    -23.89548, -23.72257, -23.54916, -23.37523, -23.2008, -23.02585, 
    -22.85039, -22.67441, -22.49792, -22.32092, -22.1434, -21.96536, 
    -21.7868, -21.60772, -21.42812, -21.248, -21.06736, -20.88619, -20.7045, 
    -20.52229, -20.33955, -20.15629, -19.9725, -19.78819, -19.60334, 
    -19.41797, -19.23207, -19.04564, -18.85868, -18.67119, -18.48317, 
    -18.29462, -18.10554, -17.91593, -17.72579, -17.53511, -17.3439, 
    -17.15216, -16.95989, -16.76708, -16.57374, -16.37987, -16.18546, 
    -15.99053, -15.79505, -15.59905, -15.40251, -15.20544, -15.00784, 
    -14.80971, -14.61104, -14.41185, -14.21212, -14.01186, -13.81107, 
    -13.60975, -13.4079, -13.20552, -13.00262, -12.79918, -12.59522, 
    -12.39073, -12.18572, -11.98018, -11.77412, -11.56754, -11.36043, 
    -11.15281, -10.94466, -10.73599, -10.52681, -10.31711, -10.10689, 
    -9.896166, -9.684923, -9.47317, -9.260907, -9.048135, -8.834857, 
    -8.621073, -8.406785, -8.191996, -7.976706, -7.760918, -7.544633, 
    -7.327853, -7.110581, -6.892817, -6.674565, -6.455827, -6.236604, 
    -6.016898, -5.796712, -5.576049, -5.35491, -5.133299, -4.911217, 
    -4.688667, -4.465652, -4.242174, -4.018236, -3.793841, -3.568991, 
    -3.343691, -3.117941, -2.891746, -2.665108, -2.438031, -2.210518, 
    -1.982571, -1.754195, -1.525392, -1.296166, -1.06652, -0.836458, 
    -0.6059834, -0.3750996, -0.1438104, 0.08788048, 0.3199694, 0.5524523, 
    0.7853256, 1.018585, 1.252227, 1.486247, 1.720642, 1.955406, 2.190536, 
    2.426028, 2.661878, 2.89808, 3.134631, 3.371526, 3.60876, 3.846329, 
    4.084229, 4.322454, 4.561001, 4.799864, 5.039038, 5.278519, 5.518301, 
    5.75838, 5.998751, 6.239408, 6.480348, 6.721563, 6.96305, 7.204803, 
    7.446816, 7.689085, 7.931604, 8.174368, 8.417371, 8.660607, 8.904073, 
    9.14776, 9.391665, 9.635782, 9.880105, 10.12463, 10.36935, 10.61425, 
    10.85934, 11.10461, 11.35004, 11.59565, 11.84141, 12.08733, 12.33339, 
    12.57959, 12.82594, 13.07241, 13.319, 13.56571, 13.81254, 14.05946, 
    14.30649, 14.55361, 14.80082, 15.04811, 15.29547, 15.5429, 15.79039, 
    16.03794, 16.28554, 16.53318, 16.78086, 17.02857, 17.27631, 17.52406, 
    17.77183, 18.0196, 18.26737, 18.51513, 18.76288, 19.01061, 19.25832, 
    19.50599, 19.75363, 20.00122, 20.24876, 20.49624, 20.74366, 20.99101, 
    21.23829, 21.48548, 21.73259, 21.9796, 22.22651, 22.47332, 22.72001, 
    22.96659, 23.21304, 23.45936, 23.70554, 23.95158, 24.19748, 24.44321, 
    24.68879, 24.9342, 25.17944, 25.4245, 25.66938, 25.91406, 26.15856, 
    26.40285, 26.64693, 26.8908, 27.13445, 27.37788, 27.62108, 27.86405, 
    28.10678, 28.34925, 28.59148, 28.83346, 29.07517, 29.31661, 29.55778, 
    29.79868, 30.03929, 30.27962, 30.51965, 30.75938, 30.99882, 31.23794, 
    31.47675, 31.71525, 31.95342, 32.19127, 32.42879, 32.66597, 32.90281, 
    33.13931, 33.37545, 33.61125, 33.84668, 34.08175, 34.31646, 34.5508, 
    34.78476, 35.01834, 35.25154, 35.48435, 35.71677, 35.9488, 36.18042, 
    36.41165, 36.64247, 36.87288, 37.10287, 37.33245, 37.56161, 37.79035, 
    38.01866, 38.24654, 38.47398, 38.70099, 38.92756, 39.15368, 39.37936, 
    39.60459, 39.82937, 40.05369, 40.27755, 40.50096, 40.7239, 40.94638, 
    41.16838, 41.38992, 41.61098, 41.83157, 42.05169, 42.27131, 42.49046, 
    42.70912, 42.9273, 43.14498, 43.36218, 43.57888, 43.79509, 44.0108, 
    44.22601, 44.44072, 44.65492, 44.86863, 45.08183, 45.29452, 45.5067, 
    45.71837, 45.92953, 46.14018, 46.35032, 46.55993, 46.76904, 46.97762, 
    47.18568, 47.39323, 47.60025, 47.80676, 48.01273, 48.21819, 48.42311, 
    48.62752, 48.8314, 49.03475, 49.23757, 49.43987, 49.64163, 49.84286, 
    50.04357, 50.24375, 50.44339, 50.64251, 50.84109, 51.03913, 51.23665, 
    51.43364, 51.63009, 51.82601, 52.0214, 52.21625, 52.41057, 52.60436, 
    52.79762, 52.99034, 53.18253, 53.37418, 53.56531, 53.7559, 53.94596, 
    54.13549, 54.32449, 54.51295, 54.70089, 54.88829, 55.07516, 55.26151, 
    55.44733, 55.63261, 55.81738, 56.00161, 56.18531,
  -35.21182, -35.07193, -34.93163, -34.79093, -34.64981, -34.50829, 
    -34.36636, -34.22401, -34.08124, -33.93806, -33.79446, -33.65044, 
    -33.50599, -33.36113, -33.21584, -33.07012, -32.92397, -32.77739, 
    -32.63038, -32.48294, -32.33506, -32.18675, -32.03799, -31.8888, 
    -31.73917, -31.58909, -31.43857, -31.2876, -31.13619, -30.98432, 
    -30.83201, -30.67924, -30.52601, -30.37234, -30.2182, -30.0636, 
    -29.90855, -29.75303, -29.59705, -29.44061, -29.28369, -29.12631, 
    -28.96846, -28.81014, -28.65135, -28.49208, -28.33234, -28.17212, 
    -28.01142, -27.85024, -27.68858, -27.52644, -27.36381, -27.2007, 
    -27.0371, -26.87301, -26.70843, -26.54336, -26.3778, -26.21174, 
    -26.04519, -25.87815, -25.7106, -25.54256, -25.37401, -25.20497, 
    -25.03542, -24.86537, -24.69481, -24.52374, -24.35217, -24.18009, 
    -24.0075, -23.8344, -23.66078, -23.48666, -23.31202, -23.13686, 
    -22.96119, -22.78499, -22.60829, -22.43106, -22.25331, -22.07504, 
    -21.89624, -21.71693, -21.53709, -21.35672, -21.17583, -20.99442, 
    -20.81247, -20.63, -20.447, -20.26347, -20.07941, -19.89482, -19.7097, 
    -19.52405, -19.33786, -19.15114, -18.96389, -18.7761, -18.58778, 
    -18.39893, -18.20954, -18.01961, -17.82915, -17.63815, -17.44662, 
    -17.25454, -17.06194, -16.86879, -16.67511, -16.48089, -16.28613, 
    -16.09084, -15.89501, -15.69864, -15.50174, -15.30429, -15.10632, 
    -14.9078, -14.70875, -14.50916, -14.30904, -14.10838, -13.90719, 
    -13.70546, -13.5032, -13.3004, -13.09707, -12.89321, -12.68882, -12.4839, 
    -12.27845, -12.07246, -11.86595, -11.65891, -11.45135, -11.24326, 
    -11.03464, -10.82551, -10.61584, -10.40566, -10.19496, -9.98374, 
    -9.772001, -9.559747, -9.346978, -9.133696, -8.919902, -8.705598, 
    -8.490786, -8.275467, -8.059643, -7.843316, -7.626487, -7.409159, 
    -7.191333, -6.973011, -6.754197, -6.53489, -6.315094, -6.094812, 
    -5.874044, -5.652795, -5.431065, -5.208857, -4.986175, -4.763019, 
    -4.539394, -4.315301, -4.090744, -3.865725, -3.640246, -3.414312, 
    -3.187925, -2.961087, -2.733802, -2.506073, -2.277904, -2.049296, 
    -1.820254, -1.590782, -1.360881, -1.130557, -0.8998119, -0.6686497, 
    -0.4370742, -0.2050888, 0.0273026, 0.2600962, 0.4932882, 0.7268746, 
    0.9608517, 1.195215, 1.429961, 1.665085, 1.900584, 2.136452, 2.372685, 
    2.609281, 2.846232, 3.083537, 3.321189, 3.559184, 3.797518, 4.036187, 
    4.275185, 4.514507, 4.754149, 4.994106, 5.234373, 5.474945, 5.715817, 
    5.956985, 6.198442, 6.440184, 6.682205, 6.924501, 7.167066, 7.409894, 
    7.652982, 7.896322, 8.13991, 8.383739, 8.627805, 8.872103, 9.116625, 
    9.361367, 9.606323, 9.851488, 10.09686, 10.34242, 10.58817, 10.83411, 
    11.08023, 11.32652, 11.57298, 11.81961, 12.06638, 12.31331, 12.56038, 
    12.80758, 13.05492, 13.30239, 13.54997, 13.79766, 14.04546, 14.29336, 
    14.54136, 14.78944, 15.03761, 15.28585, 15.53416, 15.78253, 16.03096, 
    16.27944, 16.52796, 16.77652, 17.02511, 17.27373, 17.52237, 17.77101, 
    18.01967, 18.26832, 18.51697, 18.7656, 19.01421, 19.2628, 19.51135, 
    19.75987, 20.00834, 20.25676, 20.50513, 20.75342, 21.00165, 21.24981, 
    21.49788, 21.74586, 21.99374, 22.24153, 22.4892, 22.73677, 22.98421, 
    23.23153, 23.47871, 23.72576, 23.97266, 24.21942, 24.46601, 24.71245, 
    24.95871, 25.2048, 25.45071, 25.69644, 25.94197, 26.18731, 26.43244, 
    26.67736, 26.92207, 27.16656, 27.41082, 27.65485, 27.89864, 28.14219, 
    28.38549, 28.62853, 28.87132, 29.11384, 29.3561, 29.59807, 29.83977, 
    30.08118, 30.3223, 30.56313, 30.80365, 31.04387, 31.28378, 31.52337, 
    31.76264, 32.00159, 32.2402, 32.47849, 32.71643, 32.95403, 33.19127, 
    33.42817, 33.66471, 33.90088, 34.13669, 34.37213, 34.6072, 34.84188, 
    35.07619, 35.3101, 35.54362, 35.77676, 36.00948, 36.24181, 36.47373, 
    36.70524, 36.93634, 37.16702, 37.39728, 37.62711, 37.85651, 38.08549, 
    38.31403, 38.54213, 38.76978, 38.997, 39.22377, 39.45008, 39.67595, 
    39.90135, 40.1263, 40.35078, 40.5748, 40.79835, 41.02143, 41.24404, 
    41.46617, 41.68782, 41.909, 42.12969, 42.3499, 42.56961, 42.78884, 
    43.00758, 43.22582, 43.44357, 43.66082, 43.87757, 44.09381, 44.30956, 
    44.5248, 44.73953, 44.95375, 45.16747, 45.38067, 45.59336, 45.80553, 
    46.01719, 46.22832, 46.43895, 46.64904, 46.85862, 47.06768, 47.27621, 
    47.48422, 47.6917, 47.89865, 48.10508, 48.31098, 48.51635, 48.72119, 
    48.9255, 49.12927, 49.33252, 49.53522, 49.7374, 49.93905, 50.14016, 
    50.34073, 50.54077, 50.74027, 50.93924, 51.13767, 51.33556, 51.53292, 
    51.72974, 51.92602, 52.12177, 52.31698, 52.51165, 52.70578, 52.89938, 
    53.09244, 53.28496, 53.47695, 53.6684, 53.85931, 54.04969, 54.23953, 
    54.42884, 54.61761, 54.80584, 54.99355, 55.18071, 55.36735, 55.55345, 
    55.73902, 55.92406, 56.10856, 56.29254,
  -35.33144, -35.19153, -35.05121, -34.91048, -34.76934, -34.62779, 
    -34.48582, -34.34344, -34.20064, -34.05742, -33.91378, -33.76973, 
    -33.62524, -33.48033, -33.33499, -33.18923, -33.04303, -32.8964, 
    -32.74934, -32.60184, -32.45391, -32.30554, -32.15673, -32.00747, 
    -31.85777, -31.70763, -31.55704, -31.406, -31.25451, -31.10257, 
    -30.95018, -30.79733, -30.64402, -30.49026, -30.33604, -30.18135, 
    -30.02621, -29.8706, -29.71452, -29.55798, -29.40096, -29.24348, 
    -29.08553, -28.9271, -28.76819, -28.60881, -28.44895, -28.28861, 
    -28.12779, -27.96649, -27.8047, -27.64243, -27.47967, -27.31643, 
    -27.15269, -26.98846, -26.82374, -26.65853, -26.49282, -26.32661, 
    -26.1599, -25.9927, -25.82499, -25.65679, -25.48808, -25.31886, 
    -25.14914, -24.97891, -24.80817, -24.63693, -24.46517, -24.2929, 
    -24.12012, -23.94682, -23.77301, -23.59868, -23.42383, -23.24847, 
    -23.07258, -22.89618, -22.71925, -22.5418, -22.36382, -22.18532, 
    -22.0063, -21.82675, -21.64667, -21.46606, -21.28492, -21.10325, 
    -20.92105, -20.73832, -20.55506, -20.37127, -20.18694, -20.00207, 
    -19.81667, -19.63074, -19.44427, -19.25726, -19.06971, -18.88163, 
    -18.69301, -18.50385, -18.31415, -18.12391, -17.93313, -17.74181, 
    -17.54995, -17.35755, -17.1646, -16.97112, -16.7771, -16.58253, 
    -16.38742, -16.19177, -15.99558, -15.79885, -15.60157, -15.40376, 
    -15.2054, -15.00651, -14.80707, -14.60709, -14.40657, -14.20551, 
    -14.00391, -13.80178, -13.5991, -13.39589, -13.19214, -12.98785, 
    -12.78303, -12.57767, -12.37177, -12.16535, -11.95838, -11.75089, 
    -11.54287, -11.33431, -11.12523, -10.91561, -10.70547, -10.49481, 
    -10.28362, -10.0719, -9.859668, -9.646911, -9.433634, -9.219839, 
    -9.005528, -8.790703, -8.575363, -8.359512, -8.143152, -7.926284, 
    -7.708909, -7.49103, -7.272648, -7.053766, -6.834386, -6.61451, 
    -6.394139, -6.173277, -5.951925, -5.730086, -5.507761, -5.284955, 
    -5.061668, -4.837905, -4.613666, -4.388956, -4.163775, -3.938129, 
    -3.712019, -3.485448, -3.258419, -3.030935, -2.802999, -2.574615, 
    -2.345785, -2.116513, -1.886802, -1.656656, -1.426077, -1.19507, 
    -0.963638, -0.7317842, -0.4995126, -0.2668267, -0.03373052, 0.1997723, 
    0.4336777, 0.667982, 0.9026809, 1.137771, 1.373247, 1.609106, 1.845343, 
    2.081954, 2.318934, 2.55628, 2.793987, 3.032049, 3.270464, 3.509226, 
    3.74833, 3.987772, 4.227548, 4.467651, 4.708078, 4.948824, 5.189883, 
    5.43125, 5.672921, 5.914891, 6.157154, 6.399704, 6.642538, 6.885649, 
    7.129032, 7.372682, 7.616593, 7.86076, 8.105178, 8.34984, 8.594742, 
    8.839878, 9.085241, 9.330827, 9.576629, 9.822641, 10.06886, 10.31528, 
    10.56189, 10.80868, 11.05566, 11.30282, 11.55014, 11.79763, 12.04527, 
    12.29307, 12.54101, 12.78909, 13.0373, 13.28564, 13.53409, 13.78267, 
    14.03135, 14.28013, 14.52901, 14.77797, 15.02702, 15.27615, 15.52534, 
    15.7746, 16.02392, 16.27328, 16.5227, 16.77214, 17.02163, 17.27113, 
    17.52066, 17.77019, 18.01974, 18.26928, 18.51881, 18.76834, 19.01784, 
    19.26731, 19.51676, 19.76616, 20.01552, 20.26483, 20.51408, 20.76326, 
    21.01238, 21.26141, 21.51037, 21.75923, 22.008, 22.25666, 22.50521, 
    22.75365, 23.00197, 23.25017, 23.49822, 23.74614, 23.99391, 24.24153, 
    24.48899, 24.73629, 24.98342, 25.23037, 25.47713, 25.72371, 25.9701, 
    26.21629, 26.46227, 26.70803, 26.95359, 27.19891, 27.44401, 27.68888, 
    27.9335, 28.17788, 28.42201, 28.66588, 28.90948, 29.15283, 29.39589, 
    29.63868, 29.88119, 30.1234, 30.36533, 30.60695, 30.84827, 31.08928, 
    31.32998, 31.57035, 31.8104, 32.05013, 32.28952, 32.52856, 32.76727, 
    33.00563, 33.24364, 33.48129, 33.71858, 33.9555, 34.19205, 34.42823, 
    34.66403, 34.89944, 35.13447, 35.36911, 35.60335, 35.83719, 36.07063, 
    36.30366, 36.53628, 36.76849, 37.00027, 37.23164, 37.46258, 37.69309, 
    37.92317, 38.15281, 38.38201, 38.61077, 38.83908, 39.06695, 39.29436, 
    39.52132, 39.74782, 39.97385, 40.19942, 40.42453, 40.64917, 40.87333, 
    41.09702, 41.32023, 41.54296, 41.76521, 41.98697, 42.20825, 42.42903, 
    42.64932, 42.86912, 43.08842, 43.30722, 43.52553, 43.74333, 43.96062, 
    44.17741, 44.39369, 44.60946, 44.82472, 45.03946, 45.25369, 45.4674, 
    45.6806, 45.89328, 46.10543, 46.31706, 46.52817, 46.73875, 46.94881, 
    47.15834, 47.36734, 47.57581, 47.78375, 47.99116, 48.19804, 48.40438, 
    48.61019, 48.81546, 49.0202, 49.2244, 49.42807, 49.6312, 49.83379, 
    50.03584, 50.23735, 50.43833, 50.63876, 50.83865, 51.03801, 51.23682, 
    51.43509, 51.63282, 51.83001, 52.02665, 52.22276, 52.41832, 52.61334, 
    52.80782, 53.00176, 53.19516, 53.38802, 53.58033, 53.77211, 53.96334, 
    54.15403, 54.34419, 54.53381, 54.72288, 54.91142, 55.09941, 55.28688, 
    55.4738, 55.66019, 55.84604, 56.03135, 56.21613, 56.40038,
  -35.45156, -35.31162, -35.17128, -35.03053, -34.88936, -34.74778, 
    -34.60579, -34.46337, -34.32054, -34.17729, -34.03362, -33.88952, 
    -33.74499, -33.60004, -33.45466, -33.30885, -33.16261, -33.01593, 
    -32.86882, -32.72127, -32.57328, -32.42485, -32.27598, -32.12666, 
    -31.9769, -31.82669, -31.67604, -31.52493, -31.37337, -31.22136, 
    -31.06889, -30.91596, -30.76258, -30.60873, -30.45442, -30.29965, 
    -30.14442, -29.98871, -29.83254, -29.6759, -29.51879, -29.36121, 
    -29.20315, -29.04461, -28.8856, -28.7261, -28.56613, -28.40568, 
    -28.24474, -28.08331, -27.9214, -27.759, -27.59611, -27.43273, -27.26886, 
    -27.10449, -26.93963, -26.77427, -26.60841, -26.44205, -26.2752, 
    -26.10784, -25.93997, -25.7716, -25.60273, -25.43334, -25.26345, 
    -25.09305, -24.92213, -24.75071, -24.57876, -24.40631, -24.23333, 
    -24.05984, -23.88583, -23.7113, -23.53625, -23.36068, -23.18459, 
    -23.00797, -22.83082, -22.65315, -22.47495, -22.29622, -22.11696, 
    -21.93717, -21.75686, -21.576, -21.39462, -21.2127, -21.03025, -20.84726, 
    -20.66374, -20.47968, -20.29508, -20.10994, -19.92426, -19.73805, 
    -19.55129, -19.364, -19.17616, -18.98778, -18.79885, -18.60939, 
    -18.41938, -18.22883, -18.03773, -17.84609, -17.6539, -17.46117, 
    -17.26789, -17.07407, -16.8797, -16.68479, -16.48933, -16.29333, 
    -16.09678, -15.89968, -15.70204, -15.50385, -15.30511, -15.10583, 
    -14.90601, -14.70564, -14.50472, -14.30326, -14.10126, -13.89872, 
    -13.69563, -13.49199, -13.28782, -13.0831, -12.87785, -12.67205, 
    -12.46571, -12.25884, -12.05143, -11.84348, -11.63499, -11.42597, 
    -11.21641, -11.00632, -10.7957, -10.58455, -10.37287, -10.16066, 
    -9.947928, -9.734667, -9.520881, -9.306572, -9.091742, -8.876392, 
    -8.660524, -8.444139, -8.227241, -8.009829, -7.791906, -7.573473, 
    -7.354534, -7.135089, -6.915141, -6.694692, -6.473744, -6.252299, 
    -6.03036, -5.807928, -5.585007, -5.361598, -5.137705, -4.91333, 
    -4.688475, -4.463143, -4.237338, -4.01106, -3.784315, -3.557103, 
    -3.329429, -3.101296, -2.872706, -2.643662, -2.414169, -2.184228, 
    -1.953844, -1.72302, -1.49176, -1.260066, -1.027942, -0.7953924, 
    -0.5624204, -0.3290298, -0.09522434, 0.1389921, 0.3736156, 0.6086421, 
    0.8440678, 1.079888, 1.3161, 1.552698, 1.789678, 2.027037, 2.264769, 
    2.502871, 2.741338, 2.980164, 3.219347, 3.45888, 3.69876, 3.938982, 
    4.17954, 4.42043, 4.661648, 4.903187, 5.145044, 5.387212, 5.629688, 
    5.872466, 6.11554, 6.358905, 6.602557, 6.846489, 7.090696, 7.335174, 
    7.579916, 7.824916, 8.07017, 8.315672, 8.561416, 8.807396, 9.053606, 
    9.300042, 9.546697, 9.793565, 10.04064, 10.28792, 10.53539, 10.78305, 
    11.0309, 11.27892, 11.52711, 11.77547, 12.02399, 12.27266, 12.52148, 
    12.77044, 13.01953, 13.26875, 13.51809, 13.76755, 14.01712, 14.26679, 
    14.51656, 14.76641, 15.01635, 15.26637, 15.51646, 15.76661, 16.01682, 
    16.26708, 16.51739, 16.76773, 17.01811, 17.26851, 17.51893, 17.76937, 
    18.01981, 18.27025, 18.52068, 18.7711, 19.0215, 19.27187, 19.52221, 
    19.77251, 20.02276, 20.27296, 20.52311, 20.77318, 21.02319, 21.27312, 
    21.52296, 21.77271, 22.02237, 22.27192, 22.52136, 22.77068, 23.01988, 
    23.26895, 23.51789, 23.76669, 24.01533, 24.26383, 24.51216, 24.76033, 
    25.00832, 25.25614, 25.50377, 25.75121, 25.99846, 26.2455, 26.49233, 
    26.73895, 26.98536, 27.23153, 27.47747, 27.72318, 27.96864, 28.21386, 
    28.45882, 28.70352, 28.94795, 29.19212, 29.436, 29.67961, 29.92293, 
    30.16596, 30.40869, 30.65112, 30.89323, 31.13504, 31.37653, 31.6177, 
    31.85853, 32.09904, 32.33921, 32.57903, 32.81851, 33.05764, 33.29641, 
    33.53482, 33.77286, 34.01053, 34.24783, 34.48475, 34.72129, 34.95744, 
    35.1932, 35.42856, 35.66352, 35.89808, 36.13224, 36.36597, 36.5993, 
    36.83221, 37.06469, 37.29675, 37.52837, 37.75956, 37.99032, 38.22063, 
    38.4505, 38.67992, 38.90889, 39.13741, 39.36547, 39.59307, 39.82021, 
    40.04689, 40.27309, 40.49882, 40.72408, 40.94886, 41.17315, 41.39697, 
    41.6203, 41.84315, 42.0655, 42.28736, 42.50873, 42.7296, 42.94997, 
    43.16983, 43.3892, 43.60806, 43.82641, 44.04425, 44.26159, 44.4784, 
    44.69471, 44.91049, 45.12576, 45.34051, 45.55473, 45.76844, 45.98161, 
    46.19427, 46.40639, 46.61799, 46.82906, 47.03959, 47.2496, 47.45907, 
    47.668, 47.8764, 48.08427, 48.2916, 48.49839, 48.70464, 48.91035, 
    49.11552, 49.32015, 49.52424, 49.72779, 49.93079, 50.13325, 50.33517, 
    50.53654, 50.73737, 50.93765, 51.13739, 51.33659, 51.53523, 51.73334, 
    51.93089, 52.1279, 52.32437, 52.52029, 52.71566, 52.91048, 53.10477, 
    53.2985, 53.49169, 53.68434, 53.87644, 54.06799, 54.25901, 54.44947, 
    54.6394, 54.82877, 55.01761, 55.20591, 55.39366, 55.58087, 55.76754, 
    55.95367, 56.13926, 56.32431, 56.50883,
  -35.57216, -35.43221, -35.29184, -35.15107, -35.00988, -34.86827, 
    -34.72625, -34.58381, -34.44094, -34.29766, -34.15395, -34.00982, 
    -33.86526, -33.72027, -33.57485, -33.42899, -33.2827, -33.13598, 
    -32.98882, -32.84122, -32.69318, -32.54469, -32.39576, -32.24639, 
    -32.09657, -31.9463, -31.79557, -31.6444, -31.49277, -31.34068, 
    -31.18814, -31.03514, -30.88167, -30.72775, -30.57336, -30.4185, 
    -30.26318, -30.10738, -29.95112, -29.79439, -29.63718, -29.47949, 
    -29.32133, -29.16269, -29.00357, -28.84397, -28.68388, -28.52331, 
    -28.36225, -28.20071, -28.03867, -27.87615, -27.71313, -27.54962, 
    -27.38561, -27.2211, -27.0561, -26.8906, -26.7246, -26.55809, -26.39108, 
    -26.22356, -26.05554, -25.88701, -25.71797, -25.54842, -25.37836, 
    -25.20778, -25.03669, -24.86509, -24.69296, -24.52032, -24.34715, 
    -24.17347, -23.99927, -23.82454, -23.64928, -23.47351, -23.2972, 
    -23.12037, -22.943, -22.76511, -22.58669, -22.40773, -22.22824, 
    -22.04822, -21.86766, -21.68657, -21.50494, -21.32277, -21.14007, 
    -20.95682, -20.77304, -20.58871, -20.40384, -20.21844, -20.03248, 
    -19.84599, -19.65895, -19.47136, -19.28323, -19.09455, -18.90533, 
    -18.71556, -18.52524, -18.33437, -18.14296, -17.951, -17.75849, 
    -17.56542, -17.37181, -17.17765, -16.98294, -16.78768, -16.59187, 
    -16.39551, -16.1986, -16.00114, -15.80312, -15.60456, -15.40545, 
    -15.20579, -15.00558, -14.80481, -14.6035, -14.40164, -14.19923, 
    -13.99628, -13.79277, -13.58872, -13.38412, -13.17898, -12.97329, 
    -12.76705, -12.56027, -12.35295, -12.14508, -11.93667, -11.72773, 
    -11.51824, -11.30821, -11.09764, -10.88654, -10.6749, -10.46273, 
    -10.25003, -10.03679, -9.823022, -9.608726, -9.3939, -9.17855, -8.962673, 
    -8.746275, -8.529355, -8.311915, -8.093957, -7.875484, -7.656496, 
    -7.436996, -7.216986, -6.996467, -6.775443, -6.553914, -6.331884, 
    -6.109355, -5.886328, -5.662807, -5.438794, -5.214292, -4.989301, 
    -4.763827, -4.537871, -4.311436, -4.084525, -3.85714, -3.629285, 
    -3.400962, -3.172175, -2.942927, -2.713221, -2.48306, -2.252447, 
    -2.021386, -1.789881, -1.557934, -1.325549, -1.09273, -0.85948, 
    -0.6258033, -0.3917035, -0.1571844, 0.07775015, 0.3130962, 0.5488497, 
    0.7850067, 1.021563, 1.258514, 1.495857, 1.733586, 1.971697, 2.210186, 
    2.449049, 2.68828, 2.927876, 3.167831, 3.408142, 3.648803, 3.889809, 
    4.131156, 4.372839, 4.614852, 4.857192, 5.099852, 5.342827, 5.586113, 
    5.829705, 6.073596, 6.317782, 6.562258, 6.807017, 7.052055, 7.297367, 
    7.542945, 7.788785, 8.034883, 8.281229, 8.527822, 8.774652, 9.021717, 
    9.26901, 9.516523, 9.764253, 10.01219, 10.26034, 10.50868, 10.75721, 
    11.00593, 11.25483, 11.5039, 11.75314, 12.00253, 12.25209, 12.50179, 
    12.75164, 13.00162, 13.25173, 13.50196, 13.75231, 14.00277, 14.25334, 
    14.504, 14.75476, 15.00559, 15.25651, 15.5075, 15.75855, 16.00966, 
    16.26083, 16.51204, 16.76328, 17.01456, 17.26587, 17.5172, 17.76854, 
    18.01988, 18.27122, 18.52256, 18.77388, 19.02518, 19.27646, 19.5277, 
    19.77891, 20.03006, 20.28116, 20.53221, 20.78319, 21.03409, 21.28492, 
    21.53565, 21.7863, 22.03685, 22.2873, 22.53763, 22.78784, 23.03793, 
    23.28789, 23.53772, 23.7874, 24.03693, 24.2863, 24.53551, 24.78456, 
    25.03343, 25.28212, 25.53062, 25.77893, 26.02704, 26.27495, 26.52264, 
    26.77012, 27.01738, 27.26441, 27.5112, 27.75776, 28.00406, 28.25012, 
    28.49592, 28.74146, 28.98672, 29.23172, 29.47643, 29.72086, 29.965, 
    30.20885, 30.45239, 30.69563, 30.93855, 31.18116, 31.42345, 31.66541, 
    31.90704, 32.14834, 32.38929, 32.62989, 32.87015, 33.11005, 33.34959, 
    33.58876, 33.82756, 34.06599, 34.30404, 34.54171, 34.77899, 35.01588, 
    35.25238, 35.48847, 35.72416, 35.95944, 36.19431, 36.42876, 36.6628, 
    36.8964, 37.12959, 37.36234, 37.59465, 37.82653, 38.05796, 38.28896, 
    38.5195, 38.74959, 38.97922, 39.2084, 39.43711, 39.66536, 39.89314, 
    40.12045, 40.34729, 40.57365, 40.79953, 41.02493, 41.24984, 41.47426, 
    41.6982, 41.92164, 42.14459, 42.36704, 42.58899, 42.81044, 43.03138, 
    43.25182, 43.47175, 43.69117, 43.91008, 44.12847, 44.34634, 44.5637, 
    44.78054, 44.99686, 45.21265, 45.42792, 45.64266, 45.85687, 46.07056, 
    46.28371, 46.49633, 46.70842, 46.91997, 47.13099, 47.34147, 47.55141, 
    47.76081, 47.96968, 48.178, 48.38578, 48.59302, 48.79971, 49.00586, 
    49.21146, 49.41652, 49.62103, 49.825, 50.02842, 50.23129, 50.43361, 
    50.63538, 50.83661, 51.03728, 51.23741, 51.43698, 51.63601, 51.83448, 
    52.03241, 52.22978, 52.42661, 52.62288, 52.81861, 53.01378, 53.2084, 
    53.40248, 53.596, 53.78897, 53.9814, 54.17327, 54.3646, 54.55538, 
    54.74561, 54.9353, 55.12444, 55.31303, 55.50107, 55.68857, 55.87552, 
    56.06194, 56.2478, 56.43312, 56.6179,
  -35.69325, -35.55328, -35.4129, -35.2721, -35.13089, -34.98927, -34.84722, 
    -34.70475, -34.56186, -34.41854, -34.2748, -34.13063, -33.98604, 
    -33.84101, -33.69555, -33.54966, -33.40332, -33.25655, -33.10934, 
    -32.9617, -32.8136, -32.66507, -32.51608, -32.36665, -32.21677, 
    -32.06643, -31.91565, -31.76441, -31.61271, -31.46055, -31.30794, 
    -31.15486, -31.00132, -30.84732, -30.69284, -30.5379, -30.38249, 
    -30.22661, -30.07026, -29.91343, -29.75612, -29.59834, -29.44008, 
    -29.28133, -29.12211, -28.9624, -28.8022, -28.64152, -28.48034, 
    -28.31868, -28.15652, -27.99387, -27.83073, -27.66708, -27.50294, 
    -27.3383, -27.17316, -27.00752, -26.84137, -26.67472, -26.50756, 
    -26.33989, -26.17171, -26.00302, -25.83382, -25.6641, -25.49387, 
    -25.32312, -25.15186, -24.98007, -24.80776, -24.63494, -24.46159, 
    -24.28771, -24.11331, -23.93838, -23.76293, -23.58694, -23.41043, 
    -23.23338, -23.05581, -22.87769, -22.69905, -22.51987, -22.34015, 
    -22.15989, -21.9791, -21.79776, -21.61589, -21.43347, -21.25051, 
    -21.06701, -20.88297, -20.69838, -20.51324, -20.32756, -20.14133, 
    -19.95456, -19.76723, -19.57936, -19.39093, -19.20196, -19.01244, 
    -18.82236, -18.63173, -18.44056, -18.24883, -18.05654, -17.8637, 
    -17.67031, -17.47637, -17.28187, -17.08681, -16.89121, -16.69505, 
    -16.49833, -16.30106, -16.10323, -15.90485, -15.70591, -15.50642, 
    -15.30637, -15.10577, -14.90462, -14.70291, -14.50065, -14.29784, 
    -14.09447, -13.89055, -13.68608, -13.48105, -13.27548, -13.06935, 
    -12.86268, -12.65545, -12.44768, -12.23936, -12.03049, -11.82108, 
    -11.61112, -11.40062, -11.18958, -10.97799, -10.76587, -10.5532, -10.34, 
    -10.12626, -9.911983, -9.697173, -9.481831, -9.265957, -9.049553, 
    -8.832622, -8.615164, -8.397181, -8.178676, -7.959649, -7.740103, 
    -7.52004, -7.299462, -7.078371, -6.856769, -6.634657, -6.412039, 
    -6.188917, -5.965293, -5.741169, -5.516548, -5.291432, -5.065825, 
    -4.839728, -4.613144, -4.386076, -4.158527, -3.930501, -3.701998, 
    -3.473024, -3.24358, -3.01367, -2.783297, -2.552465, -2.321176, 
    -2.089434, -1.857243, -1.624606, -1.391526, -1.158007, -0.9240526, 
    -0.6896669, -0.4548536, -0.2196163, 0.01604087, 0.2521141, 0.4885992, 
    0.7254923, 0.9627891, 1.200485, 1.438577, 1.677059, 1.915928, 2.15518, 
    2.394808, 2.63481, 2.87518, 3.115914, 3.357007, 3.598454, 3.840251, 
    4.082392, 4.324872, 4.567688, 4.810833, 5.054302, 5.29809, 5.542193, 
    5.786604, 6.031319, 6.276332, 6.521638, 6.767231, 7.013106, 7.259257, 
    7.505678, 7.752365, 7.99931, 8.24651, 8.493957, 8.741646, 8.989572, 
    9.237726, 9.486106, 9.734704, 9.983515, 10.23253, 10.48175, 10.73116, 
    10.98076, 11.23054, 11.48049, 11.73062, 11.98091, 12.23135, 12.48195, 
    12.73268, 12.98356, 13.23457, 13.4857, 13.73695, 13.98831, 14.23978, 
    14.49135, 14.743, 14.99475, 15.24657, 15.49847, 15.75043, 16.00245, 
    16.25452, 16.50664, 16.7588, 17.01099, 17.26321, 17.51545, 17.76769, 
    18.01995, 18.27221, 18.52446, 18.77669, 19.0289, 19.28109, 19.53324, 
    19.78536, 20.03742, 20.28943, 20.54138, 20.79327, 21.04508, 21.29681, 
    21.54845, 21.8, 22.05146, 22.3028, 22.55403, 22.80515, 23.05613, 
    23.30699, 23.5577, 23.80828, 24.0587, 24.30896, 24.55906, 24.80899, 
    25.05874, 25.30831, 25.55769, 25.80687, 26.05586, 26.30463, 26.5532, 
    26.80154, 27.04966, 27.29755, 27.5452, 27.79261, 28.03977, 28.28667, 
    28.53332, 28.7797, 29.02581, 29.27164, 29.51719, 29.76244, 30.00741, 
    30.25208, 30.49644, 30.74049, 30.98423, 31.22765, 31.47074, 31.71351, 
    31.95593, 32.19802, 32.43976, 32.68115, 32.92219, 33.16287, 33.40318, 
    33.64312, 33.88269, 34.12188, 34.36069, 34.59911, 34.83714, 35.07478, 
    35.31201, 35.54884, 35.78526, 36.02126, 36.25686, 36.49203, 36.72677, 
    36.96109, 37.19497, 37.42842, 37.66143, 37.894, 38.12612, 38.35779, 
    38.58901, 38.81977, 39.05007, 39.2799, 39.50927, 39.73817, 39.9666, 
    40.19455, 40.42203, 40.64902, 40.87553, 41.10154, 41.32708, 41.55211, 
    41.77665, 42.0007, 42.22424, 42.44729, 42.66983, 42.89186, 43.11338, 
    43.33439, 43.55489, 43.77487, 43.99433, 44.21328, 44.4317, 44.6496, 
    44.86697, 45.08382, 45.30014, 45.51593, 45.73119, 45.94592, 46.16011, 
    46.37376, 46.58688, 46.79946, 47.0115, 47.223, 47.43396, 47.64437, 
    47.85424, 48.06357, 48.27235, 48.48058, 48.68827, 48.8954, 49.10199, 
    49.30803, 49.51352, 49.71846, 49.92284, 50.12667, 50.32996, 50.53268, 
    50.73486, 50.93648, 51.13754, 51.33805, 51.53801, 51.73742, 51.93626, 
    52.13456, 52.3323, 52.52948, 52.72611, 52.92219, 53.11771, 53.31267, 
    53.50708, 53.70094, 53.89425, 54.08699, 54.27919, 54.47084, 54.66193, 
    54.85247, 55.04245, 55.23189, 55.42078, 55.60911, 55.7969, 55.98414, 
    56.17083, 56.35697, 56.54256, 56.72761,
  -35.81484, -35.67486, -35.53446, -35.39364, -35.25241, -35.11076, 
    -34.96869, -34.8262, -34.68328, -34.53994, -34.39617, -34.25197, 
    -34.10733, -33.96227, -33.81677, -33.67084, -33.52446, -33.37765, 
    -33.2304, -33.0827, -32.93456, -32.78597, -32.63693, -32.48745, 
    -32.33751, -32.18711, -32.03627, -31.88496, -31.7332, -31.58097, 
    -31.42829, -31.27514, -31.12152, -30.96744, -30.81289, -30.65787, 
    -30.50237, -30.34641, -30.18996, -30.03304, -29.87564, -29.71776, 
    -29.5594, -29.40055, -29.24122, -29.0814, -28.9211, -28.7603, -28.59901, 
    -28.43723, -28.27495, -28.11218, -27.94891, -27.78514, -27.62087, 
    -27.45609, -27.29082, -27.12503, -26.95874, -26.79194, -26.62463, 
    -26.45681, -26.28848, -26.11963, -25.95027, -25.78039, -25.60999, 
    -25.43907, -25.26763, -25.09566, -24.92318, -24.75017, -24.57663, 
    -24.40257, -24.22797, -24.05285, -23.87719, -23.701, -23.52428, 
    -23.34702, -23.16923, -22.9909, -22.81203, -22.63263, -22.45268, 
    -22.27219, -22.09116, -21.90958, -21.72746, -21.5448, -21.36159, 
    -21.17783, -20.99353, -20.80868, -20.62327, -20.43732, -20.25082, 
    -20.06376, -19.87615, -19.68799, -19.49928, -19.31001, -19.12018, 
    -18.92981, -18.73887, -18.54738, -18.35533, -18.16273, -17.96956, 
    -17.77584, -17.58156, -17.38673, -17.19133, -16.99537, -16.79886, 
    -16.60179, -16.40416, -16.20596, -16.00721, -15.8079, -15.60803, 
    -15.4076, -15.20661, -15.00507, -14.80296, -14.6003, -14.39707, -14.1933, 
    -13.98896, -13.78406, -13.57861, -13.37261, -13.16605, -12.95893, 
    -12.75126, -12.54304, -12.33427, -12.12494, -11.91506, -11.70464, 
    -11.49366, -11.28214, -11.07007, -10.85745, -10.64429, -10.43059, 
    -10.21634, -10.00156, -9.786232, -9.57037, -9.353971, -9.137037, 
    -8.919571, -8.701573, -8.483046, -8.263989, -8.044408, -7.824302, 
    -7.603674, -7.382525, -7.160859, -6.938676, -6.715979, -6.492771, 
    -6.269053, -6.044827, -5.820098, -5.594866, -5.369135, -5.142907, 
    -4.916183, -4.688969, -4.461266, -4.233076, -4.004403, -3.77525, 
    -3.54562, -3.315516, -3.08494, -2.853897, -2.62239, -2.390421, -2.157994, 
    -1.925113, -1.691781, -1.458002, -1.223779, -0.9891162, -0.7540172, 
    -0.5184858, -0.2825259, -0.04614144, 0.1906636, 0.4278851, 0.6655189, 
    0.9035611, 1.142007, 1.380853, 1.620094, 1.859725, 2.099744, 2.340144, 
    2.580921, 2.822071, 3.063589, 3.30547, 3.547709, 3.790301, 4.033242, 
    4.276526, 4.52015, 4.764106, 5.00839, 5.252997, 5.497922, 5.74316, 
    5.988704, 6.23455, 6.480692, 6.727125, 6.973843, 7.22084, 7.468111, 
    7.71565, 7.963451, 8.21151, 8.459818, 8.708372, 8.957164, 9.206189, 
    9.455441, 9.704915, 9.954603, 10.2045, 10.4546, 10.7049, 10.95538, 
    11.20605, 11.4569, 11.70792, 11.9591, 12.21044, 12.46194, 12.71357, 
    12.96535, 13.21726, 13.4693, 13.72146, 13.97373, 14.22611, 14.47858, 
    14.73115, 14.98381, 15.23655, 15.48936, 15.74224, 15.99517, 16.24816, 
    16.5012, 16.75428, 17.00739, 17.26052, 17.51368, 17.76685, 18.02002, 
    18.2732, 18.52637, 18.77952, 19.03265, 19.28576, 19.53883, 19.79186, 
    20.04484, 20.29777, 20.55064, 20.80344, 21.05616, 21.3088, 21.56136, 
    21.81382, 22.06618, 22.31844, 22.57057, 22.82259, 23.07448, 23.32624, 
    23.57786, 23.82933, 24.08064, 24.3318, 24.58279, 24.83361, 25.08426, 
    25.33471, 25.58498, 25.83504, 26.08491, 26.33456, 26.584, 26.83322, 
    27.08221, 27.33096, 27.57948, 27.82775, 28.07576, 28.32352, 28.57102, 
    28.81825, 29.0652, 29.31188, 29.55826, 29.80436, 30.05016, 30.29565, 
    30.54084, 30.78572, 31.03027, 31.27451, 31.51841, 31.76198, 32.00521, 
    32.2481, 32.49063, 32.73281, 32.97464, 33.2161, 33.45719, 33.69791, 
    33.93825, 34.17821, 34.41778, 34.65696, 34.89574, 35.13412, 35.3721, 
    35.60967, 35.84682, 36.08356, 36.31988, 36.55577, 36.79123, 37.02626, 
    37.26086, 37.49501, 37.72872, 37.96198, 38.19479, 38.42714, 38.65904, 
    38.89048, 39.12144, 39.35194, 39.58197, 39.81153, 40.04061, 40.2692, 
    40.49732, 40.72495, 40.95208, 41.17873, 41.40488, 41.63053, 41.85568, 
    42.08033, 42.30447, 42.52811, 42.75124, 42.97385, 43.19596, 43.41754, 
    43.63861, 43.85915, 44.07918, 44.29868, 44.51765, 44.73609, 44.95401, 
    45.17139, 45.38824, 45.60455, 45.82033, 46.03557, 46.25027, 46.46443, 
    46.67805, 46.89112, 47.10365, 47.31563, 47.52707, 47.73796, 47.9483, 
    48.15809, 48.36733, 48.57602, 48.78415, 48.99173, 49.19876, 49.40523, 
    49.61115, 49.81651, 50.02132, 50.22557, 50.42926, 50.63239, 50.83497, 
    51.03698, 51.23845, 51.43934, 51.63968, 51.83947, 52.03869, 52.23735, 
    52.43546, 52.633, 52.82998, 53.02641, 53.22227, 53.41758, 53.61233, 
    53.80652, 54.00016, 54.19323, 54.38575, 54.57771, 54.76911, 54.95996, 
    55.15025, 55.33998, 55.52917, 55.71779, 55.90586, 56.09339, 56.28035, 
    56.46677, 56.65264, 56.83795,
  -35.93693, -35.79693, -35.65652, -35.51569, -35.37444, -35.23277, 
    -35.09068, -34.94816, -34.80522, -34.66185, -34.51805, -34.37382, 
    -34.22915, -34.08406, -33.93852, -33.79255, -33.64614, -33.49928, 
    -33.35199, -33.20424, -33.05605, -32.90741, -32.75832, -32.60878, 
    -32.45879, -32.30834, -32.15743, -32.00606, -31.85423, -31.70194, 
    -31.54919, -31.39597, -31.24228, -31.08812, -30.93349, -30.77839, 
    -30.62281, -30.46676, -30.31023, -30.15322, -29.99573, -29.83775, 
    -29.67929, -29.52035, -29.36091, -29.20099, -29.04058, -28.87967, 
    -28.71827, -28.55637, -28.39397, -28.23108, -28.06768, -27.90379, 
    -27.73939, -27.57448, -27.40907, -27.24314, -27.07671, -26.90977, 
    -26.74231, -26.57434, -26.40585, -26.23685, -26.06732, -25.89728, 
    -25.72672, -25.55563, -25.38401, -25.21188, -25.03921, -24.86602, 
    -24.69229, -24.51804, -24.34325, -24.16793, -23.99208, -23.81569, 
    -23.63876, -23.46129, -23.28328, -23.10474, -22.92565, -22.74602, 
    -22.56584, -22.38512, -22.20385, -22.02204, -21.83968, -21.65676, 
    -21.4733, -21.28929, -21.10473, -20.91961, -20.73394, -20.54772, 
    -20.36094, -20.17361, -19.98572, -19.79727, -19.60826, -19.4187, 
    -19.22858, -19.03789, -18.84665, -18.65485, -18.46248, -18.26956, 
    -18.07607, -17.88202, -17.68741, -17.49223, -17.29649, -17.10019, 
    -16.90332, -16.70589, -16.5079, -16.30934, -16.11022, -15.91054, 
    -15.71029, -15.50947, -15.3081, -15.10616, -14.90365, -14.70059, 
    -14.49696, -14.29276, -14.08801, -13.8827, -13.67682, -13.47038, 
    -13.26338, -13.05583, -12.84771, -12.63904, -12.42981, -12.22002, 
    -12.00968, -11.79878, -11.58733, -11.37532, -11.16277, -10.94966, 
    -10.736, -10.5218, -10.30705, -10.09175, -9.875908, -9.659524, -9.442598, 
    -9.225133, -9.00713, -8.788589, -8.569514, -8.349907, -8.129767, 
    -7.909099, -7.687903, -7.466182, -7.243937, -7.021171, -6.797886, 
    -6.574084, -6.349768, -6.124939, -5.899601, -5.673756, -5.447405, 
    -5.220553, -4.993201, -4.765352, -4.53701, -4.308176, -4.078854, 
    -3.849047, -3.618757, -3.387989, -3.156744, -2.925027, -2.69284, 
    -2.460187, -2.227072, -1.993497, -1.759466, -1.524984, -1.290053, 
    -1.054677, -0.8188599, -0.582606, -0.3459189, -0.1088025, 0.128739, 
    0.3667016, 0.6050811, 0.8438734, 1.083074, 1.322679, 1.562683, 1.803083, 
    2.043874, 2.28505, 2.526609, 2.768544, 3.010851, 3.253525, 3.496562, 
    3.739956, 3.983702, 4.227796, 4.472233, 4.717006, 4.962111, 5.207543, 
    5.453297, 5.699367, 5.945746, 6.192432, 6.439417, 6.686696, 6.934263, 
    7.182113, 7.43024, 7.678638, 7.927301, 8.176225, 8.425402, 8.674827, 
    8.924493, 9.174395, 9.424527, 9.674882, 9.925455, 10.17624, 10.42723, 
    10.67842, 10.9298, 11.18136, 11.43311, 11.68503, 11.93711, 12.18936, 
    12.44176, 12.69431, 12.947, 13.19982, 13.45277, 13.70584, 13.95903, 
    14.21232, 14.46572, 14.71921, 14.97278, 15.22644, 15.48018, 15.73398, 
    15.98784, 16.24175, 16.49571, 16.74972, 17.00375, 17.25782, 17.5119, 
    17.766, 18.0201, 18.2742, 18.52829, 18.78237, 19.03643, 19.29046, 
    19.54446, 19.79842, 20.05232, 20.30618, 20.55997, 20.81369, 21.06733, 
    21.3209, 21.57437, 21.82775, 22.08103, 22.3342, 22.58725, 22.84018, 
    23.09299, 23.34565, 23.59818, 23.85055, 24.10277, 24.35483, 24.60673, 
    24.85844, 25.10998, 25.36133, 25.61249, 25.86345, 26.11419, 26.36473, 
    26.61506, 26.86515, 27.11502, 27.36465, 27.61403, 27.86317, 28.11205, 
    28.36067, 28.60903, 28.85711, 29.10492, 29.35244, 29.59967, 29.84661, 
    30.09325, 30.33958, 30.5856, 30.8313, 31.07668, 31.32174, 31.56646, 
    31.81084, 32.05488, 32.29857, 32.54191, 32.78489, 33.0275, 33.26975, 
    33.51163, 33.75312, 33.99424, 34.23497, 34.47531, 34.71525, 34.95479, 
    35.19393, 35.43266, 35.67097, 35.90886, 36.14634, 36.38339, 36.62001, 
    36.85619, 37.09194, 37.32724, 37.5621, 37.79652, 38.03048, 38.26398, 
    38.49702, 38.7296, 38.96171, 39.19336, 39.42452, 39.65522, 39.88543, 
    40.11516, 40.34441, 40.57316, 40.80143, 41.0292, 41.25647, 41.48324, 
    41.70951, 41.93528, 42.16054, 42.38528, 42.60952, 42.83324, 43.05644, 
    43.27913, 43.50129, 43.72293, 43.94404, 44.16462, 44.38468, 44.6042, 
    44.82319, 45.04165, 45.25957, 45.47695, 45.69379, 45.91009, 46.12584, 
    46.34105, 46.55572, 46.76984, 46.98341, 47.19643, 47.40889, 47.62081, 
    47.83218, 48.04298, 48.25324, 48.46294, 48.67208, 48.88067, 49.0887, 
    49.29617, 49.50307, 49.70942, 49.91521, 50.12044, 50.3251, 50.52921, 
    50.73275, 50.93572, 51.13814, 51.33999, 51.54128, 51.742, 51.94216, 
    52.14176, 52.34079, 52.53926, 52.73716, 52.9345, 53.13128, 53.32749, 
    53.52314, 53.71823, 53.91275, 54.10671, 54.30011, 54.49295, 54.68523, 
    54.87694, 55.06809, 55.25869, 55.44872, 55.6382, 55.82711, 56.01548, 
    56.20328, 56.39053, 56.57721, 56.76335, 56.94893,
  -36.05952, -35.91951, -35.77909, -35.63824, -35.49697, -35.35529, 
    -35.21317, -35.07064, -34.92767, -34.78428, -34.64045, -34.49619, 
    -34.3515, -34.20637, -34.0608, -33.91479, -33.76834, -33.62144, 
    -33.47411, -33.32632, -33.17809, -33.0294, -32.88026, -32.73067, 
    -32.58062, -32.43011, -32.27914, -32.12772, -31.97583, -31.82347, 
    -31.67065, -31.51736, -31.3636, -31.20937, -31.05466, -30.89948, 
    -30.74382, -30.58769, -30.43107, -30.27397, -30.11639, -29.95832, 
    -29.79976, -29.64072, -29.48119, -29.32116, -29.16064, -28.99962, 
    -28.83811, -28.6761, -28.51359, -28.35057, -28.18706, -28.02303, 
    -27.8585, -27.69346, -27.52792, -27.36186, -27.19529, -27.0282, -26.8606, 
    -26.69247, -26.52384, -26.35468, -26.18499, -26.01479, -25.84406, 
    -25.6728, -25.50102, -25.32871, -25.15586, -24.98249, -24.80858, 
    -24.63414, -24.45916, -24.28365, -24.10759, -23.931, -23.75386, 
    -23.57619, -23.39797, -23.21921, -23.0399, -22.86004, -22.67964, 
    -22.49869, -22.31719, -22.13513, -21.95253, -21.76937, -21.58566, 
    -21.4014, -21.21658, -21.0312, -20.84526, -20.65877, -20.47172, -20.2841, 
    -20.09593, -19.9072, -19.7179, -19.52804, -19.33762, -19.14663, 
    -18.95508, -18.76297, -18.57029, -18.37704, -18.18323, -17.98885, 
    -17.7939, -17.59839, -17.40231, -17.20566, -17.00844, -16.81065, 
    -16.6123, -16.41338, -16.21388, -16.01382, -15.8132, -15.612, -15.41023, 
    -15.2079, -15.005, -14.80153, -14.59749, -14.39288, -14.18771, -13.98197, 
    -13.77567, -13.5688, -13.36136, -13.15337, -12.9448, -12.73568, 
    -12.52599, -12.31574, -12.10493, -11.89356, -11.68163, -11.46914, 
    -11.2561, -11.0425, -10.82834, -10.61364, -10.39838, -10.18257, 
    -9.966207, -9.749299, -9.531845, -9.313846, -9.095304, -8.87622, 
    -8.656595, -8.436433, -8.215734, -7.994501, -7.772735, -7.550438, 
    -7.327612, -7.104261, -6.880385, -6.655987, -6.43107, -6.205635, 
    -5.979685, -5.753222, -5.52625, -5.298771, -5.070787, -4.842301, 
    -4.613316, -4.383834, -4.15386, -3.923394, -3.692442, -3.461005, 
    -3.229088, -2.996693, -2.763823, -2.530482, -2.296674, -2.062401, 
    -1.827667, -1.592477, -1.356833, -1.12074, -0.884201, -0.6472201, 
    -0.4098012, -0.1719483, 0.0663344, 0.3050429, 0.544173, 0.7837204, 
    1.023681, 1.26405, 1.504823, 1.745996, 1.987564, 2.229523, 2.471867, 
    2.714593, 2.957695, 3.201168, 3.445008, 3.689209, 3.933767, 4.178677, 
    4.423932, 4.669529, 4.915462, 5.161724, 5.408312, 5.65522, 5.902442, 
    6.149973, 6.397807, 6.645938, 6.894361, 7.143071, 7.39206, 7.641324, 
    7.890857, 8.140652, 8.390704, 8.641006, 8.891554, 9.14234, 9.393358, 
    9.644603, 9.896067, 10.14775, 10.39963, 10.65172, 10.904, 11.15647, 
    11.40912, 11.66195, 11.91494, 12.1681, 12.42142, 12.67488, 12.92849, 
    13.18223, 13.4361, 13.69009, 13.9442, 14.19842, 14.45274, 14.70716, 
    14.96167, 15.21625, 15.47092, 15.72565, 15.98044, 16.23529, 16.49018, 
    16.74512, 17.00009, 17.25509, 17.5101, 17.76513, 18.02017, 18.27521, 
    18.53024, 18.78525, 19.04025, 19.29521, 19.55014, 19.80503, 20.05987, 
    20.31465, 20.56937, 20.82402, 21.0786, 21.33309, 21.58749, 21.8418, 
    22.096, 22.35009, 22.60407, 22.85792, 23.11164, 23.36522, 23.61866, 
    23.87195, 24.12509, 24.37806, 24.63086, 24.88348, 25.13592, 25.38817, 
    25.64023, 25.89208, 26.14372, 26.39515, 26.64636, 26.89735, 27.14809, 
    27.3986, 27.64887, 27.89888, 28.14863, 28.39812, 28.64734, 28.89629, 
    29.14495, 29.39333, 29.64142, 29.8892, 30.13668, 30.38386, 30.63071, 
    30.87725, 31.12346, 31.36934, 31.61489, 31.86009, 32.10494, 32.34944, 
    32.59359, 32.83737, 33.08078, 33.32383, 33.56649, 33.80878, 34.05067, 
    34.29218, 34.53329, 34.774, 35.01431, 35.2542, 35.49368, 35.73275, 
    35.97139, 36.2096, 36.44739, 36.68473, 36.92165, 37.15812, 37.39414, 
    37.62971, 37.86483, 38.09949, 38.33369, 38.56742, 38.80069, 39.03349, 
    39.2658, 39.49765, 39.72901, 39.95988, 40.19027, 40.42017, 40.64957, 
    40.87848, 41.10688, 41.33479, 41.56219, 41.78908, 42.01546, 42.24133, 
    42.46668, 42.69152, 42.91583, 43.13963, 43.3629, 43.58564, 43.80785, 
    44.02953, 44.25068, 44.47129, 44.69137, 44.91091, 45.12991, 45.34837, 
    45.56628, 45.78365, 46.00047, 46.21674, 46.43246, 46.64764, 46.86226, 
    47.07632, 47.28983, 47.50279, 47.71519, 47.92703, 48.13831, 48.34903, 
    48.55919, 48.7688, 48.97783, 49.18631, 49.39421, 49.60156, 49.80834, 
    50.01456, 50.2202, 50.42529, 50.6298, 50.83375, 51.03713, 51.23994, 
    51.44218, 51.64386, 51.84497, 52.04551, 52.24548, 52.44488, 52.64371, 
    52.84198, 53.03967, 53.2368, 53.43336, 53.62935, 53.82478, 54.01963, 
    54.21392, 54.40765, 54.6008, 54.7934, 54.98542, 55.17688, 55.36778, 
    55.55811, 55.74788, 55.93709, 56.12573, 56.31382, 56.50134, 56.6883, 
    56.87471, 57.06056,
  -36.18262, -36.0426, -35.90216, -35.7613, -35.62002, -35.47832, -35.33619, 
    -35.19363, -35.05064, -34.90723, -34.76337, -34.61909, -34.47437, 
    -34.3292, -34.18361, -34.03756, -33.89108, -33.74414, -33.59676, 
    -33.44894, -33.30066, -33.15192, -33.00274, -32.8531, -32.703, -32.55243, 
    -32.40141, -32.24993, -32.09797, -31.94556, -31.79267, -31.63931, 
    -31.48548, -31.33118, -31.1764, -31.02114, -30.8654, -30.70918, 
    -30.55248, -30.3953, -30.23763, -30.07947, -29.92082, -29.76168, 
    -29.60205, -29.44192, -29.28129, -29.12017, -28.95855, -28.79642, 
    -28.63379, -28.47066, -28.30702, -28.14288, -27.97822, -27.81305, 
    -27.64737, -27.48118, -27.31447, -27.14724, -26.97949, -26.81122, 
    -26.64244, -26.47312, -26.30328, -26.13292, -25.96202, -25.7906, 
    -25.61865, -25.44616, -25.27314, -25.09959, -24.9255, -24.75087, 
    -24.5757, -24.39999, -24.22374, -24.04695, -23.86961, -23.69172, 
    -23.51329, -23.33432, -23.15479, -22.97471, -22.79408, -22.6129, 
    -22.43117, -22.24888, -22.06603, -21.88263, -21.69867, -21.51415, 
    -21.32907, -21.14343, -20.95723, -20.77047, -20.58314, -20.39525, 
    -20.2068, -20.01778, -19.82819, -19.63804, -19.44732, -19.25603, 
    -19.06417, -18.87175, -18.67875, -18.48518, -18.29105, -18.09634, 
    -17.90106, -17.7052, -17.50878, -17.31178, -17.11421, -16.91607, 
    -16.71736, -16.51807, -16.31821, -16.11777, -15.91676, -15.71518, 
    -15.51303, -15.3103, -15.107, -14.90312, -14.69868, -14.49366, -14.28807, 
    -14.08191, -13.87517, -13.66787, -13.46, -13.25155, -13.04254, -12.83296, 
    -12.62282, -12.4121, -12.20082, -11.98898, -11.77657, -11.5636, 
    -11.35007, -11.13598, -10.92132, -10.70611, -10.49034, -10.27402, 
    -10.05714, -9.839704, -9.621718, -9.403184, -9.1841, -8.96447, -8.744294, 
    -8.523575, -8.302314, -8.080513, -7.858175, -7.635301, -7.411892, 
    -7.187953, -6.963483, -6.738486, -6.512965, -6.286921, -6.060356, 
    -5.833274, -5.605677, -5.377567, -5.148947, -4.91982, -4.690189, 
    -4.460057, -4.229426, -3.9983, -3.766681, -3.534572, -3.301978, 
    -3.068901, -2.835344, -2.601311, -2.366806, -2.131831, -1.896391, 
    -1.660488, -1.424128, -1.187312, -0.9500467, -0.7123342, -0.4741789, 
    -0.2355848, 0.003443994, 0.2429032, 0.4827888, 0.7230963, 0.9638215, 
    1.20496, 1.446507, 1.688458, 1.930809, 2.173555, 2.416692, 2.660213, 
    2.904116, 3.148394, 3.393042, 3.638057, 3.883432, 4.129162, 4.375243, 
    4.621669, 4.868435, 5.115535, 5.362964, 5.610716, 5.858787, 6.107169, 
    6.355859, 6.604849, 6.854135, 7.10371, 7.353569, 7.603705, 7.854113, 
    8.104787, 8.355721, 8.606909, 8.858344, 9.110021, 9.361932, 9.614073, 
    9.866436, 10.11902, 10.37181, 10.6248, 10.87799, 11.13137, 11.38493, 
    11.63868, 11.89259, 12.14667, 12.4009, 12.65529, 12.90982, 13.16449, 
    13.41929, 13.67421, 13.92925, 14.18441, 14.43966, 14.69501, 14.95045, 
    15.20598, 15.46158, 15.71725, 15.97298, 16.22877, 16.48461, 16.74048, 
    16.9964, 17.25233, 17.50829, 17.76427, 18.02025, 18.27622, 18.5322, 
    18.78815, 19.04409, 19.3, 19.55587, 19.8117, 20.06747, 20.3232, 20.57886, 
    20.83445, 21.08996, 21.34539, 21.60072, 21.85596, 22.1111, 22.36612, 
    22.62102, 22.8758, 23.13045, 23.38496, 23.63932, 23.89353, 24.14758, 
    24.40147, 24.65519, 24.90872, 25.16208, 25.41523, 25.6682, 25.92095, 
    26.1735, 26.42583, 26.67793, 26.92981, 27.18145, 27.43284, 27.68399, 
    27.93488, 28.18551, 28.43588, 28.68597, 28.93579, 29.18532, 29.43456, 
    29.6835, 29.93214, 30.18048, 30.4285, 30.6762, 30.92357, 31.17062, 
    31.41733, 31.66371, 31.90973, 32.15541, 32.40073, 32.64568, 32.89027, 
    33.13449, 33.37833, 33.6218, 33.86487, 34.10755, 34.34984, 34.59173, 
    34.83321, 35.07428, 35.31495, 35.55518, 35.795, 36.03439, 36.27335, 
    36.51188, 36.74997, 36.98761, 37.2248, 37.46155, 37.69783, 37.93366, 
    38.16903, 38.40393, 38.63836, 38.87232, 39.1058, 39.3388, 39.57132, 
    39.80335, 40.03489, 40.26594, 40.49649, 40.72655, 40.9561, 41.18515, 
    41.41368, 41.64171, 41.86923, 42.09623, 42.32271, 42.54867, 42.77411, 
    42.99903, 43.22341, 43.44727, 43.67059, 43.89338, 44.11563, 44.33735, 
    44.55853, 44.77916, 44.99925, 45.21879, 45.43779, 45.65624, 45.87413, 
    46.09148, 46.30827, 46.52451, 46.74019, 46.95531, 47.16988, 47.38388, 
    47.59733, 47.81021, 48.02253, 48.23428, 48.44547, 48.6561, 48.86615, 
    49.07564, 49.28456, 49.49292, 49.7007, 49.90791, 50.11456, 50.32063, 
    50.52613, 50.73106, 50.93541, 51.13919, 51.3424, 51.54504, 51.7471, 
    51.9486, 52.14951, 52.34986, 52.54963, 52.74883, 52.94745, 53.1455, 
    53.34298, 53.53989, 53.73623, 53.93198, 54.12717, 54.32179, 54.51584, 
    54.70932, 54.90222, 55.09456, 55.28633, 55.47752, 55.66816, 55.85822, 
    56.04771, 56.23664, 56.42501, 56.61281, 56.80005, 56.98672, 57.17283,
  -36.30622, -36.16619, -36.02575, -35.88488, -35.74358, -35.60186, 
    -35.45972, -35.31714, -35.17414, -35.0307, -34.88683, -34.74252, 
    -34.59777, -34.45258, -34.30695, -34.16087, -34.01435, -33.86738, 
    -33.71997, -33.5721, -33.42378, -33.275, -33.12577, -32.97608, -32.82593, 
    -32.67531, -32.52423, -32.37269, -32.22068, -32.0682, -31.91525, 
    -31.76183, -31.60793, -31.45356, -31.29871, -31.14337, -30.98756, 
    -30.83126, -30.67448, -30.51721, -30.35945, -30.2012, -30.04246, 
    -29.88322, -29.72349, -29.56326, -29.40254, -29.24131, -29.07958, 
    -28.91734, -28.7546, -28.59135, -28.4276, -28.26333, -28.09855, 
    -27.93325, -27.76744, -27.60111, -27.43426, -27.2669, -27.099, -26.93059, 
    -26.76165, -26.59219, -26.42219, -26.25167, -26.08061, -25.90903, 
    -25.7369, -25.56425, -25.39105, -25.21732, -25.04305, -24.86823, 
    -24.69287, -24.51697, -24.34053, -24.16353, -23.98599, -23.8079, 
    -23.62926, -23.45007, -23.27033, -23.09003, -22.90917, -22.72776, 
    -22.5458, -22.36327, -22.18018, -21.99654, -21.81233, -21.62756, 
    -21.44222, -21.25632, -21.06986, -20.88283, -20.69523, -20.50706, 
    -20.31833, -20.12902, -19.93915, -19.7487, -19.55768, -19.36609, 
    -19.17393, -18.98119, -18.78788, -18.59399, -18.39953, -18.20449, 
    -18.00888, -17.81269, -17.61592, -17.41858, -17.22066, -17.02216, 
    -16.82308, -16.62343, -16.42319, -16.22238, -16.02099, -15.81903, 
    -15.61648, -15.41336, -15.20966, -15.00538, -14.80053, -14.59509, 
    -14.38908, -14.1825, -13.97534, -13.7676, -13.55929, -13.3504, -13.14094, 
    -12.93091, -12.7203, -12.50912, -12.29737, -12.08506, -11.87217, 
    -11.65871, -11.44469, -11.2301, -11.01494, -10.79923, -10.58295, 
    -10.3661, -10.1487, -9.930742, -9.712226, -9.493153, -9.273526, 
    -9.053348, -8.832619, -8.611341, -8.389515, -8.167145, -7.944231, 
    -7.720777, -7.496783, -7.272252, -7.047186, -6.821588, -6.595459, 
    -6.368803, -6.141621, -5.913916, -5.68569, -5.456947, -5.227689, 
    -4.997918, -4.767638, -4.536851, -4.30556, -4.073769, -3.84148, 
    -3.608696, -3.375421, -3.141658, -2.907411, -2.672682, -2.437475, 
    -2.201794, -1.965642, -1.729024, -1.491942, -1.2544, -1.016403, 
    -0.7779544, -0.5390579, -0.2997179, -0.05993829, 0.1802766, 0.4209225, 
    0.6619952, 0.9034902, 1.145403, 1.38773, 1.630465, 1.873604, 2.117143, 
    2.361076, 2.6054, 2.850108, 3.095196, 3.34066, 3.586493, 3.832691, 
    4.079249, 4.326161, 4.573422, 4.821027, 5.068971, 5.317247, 5.56585, 
    5.814775, 6.064016, 6.313568, 6.563424, 6.813578, 7.064026, 7.314761, 
    7.565776, 7.817067, 8.068626, 8.32045, 8.572529, 8.824859, 9.077434, 
    9.330246, 9.58329, 9.836559, 10.09005, 10.34375, 10.59766, 10.85176, 
    11.10606, 11.36055, 11.61521, 11.87005, 12.12506, 12.38022, 12.63554, 
    12.891, 13.1466, 13.40234, 13.6582, 13.91418, 14.17027, 14.42647, 
    14.68276, 14.93915, 15.19562, 15.45216, 15.70878, 15.96546, 16.2222, 
    16.47898, 16.73581, 16.99267, 17.24956, 17.50647, 17.76339, 18.02032, 
    18.27725, 18.53417, 18.79108, 19.04796, 19.30482, 19.56164, 19.81842, 
    20.07515, 20.33182, 20.58842, 20.84496, 21.10141, 21.35778, 21.61407, 
    21.87024, 22.12632, 22.38228, 22.63812, 22.89384, 23.14942, 23.40486, 
    23.66015, 23.91529, 24.17027, 24.42508, 24.67972, 24.93418, 25.18845, 
    25.44252, 25.6964, 25.95006, 26.20352, 26.45675, 26.70976, 26.96254, 
    27.21507, 27.46736, 27.7194, 27.97118, 28.2227, 28.47395, 28.72492, 
    28.97561, 29.22601, 29.47612, 29.72593, 29.97543, 30.22462, 30.4735, 
    30.72205, 30.97027, 31.21816, 31.46571, 31.71292, 31.95978, 32.20628, 
    32.45242, 32.69819, 32.9436, 33.18863, 33.43327, 33.67754, 33.92141, 
    34.16488, 34.40796, 34.65063, 34.89289, 35.13474, 35.37617, 35.61717, 
    35.85775, 36.0979, 36.33761, 36.57688, 36.8157, 37.05408, 37.29201, 
    37.52948, 37.76648, 38.00303, 38.23911, 38.47471, 38.70984, 38.9445, 
    39.17867, 39.41235, 39.64555, 39.87826, 40.11047, 40.34218, 40.57339, 
    40.8041, 41.0343, 41.26399, 41.49316, 41.72182, 41.94997, 42.17759, 
    42.40469, 42.63126, 42.85731, 43.08282, 43.3078, 43.53225, 43.75616, 
    43.97953, 44.20235, 44.42464, 44.64638, 44.86757, 45.08821, 45.3083, 
    45.52784, 45.74683, 45.96526, 46.18313, 46.40044, 46.6172, 46.83339, 
    47.04902, 47.26408, 47.47858, 47.69251, 47.90588, 48.11868, 48.33091, 
    48.54256, 48.75365, 48.96417, 49.17411, 49.38348, 49.59228, 49.8005, 
    50.00814, 50.21521, 50.42171, 50.62763, 50.83297, 51.03773, 51.24192, 
    51.44553, 51.64856, 51.85101, 52.05289, 52.25418, 52.45491, 52.65504, 
    52.85461, 53.05359, 53.252, 53.44983, 53.64708, 53.84376, 54.03986, 
    54.23538, 54.43033, 54.6247, 54.81849, 55.01171, 55.20436, 55.39643, 
    55.58794, 55.77886, 55.96922, 56.159, 56.34822, 56.53687, 56.72494, 
    56.91245, 57.09939, 57.28577,
  -36.43033, -36.2903, -36.14985, -36.00897, -35.86766, -35.72593, -35.58377, 
    -35.44118, -35.29816, -35.1547, -35.01081, -34.86647, -34.7217, 
    -34.57648, -34.43082, -34.28472, -34.13817, -33.99117, -33.84371, 
    -33.69581, -33.54745, -33.39863, -33.24935, -33.09961, -32.94941, 
    -32.79875, -32.64762, -32.49603, -32.34396, -32.19142, -32.03841, 
    -31.88492, -31.73096, -31.57651, -31.42159, -31.26618, -31.11029, 
    -30.95392, -30.79706, -30.6397, -30.48186, -30.32352, -30.16469, 
    -30.00536, -29.84554, -29.68521, -29.52438, -29.36305, -29.20121, 
    -29.03887, -28.87601, -28.71265, -28.54877, -28.38439, -28.21948, 
    -28.05406, -27.88812, -27.72166, -27.55468, -27.38717, -27.21914, 
    -27.05058, -26.88149, -26.71188, -26.54173, -26.37105, -26.19983, 
    -26.02808, -25.85579, -25.68297, -25.5096, -25.33569, -25.16123, 
    -24.98624, -24.81069, -24.6346, -24.45796, -24.28077, -24.10303, 
    -23.92473, -23.74588, -23.56648, -23.38652, -23.206, -23.02492, 
    -22.84328, -22.66108, -22.47832, -22.29499, -22.1111, -21.92665, 
    -21.74162, -21.55604, -21.36988, -21.18315, -20.99585, -20.80798, 
    -20.61954, -20.43052, -20.24093, -20.05077, -19.86003, -19.66871, 
    -19.47682, -19.28435, -19.0913, -18.89767, -18.70347, -18.50868, 
    -18.31331, -18.11737, -17.92084, -17.72373, -17.52604, -17.32777, 
    -17.12891, -16.92948, -16.72946, -16.52885, -16.32767, -16.1259, 
    -15.92355, -15.72061, -15.51709, -15.31299, -15.10831, -14.90305, 
    -14.6972, -14.49077, -14.28376, -14.07617, -13.868, -13.65924, -13.44991, 
    -13.24, -13.02951, -12.81845, -12.6068, -12.39458, -12.18179, -11.96842, 
    -11.75448, -11.53996, -11.32487, -11.10922, -10.89299, -10.6762, 
    -10.45884, -10.24091, -10.02242, -9.803372, -9.58376, -9.363589, 
    -9.142859, -8.921575, -8.699735, -8.477344, -8.254401, -8.03091, 
    -7.806873, -7.582291, -7.357166, -7.131502, -6.905299, -6.678561, 
    -6.451289, -6.223487, -5.995156, -5.766299, -5.536919, -5.307019, 
    -5.076601, -4.845668, -4.614223, -4.382269, -4.149809, -3.916846, 
    -3.683383, -3.449424, -3.214971, -2.980029, -2.7446, -2.508687, 
    -2.272296, -2.035429, -1.79809, -1.560282, -1.32201, -1.083277, 
    -0.8440869, -0.6044447, -0.3643538, -0.1238185, 0.1171569, 0.3585683, 
    0.6004112, 0.8426812, 1.085374, 1.328485, 1.572009, 1.815942, 2.060279, 
    2.305015, 2.550146, 2.795666, 3.041571, 3.287855, 3.534513, 3.78154, 
    4.028931, 4.27668, 4.524784, 4.773234, 5.022027, 5.271156, 5.520617, 
    5.770403, 6.020509, 6.270929, 6.521657, 6.772688, 7.024014, 7.275632, 
    7.527534, 7.779714, 8.032166, 8.284885, 8.537864, 8.791096, 9.044575, 
    9.298295, 9.55225, 9.806433, 10.06084, 10.31546, 10.57028, 10.82531, 
    11.08054, 11.33595, 11.59155, 11.84732, 12.10326, 12.35936, 12.61562, 
    12.87202, 13.12857, 13.38525, 13.64205, 13.89898, 14.15602, 14.41316, 
    14.67041, 14.92775, 15.18517, 15.44267, 15.70024, 15.95788, 16.21557, 
    16.47331, 16.73109, 16.98891, 17.24676, 17.50463, 17.76251, 18.0204, 
    18.27828, 18.53617, 18.79403, 19.05187, 19.30969, 19.56746, 19.8252, 
    20.08288, 20.34051, 20.59807, 20.85556, 21.11296, 21.37029, 21.62752, 
    21.88465, 22.14167, 22.39858, 22.65536, 22.91202, 23.16855, 23.42493, 
    23.68116, 23.93723, 24.19315, 24.44889, 24.70446, 24.95984, 25.21504, 
    25.47004, 25.72483, 25.97942, 26.23379, 26.48794, 26.74186, 26.99554, 
    27.24898, 27.50217, 27.75511, 28.00779, 28.26019, 28.51233, 28.76419, 
    29.01576, 29.26704, 29.51802, 29.7687, 30.01908, 30.26913, 30.51887, 
    30.76827, 31.01735, 31.26609, 31.51449, 31.76253, 32.01023, 32.25756, 
    32.50453, 32.75113, 32.99735, 33.2432, 33.48866, 33.73372, 33.9784, 
    34.22267, 34.46654, 34.71, 34.95304, 35.19567, 35.43787, 35.67965, 
    35.92099, 36.1619, 36.40236, 36.64238, 36.88195, 37.12107, 37.35973, 
    37.59793, 37.83566, 38.07293, 38.30972, 38.54604, 38.78187, 39.01722, 
    39.25209, 39.48647, 39.72034, 39.95373, 40.18661, 40.41899, 40.65087, 
    40.88223, 41.11308, 41.34342, 41.57324, 41.80254, 42.03131, 42.25956, 
    42.48727, 42.71446, 42.94112, 43.16723, 43.39281, 43.61785, 43.84235, 
    44.0663, 44.2897, 44.51256, 44.73486, 44.95662, 45.17781, 45.39845, 
    45.61854, 45.83806, 46.05702, 46.27542, 46.49326, 46.71053, 46.92723, 
    47.14337, 47.35894, 47.57393, 47.78836, 48.00221, 48.21549, 48.42819, 
    48.64032, 48.85187, 49.06285, 49.27324, 49.48306, 49.6923, 49.90096, 
    50.10904, 50.31654, 50.52346, 50.7298, 50.93555, 51.14073, 51.34532, 
    51.54932, 51.75275, 51.95559, 52.15785, 52.35953, 52.56062, 52.76114, 
    52.96106, 53.16041, 53.35917, 53.55735, 53.75495, 53.95197, 54.1484, 
    54.34426, 54.53953, 54.73423, 54.92834, 55.12188, 55.31483, 55.50721, 
    55.69901, 55.89024, 56.08089, 56.27096, 56.46046, 56.64938, 56.83773, 
    57.02552, 57.21272, 57.39936,
  -36.55496, -36.41492, -36.27446, -36.13358, -35.99227, -35.85052, 
    -35.70835, -35.56575, -35.42271, -35.27924, -35.13532, -34.99097, 
    -34.84617, -34.70093, -34.55524, -34.40911, -34.26253, -34.11549, 
    -33.96801, -33.82006, -33.67167, -33.52281, -33.37349, -33.22371, 
    -33.07346, -32.92275, -32.77157, -32.61992, -32.4678, -32.3152, 
    -32.16213, -32.00858, -31.85456, -31.70004, -31.54505, -31.38958, 
    -31.23361, -31.07716, -30.92022, -30.76279, -30.60486, -30.44644, 
    -30.28752, -30.1281, -29.96818, -29.80775, -29.64683, -29.48539, 
    -29.32345, -29.161, -28.99804, -28.83456, -28.67057, -28.50606, 
    -28.34103, -28.17549, -28.00942, -27.84283, -27.67571, -27.50807, 
    -27.3399, -27.1712, -27.00197, -26.8322, -26.6619, -26.49106, -26.31969, 
    -26.14778, -25.97532, -25.80233, -25.62879, -25.4547, -25.28007, 
    -25.10489, -24.92916, -24.75287, -24.57604, -24.39865, -24.22071, 
    -24.04221, -23.86316, -23.68354, -23.50336, -23.32262, -23.14132, 
    -22.95946, -22.77703, -22.59403, -22.41047, -22.22634, -22.04163, 
    -21.85636, -21.67052, -21.4841, -21.29711, -21.10954, -20.9214, 
    -20.73268, -20.54339, -20.35351, -20.16306, -19.97203, -19.78042, 
    -19.58822, -19.39545, -19.20209, -19.00815, -18.81362, -18.61851, 
    -18.42282, -18.22654, -18.02967, -17.83222, -17.63418, -17.43556, 
    -17.23635, -17.03655, -16.83616, -16.63519, -16.43363, -16.23148, 
    -16.02874, -15.82542, -15.6215, -15.417, -15.21192, -15.00624, -14.79998, 
    -14.59313, -14.38569, -14.17767, -13.96906, -13.75987, -13.55009, 
    -13.33973, -13.12879, -12.91726, -12.70515, -12.49246, -12.27918, 
    -12.06533, -11.8509, -11.63589, -11.42031, -11.20415, -10.98741, 
    -10.77011, -10.55223, -10.33377, -10.11475, -9.895167, -9.675014, 
    -9.454295, -9.233013, -9.011169, -8.788767, -8.565806, -8.34229, 
    -8.118219, -7.893597, -7.668424, -7.442703, -7.216437, -6.989627, 
    -6.762276, -6.534387, -6.305961, -6.077001, -5.847509, -5.61749, 
    -5.386944, -5.155875, -4.924286, -4.69218, -4.459559, -4.226427, 
    -3.992786, -3.75864, -3.523993, -3.288846, -3.053205, -2.817072, 
    -2.58045, -2.343344, -2.105757, -1.867692, -1.629154, -1.390147, 
    -1.150673, -0.9107382, -0.6703454, -0.4294989, -0.188203, 0.05353804, 
    0.2957199, 0.5383382, 0.7813884, 1.024866, 1.268767, 1.513085, 1.757818, 
    2.002959, 2.248503, 2.494447, 2.740785, 2.987511, 3.234622, 3.482111, 
    3.729973, 3.978203, 4.226797, 4.475747, 4.725049, 4.974698, 5.224688, 
    5.475012, 5.725666, 5.976644, 6.227939, 6.479546, 6.731459, 6.983672, 
    7.236179, 7.488974, 7.742051, 7.995403, 8.249024, 8.502909, 8.75705, 
    9.011441, 9.266077, 9.520949, 9.776053, 10.03138, 10.28693, 10.54268, 
    10.79865, 11.0548, 11.31115, 11.56769, 11.8244, 12.08128, 12.33833, 
    12.59553, 12.85288, 13.11038, 13.36801, 13.62577, 13.88365, 14.14164, 
    14.39975, 14.65795, 14.91625, 15.17463, 15.43309, 15.69163, 15.95023, 
    16.20888, 16.46759, 16.72634, 16.98512, 17.24393, 17.50277, 17.76162, 
    18.02047, 18.27933, 18.53817, 18.79701, 19.05581, 19.31459, 19.57334, 
    19.83204, 20.09068, 20.34927, 20.6078, 20.86625, 21.12462, 21.3829, 
    21.64109, 21.89917, 22.15715, 22.41501, 22.67275, 22.93036, 23.18784, 
    23.44517, 23.70234, 23.95936, 24.21622, 24.4729, 24.72941, 24.98573, 
    25.24186, 25.49779, 25.75351, 26.00902, 26.26431, 26.51938, 26.77422, 
    27.02882, 27.28317, 27.53727, 27.79111, 28.04469, 28.298, 28.55103, 
    28.80378, 29.05624, 29.30841, 29.56027, 29.81183, 30.06308, 30.314, 
    30.56461, 30.81488, 31.06482, 31.31441, 31.56366, 31.81255, 32.06109, 
    32.30926, 32.55706, 32.80449, 33.05154, 33.29821, 33.54448, 33.79036, 
    34.03585, 34.28092, 34.52559, 34.76984, 35.01368, 35.25709, 35.50007, 
    35.74262, 35.98473, 36.2264, 36.46763, 36.7084, 36.94872, 37.18858, 
    37.42799, 37.66692, 37.90538, 38.14337, 38.38088, 38.61791, 38.85446, 
    39.09051, 39.32608, 39.56114, 39.79571, 40.02978, 40.26334, 40.49639, 
    40.72893, 40.96095, 41.19246, 41.42345, 41.65391, 41.88385, 42.11325, 
    42.34213, 42.57047, 42.79827, 43.02554, 43.25227, 43.47844, 43.70408, 
    43.92916, 44.1537, 44.37768, 44.60111, 44.82399, 45.0463, 45.26805, 
    45.48925, 45.70988, 45.92994, 46.14944, 46.36837, 46.58673, 46.80452, 
    47.02174, 47.23838, 47.45445, 47.66994, 47.88486, 48.0992, 48.31296, 
    48.52614, 48.73874, 48.95076, 49.16219, 49.37305, 49.58332, 49.793, 
    50.0021, 50.21062, 50.41854, 50.62589, 50.83265, 51.03881, 51.2444, 
    51.44939, 51.6538, 51.85762, 52.06085, 52.2635, 52.46555, 52.66702, 
    52.8679, 53.0682, 53.2679, 53.46702, 53.66555, 53.86349, 54.06085, 
    54.25763, 54.45381, 54.64941, 54.84443, 55.03886, 55.23271, 55.42598, 
    55.61866, 55.81076, 56.00229, 56.19323, 56.38359, 56.57337, 56.76257, 
    56.9512, 57.13925, 57.32673, 57.51363,
  -36.6801, -36.54006, -36.3996, -36.25871, -36.11739, -35.97564, -35.83346, 
    -35.69085, -35.54779, -35.4043, -35.26037, -35.116, -34.97118, -34.82592, 
    -34.68021, -34.53405, -34.38744, -34.24038, -34.09285, -33.94488, 
    -33.79644, -33.64755, -33.49819, -33.34837, -33.19807, -33.04732, 
    -32.89609, -32.74438, -32.59221, -32.43956, -32.28643, -32.13282, 
    -31.97873, -31.82416, -31.6691, -31.51356, -31.35752, -31.20099, 
    -31.04398, -30.88646, -30.72845, -30.56995, -30.41094, -30.25143, 
    -30.09142, -29.9309, -29.76988, -29.60834, -29.4463, -29.28374, 
    -29.12067, -28.95708, -28.79298, -28.62835, -28.46321, -28.29754, 
    -28.13134, -27.96462, -27.79738, -27.6296, -27.46129, -27.29245, 
    -27.12307, -26.95316, -26.78271, -26.61172, -26.44019, -26.26811, 
    -26.09549, -25.92233, -25.74862, -25.57436, -25.39955, -25.22419, 
    -25.04827, -24.8718, -24.69478, -24.51719, -24.33905, -24.16035, 
    -23.98109, -23.80126, -23.62087, -23.43991, -23.25839, -23.0763, 
    -22.89364, -22.71041, -22.52661, -22.34224, -22.15729, -21.97177, 
    -21.78567, -21.599, -21.41174, -21.22391, -21.0355, -20.84651, -20.65693, 
    -20.46678, -20.27604, -20.08471, -19.8928, -19.70031, -19.50723, 
    -19.31356, -19.1193, -18.92446, -18.72903, -18.533, -18.33639, -18.13919, 
    -17.9414, -17.74301, -17.54404, -17.34447, -17.14431, -16.94356, 
    -16.74221, -16.54028, -16.33775, -16.13462, -15.93091, -15.7266, 
    -15.5217, -15.31621, -15.11012, -14.90344, -14.69617, -14.48831, 
    -14.27986, -14.07081, -13.86118, -13.65095, -13.44014, -13.22874, 
    -13.01675, -12.80417, -12.591, -12.37725, -12.16292, -11.948, -11.7325, 
    -11.51641, -11.29974, -11.0825, -10.86467, -10.64627, -10.42729, 
    -10.20774, -9.987617, -9.766919, -9.545651, -9.323814, -9.101412, 
    -8.878443, -8.654911, -8.430818, -8.206165, -7.980955, -7.755188, 
    -7.528869, -7.301999, -7.074579, -6.846612, -6.618102, -6.389049, 
    -6.159457, -5.929328, -5.698666, -5.467472, -5.235749, -5.0035, 
    -4.770729, -4.537437, -4.303628, -4.069307, -3.834474, -3.599134, 
    -3.36329, -3.126946, -2.890105, -2.652769, -2.414944, -2.176633, 
    -1.937839, -1.698566, -1.458819, -1.2186, -0.9779146, -0.7367663, 
    -0.4951594, -0.2530979, -0.0105863, 0.2323711, 0.4757699, 0.7196057, 
    0.9638737, 1.208569, 1.453688, 1.699225, 1.945176, 2.191535, 2.438297, 
    2.685458, 2.933012, 3.180955, 3.429281, 3.677984, 3.92706, 4.176504, 
    4.426308, 4.676469, 4.92698, 5.177835, 5.42903, 5.680559, 5.932414, 
    6.184591, 6.437085, 6.689887, 6.942993, 7.196397, 7.450092, 7.704072, 
    7.958331, 8.212863, 8.467661, 8.722718, 8.978029, 9.233587, 9.489386, 
    9.745418, 10.00168, 10.25816, 10.51485, 10.77175, 11.02885, 11.28614, 
    11.54362, 11.80128, 12.05912, 12.31711, 12.57527, 12.83358, 13.09203, 
    13.35062, 13.60934, 13.86819, 14.12715, 14.38622, 14.64539, 14.90465, 
    15.164, 15.42344, 15.68294, 15.94251, 16.20214, 16.46182, 16.72154, 
    16.9813, 17.24109, 17.5009, 17.76072, 18.02055, 18.28038, 18.5402, 
    18.80001, 19.05979, 19.31955, 19.57926, 19.83893, 20.09855, 20.35811, 
    20.61761, 20.87703, 21.13637, 21.39562, 21.65477, 21.91382, 22.17277, 
    22.43159, 22.69029, 22.94886, 23.20729, 23.46558, 23.72371, 23.98168, 
    24.23948, 24.49712, 24.75457, 25.01183, 25.2689, 25.52577, 25.78243, 
    26.03887, 26.2951, 26.55109, 26.80685, 27.06237, 27.31764, 27.57266, 
    27.82742, 28.08191, 28.33612, 28.59006, 28.84371, 29.09706, 29.35012, 
    29.60288, 29.85532, 30.10745, 30.35925, 30.61073, 30.86187, 31.11267, 
    31.36313, 31.61323, 31.86298, 32.11236, 32.36138, 32.61002, 32.85829, 
    33.10617, 33.35366, 33.60077, 33.84746, 34.09376, 34.33964, 34.58511, 
    34.83017, 35.07479, 35.31899, 35.56276, 35.80609, 36.04898, 36.29142, 
    36.53341, 36.77494, 37.01602, 37.25663, 37.49677, 37.73645, 37.97564, 
    38.21436, 38.4526, 38.69035, 38.9276, 39.16436, 39.40063, 39.63639, 
    39.87165, 40.10641, 40.34065, 40.57438, 40.80758, 41.04027, 41.27244, 
    41.50408, 41.73519, 41.96577, 42.19581, 42.42532, 42.65429, 42.88271, 
    43.11059, 43.33792, 43.5647, 43.79094, 44.01662, 44.24174, 44.4663, 
    44.69031, 44.91375, 45.13663, 45.35894, 45.58069, 45.80187, 46.02248, 
    46.24251, 46.46197, 46.68086, 46.89917, 47.1169, 47.33406, 47.55063, 
    47.76662, 47.98203, 48.19686, 48.4111, 48.62476, 48.83783, 49.05032, 
    49.26222, 49.47353, 49.68425, 49.89438, 50.10392, 50.31287, 50.52123, 
    50.729, 50.93617, 51.14276, 51.34875, 51.55415, 51.75896, 51.96317, 
    52.16679, 52.36982, 52.57226, 52.7741, 52.97535, 53.17601, 53.37608, 
    53.57555, 53.77443, 53.97272, 54.17042, 54.36753, 54.56405, 54.75998, 
    54.95532, 55.15007, 55.34423, 55.53781, 55.7308, 55.9232, 56.11501, 
    56.30625, 56.49689, 56.68696, 56.87644, 57.06534, 57.25366, 57.4414, 
    57.62856,
  -36.80576, -36.66573, -36.52526, -36.38437, -36.24305, -36.10129, -35.9591, 
    -35.81647, -35.67341, -35.52991, -35.38596, -35.24157, -35.09674, 
    -34.95145, -34.80572, -34.65954, -34.5129, -34.36581, -34.21826, 
    -34.07025, -33.92178, -33.77285, -33.62345, -33.47359, -33.32325, 
    -33.17245, -33.02118, -32.86943, -32.7172, -32.5645, -32.41131, 
    -32.25764, -32.10349, -31.94886, -31.79374, -31.63812, -31.48202, 
    -31.32542, -31.16833, -31.01074, -30.85265, -30.69406, -30.53497, 
    -30.37537, -30.21527, -30.05466, -29.89354, -29.7319, -29.56976, 
    -29.4071, -29.24392, -29.08022, -28.91601, -28.75127, -28.586, -28.42021, 
    -28.25389, -28.08705, -27.91967, -27.75176, -27.58331, -27.41433, 
    -27.24481, -27.07475, -26.90416, -26.73301, -26.56133, -26.38909, 
    -26.21631, -26.04298, -25.8691, -25.69467, -25.51968, -25.34414, 
    -25.16805, -24.99139, -24.81417, -24.6364, -24.45806, -24.27915, 
    -24.09968, -23.91965, -23.73905, -23.55787, -23.37613, -23.19382, 
    -23.01093, -22.82747, -22.64343, -22.45881, -22.27362, -22.08785, 
    -21.9015, -21.71457, -21.52706, -21.33896, -21.15028, -20.96101, 
    -20.77116, -20.58072, -20.38969, -20.19808, -20.00587, -19.81308, 
    -19.61969, -19.42572, -19.23115, -19.03599, -18.84023, -18.64388, 
    -18.44694, -18.2494, -18.05126, -17.85253, -17.6532, -17.45328, 
    -17.25276, -17.05164, -16.84993, -16.64761, -16.4447, -16.2412, 
    -16.03709, -15.83239, -15.62708, -15.42118, -15.21469, -15.00759, 
    -14.7999, -14.59161, -14.38273, -14.17325, -13.96317, -13.7525, 
    -13.54123, -13.32937, -13.11692, -12.90387, -12.69023, -12.476, 
    -12.26118, -12.04577, -11.82977, -11.61318, -11.39601, -11.17825, 
    -10.95991, -10.74099, -10.52148, -10.30139, -10.08073, -9.859484, 
    -9.637665, -9.415272, -9.192307, -8.96877, -8.744665, -8.519993, 
    -8.294755, -8.068954, -7.842592, -7.615672, -7.388194, -7.160161, 
    -6.931576, -6.702442, -6.47276, -6.242533, -6.011763, -5.780454, 
    -5.548608, -5.316228, -5.083316, -4.849876, -4.615911, -4.381423, 
    -4.146415, -3.910892, -3.674856, -3.43831, -3.201259, -2.963705, 
    -2.725652, -2.487104, -2.248064, -2.008536, -1.768524, -1.528032, 
    -1.287063, -1.045623, -0.8037142, -0.5613418, -0.3185098, -0.07522248, 
    0.1685157, 0.4127003, 0.6573268, 0.9023905, 1.147887, 1.393811, 1.640159, 
    1.886924, 2.134103, 2.38169, 2.62968, 2.878068, 3.12685, 3.376018, 
    3.625569, 3.875497, 4.125796, 4.376461, 4.627487, 4.878866, 5.130595, 
    5.382667, 5.635077, 5.887817, 6.140883, 6.394269, 6.647968, 6.901974, 
    7.156281, 7.410884, 7.665775, 7.920948, 8.176397, 8.432116, 8.688097, 
    8.944335, 9.200824, 9.457555, 9.714522, 9.971721, 10.22914, 10.48678, 
    10.74463, 11.00268, 11.26092, 11.51935, 11.77797, 12.03676, 12.29572, 
    12.55484, 12.81411, 13.07353, 13.33309, 13.59278, 13.85259, 14.11252, 
    14.37257, 14.63271, 14.89295, 15.15328, 15.41369, 15.67418, 15.93473, 
    16.19534, 16.456, 16.7167, 16.97745, 17.23822, 17.49901, 17.75982, 
    18.02063, 18.28144, 18.54225, 18.80304, 19.0638, 19.32454, 19.58524, 
    19.84589, 20.10649, 20.36703, 20.6275, 20.8879, 21.14822, 21.40844, 
    21.66857, 21.9286, 22.18851, 22.44831, 22.70798, 22.96752, 23.22691, 
    23.48616, 23.74525, 24.00419, 24.26295, 24.52154, 24.77994, 25.03816, 
    25.29618, 25.55399, 25.81159, 26.06898, 26.32614, 26.58307, 26.83977, 
    27.09621, 27.35241, 27.60835, 27.86403, 28.11943, 28.37456, 28.62941, 
    28.88397, 29.13823, 29.39218, 29.64583, 29.89917, 30.15218, 30.40487, 
    30.65723, 30.90925, 31.16092, 31.41224, 31.66321, 31.91382, 32.16406, 
    32.41393, 32.66342, 32.91253, 33.16125, 33.40957, 33.6575, 33.90503, 
    34.15214, 34.39884, 34.64512, 34.89098, 35.1364, 35.3814, 35.62595, 
    35.87007, 36.11374, 36.35695, 36.59971, 36.84201, 37.08385, 37.32521, 
    37.5661, 37.80652, 38.04646, 38.28591, 38.52487, 38.76334, 39.00132, 
    39.23879, 39.47576, 39.71223, 39.94818, 40.18362, 40.41855, 40.65295, 
    40.88684, 41.12019, 41.35302, 41.58532, 41.81708, 42.0483, 42.27899, 
    42.50913, 42.73872, 42.96777, 43.19627, 43.42421, 43.6516, 43.87844, 
    44.10471, 44.33042, 44.55557, 44.78015, 45.00417, 45.22762, 45.45049, 
    45.67279, 45.89452, 46.11567, 46.33625, 46.55624, 46.77566, 46.99449, 
    47.21274, 47.4304, 47.64748, 47.86398, 48.07988, 48.2952, 48.50993, 
    48.72406, 48.93761, 49.15056, 49.36292, 49.57469, 49.78586, 49.99644, 
    50.20642, 50.41581, 50.6246, 50.83279, 51.04039, 51.24739, 51.45379, 
    51.6596, 51.86481, 52.06942, 52.27343, 52.47684, 52.67966, 52.88187, 
    53.0835, 53.28452, 53.48494, 53.68477, 53.88401, 54.08264, 54.28069, 
    54.47813, 54.67498, 54.87123, 55.0669, 55.26197, 55.45644, 55.65033, 
    55.84362, 56.03632, 56.22843, 56.41995, 56.61089, 56.80123, 56.99099, 
    57.18016, 57.36875, 57.55676, 57.74418,
  -36.93195, -36.79191, -36.65145, -36.51056, -36.36923, -36.22747, 
    -36.08527, -35.94264, -35.79956, -35.65605, -35.51209, -35.36769, 
    -35.22284, -35.07753, -34.93178, -34.78558, -34.63892, -34.4918, 
    -34.34422, -34.19618, -34.04768, -33.89871, -33.74928, -33.59938, 
    -33.44901, -33.29816, -33.14684, -32.99504, -32.84277, -32.69001, 
    -32.53677, -32.38305, -32.22884, -32.07415, -31.91896, -31.76328, 
    -31.60711, -31.45044, -31.29328, -31.13561, -30.97745, -30.81878, 
    -30.6596, -30.49992, -30.33973, -30.17903, -30.01781, -29.85608, 
    -29.69384, -29.53108, -29.36779, -29.20399, -29.03966, -28.87481, 
    -28.70943, -28.54352, -28.37708, -28.21011, -28.0426, -27.87456, 
    -27.70598, -27.53686, -27.3672, -27.197, -27.02625, -26.85496, -26.68312, 
    -26.51073, -26.33779, -26.16429, -25.99024, -25.81564, -25.64048, 
    -25.46476, -25.28848, -25.11164, -24.93423, -24.75626, -24.57773, 
    -24.39863, -24.21895, -24.03871, -23.8579, -23.67651, -23.49455, 
    -23.31201, -23.12889, -22.9452, -22.76093, -22.57607, -22.39064, 
    -22.20462, -22.01802, -21.83083, -21.64306, -21.4547, -21.26575, 
    -21.07621, -20.88608, -20.69536, -20.50405, -20.31214, -20.11964, 
    -19.92655, -19.73286, -19.53857, -19.34369, -19.14821, -18.95213, 
    -18.75545, -18.55818, -18.3603, -18.16183, -17.96275, -17.76307, 
    -17.56279, -17.36191, -17.16043, -16.95834, -16.75565, -16.55236, 
    -16.34846, -16.14397, -15.93887, -15.73316, -15.52686, -15.31995, 
    -15.11244, -14.90433, -14.69561, -14.48629, -14.27638, -14.06586, 
    -13.85474, -13.64301, -13.4307, -13.21778, -13.00426, -12.79015, 
    -12.57543, -12.36013, -12.14423, -11.92773, -11.71064, -11.49296, 
    -11.27469, -11.05583, -10.83638, -10.61634, -10.39571, -10.17451, 
    -9.952717, -9.730345, -9.507393, -9.283863, -9.059756, -8.835075, 
    -8.609821, -8.383997, -8.157603, -7.930643, -7.703117, -7.47503, 
    -7.246382, -7.017176, -6.787415, -6.5571, -6.326234, -6.094821, 
    -5.862863, -5.630361, -5.39732, -5.163742, -4.929629, -4.694986, 
    -4.459815, -4.224119, -3.987901, -3.751165, -3.513914, -3.276151, 
    -3.03788, -2.799105, -2.559829, -2.320056, -2.07979, -1.839034, 
    -1.597793, -1.35607, -1.113869, -0.8711954, -0.6280527, -0.384445, 
    -0.1403769, 0.1041472, 0.3491228, 0.5945454, 0.8404104, 1.086713, 
    1.333448, 1.580612, 1.828198, 2.076203, 2.32462, 2.573446, 2.822674, 
    3.072299, 3.322317, 3.572722, 3.823508, 4.074669, 4.326201, 4.578098, 
    4.830353, 5.082962, 5.335917, 5.589214, 5.842847, 6.096808, 6.351094, 
    6.605696, 6.86061, 7.115828, 7.371345, 7.627154, 7.883248, 8.139623, 
    8.39627, 8.653182, 8.910356, 9.167781, 9.425453, 9.683364, 9.941508, 
    10.19988, 10.45847, 10.71727, 10.97628, 11.23548, 11.49488, 11.75446, 
    12.01421, 12.27414, 12.53423, 12.79447, 13.05487, 13.3154, 13.57607, 
    13.83686, 14.09778, 14.3588, 14.61993, 14.88116, 15.14247, 15.40387, 
    15.66534, 15.92688, 16.18848, 16.45013, 16.71182, 16.97356, 17.23532, 
    17.4971, 17.7589, 18.02071, 18.28251, 18.54431, 18.80609, 19.06785, 
    19.32957, 19.59126, 19.85291, 20.11449, 20.37602, 20.63748, 20.89887, 
    21.16017, 21.42138, 21.6825, 21.9435, 22.2044, 22.46517, 22.72582, 
    22.98633, 23.2467, 23.50692, 23.76699, 24.02689, 24.28662, 24.54617, 
    24.80553, 25.06471, 25.32368, 25.58245, 25.84101, 26.09934, 26.35745, 
    26.61532, 26.87296, 27.13034, 27.38747, 27.64435, 27.90095, 28.15728, 
    28.41333, 28.66909, 28.92456, 29.17973, 29.4346, 29.68915, 29.94339, 
    30.1973, 30.45088, 30.70412, 30.95702, 31.20957, 31.46177, 31.71361, 
    31.96508, 32.21619, 32.46692, 32.71726, 32.96721, 33.21678, 33.46594, 
    33.7147, 33.96305, 34.21099, 34.45852, 34.70561, 34.95228, 35.19851, 
    35.44431, 35.68966, 35.93456, 36.17902, 36.42301, 36.66655, 36.90961, 
    37.15221, 37.39434, 37.63599, 37.87715, 38.11783, 38.35802, 38.59771, 
    38.83691, 39.0756, 39.31379, 39.55148, 39.78865, 40.0253, 40.26144, 
    40.49705, 40.73214, 40.9667, 41.20073, 41.43422, 41.66718, 41.89959, 
    42.13146, 42.36279, 42.59357, 42.8238, 43.05347, 43.28259, 43.51115, 
    43.73915, 43.96658, 44.19345, 44.41976, 44.64549, 44.87066, 45.09525, 
    45.31926, 45.5427, 45.76556, 45.98784, 46.20954, 46.43065, 46.65118, 
    46.87113, 47.09048, 47.30925, 47.52743, 47.74502, 47.96202, 48.17842, 
    48.39423, 48.60944, 48.82405, 49.03807, 49.2515, 49.46432, 49.67654, 
    49.88817, 50.0992, 50.30962, 50.51944, 50.72867, 50.93729, 51.14531, 
    51.35272, 51.55953, 51.76574, 51.97135, 52.17636, 52.38076, 52.58456, 
    52.78775, 52.99035, 53.19234, 53.39373, 53.59451, 53.7947, 53.99428, 
    54.19326, 54.39164, 54.58942, 54.78661, 54.98319, 55.17917, 55.37456, 
    55.56934, 55.76353, 55.95713, 56.15013, 56.34254, 56.53435, 56.72557, 
    56.91619, 57.10623, 57.29568, 57.48453, 57.6728, 57.86048,
  -37.05865, -36.91862, -36.77816, -36.63727, -36.49594, -36.35418, 
    -36.21198, -36.06934, -35.92626, -35.78274, -35.63877, -35.49435, 
    -35.34949, -35.20417, -35.0584, -34.91217, -34.76549, -34.61835, 
    -34.47075, -34.32268, -34.17414, -34.02515, -33.87568, -33.72574, 
    -33.57533, -33.42444, -33.27308, -33.12124, -32.96892, -32.81611, 
    -32.66282, -32.50905, -32.35478, -32.20003, -32.04478, -31.88904, 
    -31.7328, -31.57607, -31.41883, -31.26109, -31.10285, -30.9441, 
    -30.78485, -30.62508, -30.4648, -30.30401, -30.14271, -29.98088, 
    -29.81854, -29.65568, -29.49229, -29.32838, -29.16395, -28.99898, 
    -28.83349, -28.66746, -28.5009, -28.33381, -28.16617, -27.998, -27.82929, 
    -27.66003, -27.49024, -27.31989, -27.149, -26.97755, -26.80556, 
    -26.63302, -26.45992, -26.28626, -26.11205, -25.93727, -25.76194, 
    -25.58604, -25.40958, -25.23256, -25.05497, -24.87681, -24.69807, 
    -24.51877, -24.3389, -24.15845, -23.97742, -23.79582, -23.61364, 
    -23.43088, -23.24754, -23.06362, -22.87911, -22.69402, -22.50834, 
    -22.32208, -22.13523, -21.94779, -21.75975, -21.57113, -21.38191, 
    -21.1921, -21.0017, -20.81069, -20.6191, -20.4269, -20.23411, -20.04071, 
    -19.84672, -19.65213, -19.45693, -19.26114, -19.06474, -18.86773, 
    -18.67012, -18.47191, -18.27309, -18.07367, -17.87364, -17.67301, 
    -17.47176, -17.26991, -17.06746, -16.86439, -16.66072, -16.45644, 
    -16.25155, -16.04605, -15.83995, -15.63324, -15.42592, -15.21799, 
    -15.00945, -14.80031, -14.59056, -14.38021, -14.16924, -13.95767, 
    -13.7455, -13.53272, -13.31933, -13.10535, -12.89075, -12.67556, 
    -12.45977, -12.24337, -12.02638, -11.80878, -11.59059, -11.37181, 
    -11.15242, -10.93245, -10.71188, -10.49072, -10.26896, -10.04662, 
    -9.823696, -9.600183, -9.376087, -9.151408, -8.926149, -8.700312, 
    -8.473897, -8.246908, -8.019347, -7.791215, -7.562515, -7.333248, 
    -7.103418, -6.873027, -6.642076, -6.41057, -6.178509, -5.945898, 
    -5.712738, -5.479033, -5.244784, -5.009996, -4.774671, -4.538813, 
    -4.302424, -4.065508, -3.828068, -3.590107, -3.351629, -3.112637, 
    -2.873136, -2.633128, -2.392617, -2.151608, -1.910103, -1.668108, 
    -1.425626, -1.182661, -0.9392169, -0.6952987, -0.4509103, -0.2060563, 
    0.03925902, 0.2850311, 0.5312552, 0.7779267, 1.025041, 1.272593, 
    1.520578, 1.768991, 2.017828, 2.267081, 2.516748, 2.766822, 3.017299, 
    3.268172, 3.519436, 3.771087, 4.023118, 4.275523, 4.528297, 4.781435, 
    5.034929, 5.288775, 5.542967, 5.797498, 6.052363, 6.307555, 6.563068, 
    6.818896, 7.075032, 7.331471, 7.588205, 7.845229, 8.102535, 8.360118, 
    8.61797, 8.876084, 9.134456, 9.393076, 9.651939, 9.911037, 10.17037, 
    10.42991, 10.68968, 10.94965, 11.20982, 11.47019, 11.73074, 11.99147, 
    12.25238, 12.51344, 12.77467, 13.03605, 13.29756, 13.55922, 13.821, 
    14.0829, 14.34492, 14.60704, 14.86926, 15.13157, 15.39396, 15.65643, 
    15.91896, 16.18156, 16.44421, 16.7069, 16.96964, 17.2324, 17.49518, 
    17.75798, 18.02079, 18.28359, 18.54639, 18.80917, 19.07193, 19.33465, 
    19.59734, 19.85998, 20.12257, 20.3851, 20.64755, 20.90993, 21.17223, 
    21.43443, 21.69654, 21.95853, 22.22042, 22.48218, 22.74381, 23.00531, 
    23.26666, 23.52786, 23.78891, 24.04978, 24.31049, 24.57101, 24.83135, 
    25.09149, 25.35143, 25.61116, 25.87067, 26.12996, 26.38902, 26.64785, 
    26.90643, 27.16476, 27.42284, 27.68064, 27.93818, 28.19545, 28.45243, 
    28.70911, 28.9655, 29.22159, 29.47737, 29.73283, 29.98797, 30.24279, 
    30.49726, 30.7514, 31.00519, 31.25863, 31.51171, 31.76443, 32.01677, 
    32.26875, 32.52034, 32.77154, 33.02235, 33.27276, 33.52277, 33.77237, 
    34.02156, 34.27033, 34.51868, 34.76659, 35.01408, 35.26112, 35.50772, 
    35.75388, 35.99958, 36.24482, 36.4896, 36.73391, 36.97776, 37.22113, 
    37.46402, 37.70642, 37.94834, 38.18977, 38.43069, 38.67113, 38.91106, 
    39.15047, 39.38939, 39.62778, 39.86566, 40.10302, 40.33985, 40.57616, 
    40.81193, 41.04717, 41.28188, 41.51604, 41.74966, 41.98273, 42.21526, 
    42.44723, 42.67865, 42.90951, 43.13981, 43.36955, 43.59873, 43.82734, 
    44.05538, 44.28285, 44.50975, 44.73607, 44.96182, 45.18699, 45.41158, 
    45.63558, 45.859, 46.08183, 46.30408, 46.52574, 46.74681, 46.96728, 
    47.18716, 47.40645, 47.62515, 47.84324, 48.06074, 48.27764, 48.49394, 
    48.70964, 48.92474, 49.13924, 49.35313, 49.56642, 49.7791, 49.99118, 
    50.20265, 50.41352, 50.62378, 50.83344, 51.04248, 51.25092, 51.45876, 
    51.66598, 51.87259, 52.0786, 52.284, 52.48879, 52.69298, 52.89655, 
    53.09952, 53.30188, 53.50364, 53.70478, 53.90532, 54.10526, 54.30458, 
    54.5033, 54.70142, 54.89893, 55.09584, 55.29215, 55.48785, 55.68295, 
    55.87745, 56.07135, 56.26464, 56.45734, 56.64944, 56.84095, 57.03185, 
    57.22216, 57.41188, 57.60101, 57.78954, 57.97747,
  -37.18589, -37.04587, -36.90541, -36.76452, -36.6232, -36.48143, -36.33923, 
    -36.19659, -36.0535, -35.90997, -35.766, -35.62157, -35.47669, -35.33136, 
    -35.18557, -35.03933, -34.89262, -34.74546, -34.59783, -34.44974, 
    -34.30118, -34.15215, -34.00266, -33.85268, -33.70223, -33.55131, 
    -33.39991, -33.24802, -33.09565, -32.9428, -32.78946, -32.63564, 
    -32.48132, -32.32651, -32.1712, -32.0154, -31.85909, -31.70229, 
    -31.54499, -31.38718, -31.22886, -31.07004, -30.91071, -30.75086, 
    -30.5905, -30.42962, -30.26822, -30.10631, -29.94387, -29.78091, 
    -29.61743, -29.45341, -29.28887, -29.12379, -28.95819, -28.79205, 
    -28.62537, -28.45815, -28.29039, -28.12209, -27.95325, -27.78386, 
    -27.61392, -27.44344, -27.2724, -27.10081, -26.92867, -26.75597, 
    -26.58271, -26.40889, -26.23451, -26.05957, -25.88407, -25.708, 
    -25.53136, -25.35415, -25.17637, -24.99802, -24.8191, -24.6396, 
    -24.45953, -24.27887, -24.09764, -23.91582, -23.73343, -23.55045, 
    -23.36688, -23.18273, -22.99799, -22.81266, -22.62675, -22.44024, 
    -22.25313, -22.06544, -21.87715, -21.68826, -21.49878, -21.30869, 
    -21.11801, -20.92673, -20.73485, -20.54237, -20.34928, -20.15559, 
    -19.96129, -19.76639, -19.57088, -19.37477, -19.17805, -18.98072, 
    -18.78278, -18.58423, -18.38507, -18.1853, -17.98492, -17.78393, 
    -17.58233, -17.38011, -17.17729, -16.97385, -16.76979, -16.56513, 
    -16.35985, -16.15396, -15.94745, -15.74033, -15.5326, -15.32425, 
    -15.11529, -14.90572, -14.69554, -14.48474, -14.27333, -14.06131, 
    -13.84868, -13.63544, -13.42159, -13.20713, -12.99207, -12.77639, 
    -12.56011, -12.34322, -12.12572, -11.90762, -11.68892, -11.46962, 
    -11.24971, -11.02921, -10.8081, -10.5864, -10.3641, -10.14121, -9.917728, 
    -9.693652, -9.468987, -9.243733, -9.017894, -8.791471, -8.564465, 
    -8.336878, -8.108712, -7.879971, -7.650655, -7.420768, -7.19031, 
    -6.959287, -6.727697, -6.495546, -6.262836, -6.029568, -5.795746, 
    -5.561373, -5.326451, -5.090983, -4.854974, -4.618424, -4.381339, 
    -4.14372, -3.905572, -3.666897, -3.4277, -3.187983, -2.947751, -2.707006, 
    -2.465754, -2.223997, -1.981739, -1.738985, -1.495739, -1.252004, 
    -1.007785, -0.7630866, -0.5179124, -0.2722672, -0.02615537, 0.2204184, 
    0.4674495, 0.7149333, 0.9628649, 1.211239, 1.460052, 1.709298, 1.958971, 
    2.209068, 2.459582, 2.710508, 2.961841, 3.213576, 3.465707, 3.718228, 
    3.971134, 4.22442, 4.478078, 4.732105, 4.986493, 5.241237, 5.49633, 
    5.751767, 6.007542, 6.263647, 6.520078, 6.776828, 7.033889, 7.291257, 
    7.548924, 7.806884, 8.065131, 8.323657, 8.582456, 8.84152, 9.100844, 
    9.360421, 9.620243, 9.880304, 10.1406, 10.40111, 10.66185, 10.92279, 
    11.18394, 11.44529, 11.70682, 11.96853, 12.23042, 12.49248, 12.75469, 
    13.01706, 13.27957, 13.54222, 13.805, 14.0679, 14.33091, 14.59403, 
    14.85725, 15.12057, 15.38396, 15.64744, 15.91098, 16.17458, 16.43824, 
    16.70194, 16.96568, 17.22945, 17.49324, 17.75705, 18.02087, 18.28468, 
    18.54849, 18.81228, 19.07604, 19.33978, 19.60347, 19.86712, 20.13071, 
    20.39425, 20.65771, 20.92109, 21.18439, 21.4476, 21.7107, 21.9737, 
    22.23658, 22.49934, 22.76196, 23.02445, 23.2868, 23.54899, 23.81102, 
    24.07288, 24.33456, 24.59607, 24.85738, 25.1185, 25.37941, 25.64011, 
    25.90059, 26.16085, 26.42087, 26.68066, 26.94019, 27.19948, 27.4585, 
    27.71726, 27.97574, 28.23394, 28.49185, 28.74947, 29.00679, 29.26381, 
    29.52051, 29.77689, 30.03294, 30.28866, 30.54404, 30.79908, 31.05377, 
    31.3081, 31.56207, 31.81567, 32.0689, 32.32174, 32.5742, 32.82627, 
    33.07794, 33.32921, 33.58007, 33.83052, 34.08055, 34.33016, 34.57933, 
    34.82808, 35.07638, 35.32425, 35.57166, 35.81861, 36.06512, 36.31116, 
    36.55672, 36.80183, 37.04645, 37.29059, 37.53425, 37.77742, 38.02009, 
    38.26227, 38.50395, 38.74512, 38.98579, 39.22594, 39.46557, 39.70469, 
    39.94328, 40.18134, 40.41888, 40.65588, 40.89234, 41.12827, 41.36365, 
    41.59848, 41.83277, 42.06651, 42.29968, 42.53231, 42.76437, 42.99587, 
    43.2268, 43.45717, 43.68697, 43.91619, 44.14484, 44.37292, 44.60041, 
    44.82732, 45.05366, 45.2794, 45.50457, 45.72914, 45.95312, 46.17651, 
    46.39931, 46.62151, 46.84312, 47.06413, 47.28454, 47.50435, 47.72356, 
    47.94216, 48.16017, 48.37757, 48.59436, 48.81055, 49.02613, 49.2411, 
    49.45546, 49.66922, 49.88236, 50.09489, 50.30682, 50.51813, 50.72882, 
    50.93892, 51.14839, 51.35725, 51.5655, 51.77313, 51.98016, 52.18657, 
    52.39236, 52.59754, 52.80211, 53.00607, 53.20941, 53.41214, 53.61426, 
    53.81577, 54.01666, 54.21695, 54.41662, 54.61568, 54.81413, 55.01197, 
    55.20921, 55.40583, 55.60185, 55.79726, 55.99207, 56.18627, 56.37986, 
    56.57285, 56.76524, 56.95703, 57.14822, 57.3388, 57.52879, 57.71818, 
    57.90697, 58.09517,
  -37.31366, -37.17365, -37.0332, -36.89231, -36.75099, -36.60923, -36.46703, 
    -36.32438, -36.1813, -36.03776, -35.89378, -35.74934, -35.60445, 
    -35.45911, -35.3133, -35.16705, -35.02032, -34.87314, -34.72549, 
    -34.57738, -34.42879, -34.27974, -34.13021, -33.9802, -33.82972, 
    -33.67876, -33.52732, -33.37539, -33.22298, -33.07008, -32.9167, 
    -32.76282, -32.60845, -32.45359, -32.29822, -32.14236, -31.986, 
    -31.82913, -31.67176, -31.51388, -31.35549, -31.1966, -31.03718, 
    -30.87726, -30.71681, -30.55585, -30.39437, -30.23236, -30.06983, 
    -29.90678, -29.74319, -29.57908, -29.41443, -29.24925, -29.08353, 
    -28.91727, -28.75048, -28.58314, -28.41526, -28.24684, -28.07786, 
    -27.90834, -27.73827, -27.56764, -27.39647, -27.22473, -27.05244, 
    -26.87959, -26.70617, -26.5322, -26.35766, -26.18255, -26.00687, 
    -25.83063, -25.65381, -25.47643, -25.29846, -25.11993, -24.94081, 
    -24.76112, -24.58084, -24.39998, -24.21854, -24.03652, -23.8539, 
    -23.67071, -23.48692, -23.30254, -23.11757, -22.932, -22.74585, 
    -22.55909, -22.37174, -22.18379, -21.99524, -21.8061, -21.61635, -21.426, 
    -21.23504, -21.04348, -20.85131, -20.65854, -20.46516, -20.27117, 
    -20.07658, -19.88137, -19.68555, -19.48912, -19.29208, -19.09442, 
    -18.89615, -18.69727, -18.49777, -18.29766, -18.09693, -17.89558, 
    -17.69361, -17.49103, -17.28784, -17.08402, -16.87959, -16.67453, 
    -16.46886, -16.26257, -16.05567, -15.84814, -15.63999, -15.43123, 
    -15.22185, -15.01185, -14.80123, -14.58999, -14.37814, -14.16567, 
    -13.95259, -13.73888, -13.52457, -13.30963, -13.09409, -12.87793, 
    -12.66115, -12.44377, -12.22577, -12.00717, -11.78795, -11.56813, 
    -11.3477, -11.12666, -10.90502, -10.68278, -10.45994, -10.23649, 
    -10.01245, -9.787807, -9.562571, -9.33674, -9.110318, -8.883306, 
    -8.655705, -8.427518, -8.198747, -7.969393, -7.73946, -7.508948, 
    -7.277861, -7.046201, -6.81397, -6.581172, -6.347807, -6.11388, 
    -5.879393, -5.644348, -5.408749, -5.172599, -4.9359, -4.698656, -4.46087, 
    -4.222545, -3.983685, -3.744292, -3.504371, -3.263925, -3.022958, 
    -2.781472, -2.539473, -2.296964, -2.053949, -1.810431, -1.566416, 
    -1.321907, -1.076908, -0.8314233, -0.5854581, -0.3390164, -0.09210275, 
    0.1552782, 0.4031219, 0.6514234, 0.900178, 1.149381, 1.399027, 1.649111, 
    1.899628, 2.150573, 2.40194, 2.653725, 2.905921, 3.158525, 3.411528, 
    3.664927, 3.918715, 4.172887, 4.427437, 4.682359, 4.937647, 5.193295, 
    5.449297, 5.705647, 5.962339, 6.219366, 6.476722, 6.7344, 6.992395, 
    7.2507, 7.509307, 7.768211, 8.027405, 8.286881, 8.546636, 8.806658, 
    9.066943, 9.327484, 9.588274, 9.849305, 10.11057, 10.37206, 10.63378, 
    10.8957, 11.15784, 11.42017, 11.68269, 11.94539, 12.20828, 12.47133, 
    12.73454, 12.99791, 13.26142, 13.52507, 13.78885, 14.05276, 14.31678, 
    14.58091, 14.84514, 15.10947, 15.37388, 15.63836, 15.90292, 16.16754, 
    16.43221, 16.69693, 16.96169, 17.22648, 17.49129, 17.75611, 18.02095, 
    18.28578, 18.5506, 18.81541, 19.08019, 19.34495, 19.60966, 19.87432, 
    20.13893, 20.40348, 20.66795, 20.93235, 21.19666, 21.46088, 21.72499, 
    21.98899, 22.25288, 22.51664, 22.78027, 23.04376, 23.30711, 23.57029, 
    23.83332, 24.09617, 24.35885, 24.62134, 24.88364, 25.14574, 25.40764, 
    25.66932, 25.93077, 26.192, 26.453, 26.71375, 26.97425, 27.23449, 
    27.49447, 27.75418, 28.01361, 28.27276, 28.53162, 28.79018, 29.04844, 
    29.30638, 29.56401, 29.82131, 30.07829, 30.33493, 30.59122, 30.84717, 
    31.10276, 31.35799, 31.61285, 31.86734, 32.12146, 32.37518, 32.62852, 
    32.88146, 33.134, 33.38613, 33.63785, 33.88915, 34.14003, 34.39048, 
    34.64049, 34.89007, 35.1392, 35.38788, 35.63611, 35.88388, 36.13119, 
    36.37803, 36.6244, 36.87029, 37.1157, 37.36061, 37.60505, 37.84898, 
    38.09242, 38.33536, 38.57779, 38.81971, 39.06111, 39.30199, 39.54236, 
    39.7822, 40.0215, 40.26028, 40.49852, 40.73622, 40.97338, 41.20999, 
    41.44605, 41.68156, 41.91652, 42.15092, 42.38476, 42.61803, 42.85074, 
    43.08288, 43.31445, 43.54545, 43.77587, 44.00571, 44.23497, 44.46365, 
    44.69175, 44.91925, 45.14618, 45.3725, 45.59824, 45.82338, 46.04793, 
    46.27188, 46.49523, 46.71798, 46.94012, 47.16167, 47.38261, 47.60294, 
    47.82267, 48.04179, 48.2603, 48.4782, 48.69548, 48.91216, 49.12822, 
    49.34367, 49.55851, 49.77273, 49.98633, 50.19932, 50.41169, 50.62345, 
    50.83459, 51.04511, 51.25501, 51.46429, 51.67296, 51.88101, 52.08844, 
    52.29525, 52.50144, 52.70701, 52.91196, 53.1163, 53.32002, 53.52312, 
    53.72561, 53.92747, 54.12872, 54.32935, 54.52937, 54.72877, 54.92756, 
    55.12573, 55.32329, 55.52023, 55.71657, 55.91229, 56.1074, 56.3019, 
    56.49579, 56.68908, 56.88175, 57.07382, 57.26529, 57.45615, 57.6464, 
    57.83606, 58.02511, 58.21356,
  -37.44196, -37.30196, -37.16152, -37.02064, -36.87933, -36.73757, 
    -36.59537, -36.45273, -36.30964, -36.1661, -36.02211, -35.87767, 
    -35.73277, -35.58742, -35.4416, -35.29533, -35.14859, -35.00139, 
    -34.85372, -34.70559, -34.55698, -34.40789, -34.25834, -34.1083, 
    -33.95779, -33.8068, -33.65532, -33.50336, -33.35091, -33.19796, 
    -33.04453, -32.89061, -32.73619, -32.58127, -32.42585, -32.26993, 
    -32.11351, -31.95658, -31.79915, -31.6412, -31.48274, -31.32377, 
    -31.16429, -31.00428, -30.84376, -30.68271, -30.52115, -30.35905, 
    -30.19643, -30.03328, -29.8696, -29.70539, -29.54063, -29.37535, 
    -29.20952, -29.04315, -28.87624, -28.70879, -28.54079, -28.37224, 
    -28.20314, -28.03349, -27.86328, -27.69252, -27.5212, -27.34932, 
    -27.17688, -27.00388, -26.83031, -26.65618, -26.48147, -26.3062, 
    -26.13036, -25.95395, -25.77695, -25.59939, -25.42124, -25.24252, 
    -25.06321, -24.88332, -24.70285, -24.52179, -24.34014, -24.15791, 
    -23.97508, -23.79166, -23.60765, -23.42305, -23.23785, -23.05205, 
    -22.86565, -22.67866, -22.49106, -22.30286, -22.11406, -21.92465, 
    -21.73463, -21.54401, -21.35278, -21.16095, -20.9685, -20.77544, 
    -20.58177, -20.38748, -20.19258, -19.99707, -19.80094, -19.60419, 
    -19.40683, -19.20885, -19.01025, -18.81103, -18.61119, -18.41073, 
    -18.20965, -18.00795, -17.80563, -17.60268, -17.39911, -17.19492, 
    -16.9901, -16.78467, -16.5786, -16.37192, -16.16461, -15.95667, 
    -15.74812, -15.53893, -15.32913, -15.1187, -14.90765, -14.69597, 
    -14.48367, -14.27075, -14.05721, -13.84304, -13.62826, -13.41285, 
    -13.19682, -12.98018, -12.76291, -12.54503, -12.32653, -12.10742, 
    -11.88769, -11.66735, -11.44639, -11.22482, -11.00265, -10.77986, 
    -10.55647, -10.33247, -10.10786, -9.882655, -9.656845, -9.430436, 
    -9.203429, -8.975826, -8.747628, -8.518839, -8.289458, -8.059489, 
    -7.828935, -7.597797, -7.366077, -7.133778, -6.900903, -6.667453, 
    -6.433432, -6.198842, -5.963686, -5.727967, -5.491687, -5.25485, 
    -5.017459, -4.779517, -4.541026, -4.301991, -4.062414, -3.8223, 
    -3.581651, -3.340471, -3.098764, -2.856533, -2.613783, -2.370517, 
    -2.126739, -1.882453, -1.637664, -1.392375, -1.146591, -0.9003159, 
    -0.6535544, -0.4063109, -0.15859, 0.08960369, 0.3382654, 0.5873904, 
    0.8369737, 1.087011, 1.337496, 1.588424, 1.839791, 2.09159, 2.343818, 
    2.596467, 2.849533, 3.10301, 3.356894, 3.611176, 3.865853, 4.120919, 
    4.376367, 4.632191, 4.888387, 5.144946, 5.401864, 5.659134, 5.91675, 
    6.174705, 6.432993, 6.691608, 6.950544, 7.209793, 7.469348, 7.729204, 
    7.989353, 8.249789, 8.510505, 8.771493, 9.032747, 9.294261, 9.556026, 
    9.818036, 10.08028, 10.34276, 10.60546, 10.86838, 11.1315, 11.39483, 
    11.65835, 11.92205, 12.18594, 12.44999, 12.71421, 12.97858, 13.24311, 
    13.50777, 13.77257, 14.03749, 14.30253, 14.56768, 14.83293, 15.09827, 
    15.3637, 15.62921, 15.89479, 16.16044, 16.42613, 16.69188, 16.95766, 
    17.22348, 17.48931, 17.75517, 18.02103, 18.28689, 18.55274, 18.81857, 
    19.08438, 19.35016, 19.6159, 19.88159, 20.14722, 20.41279, 20.67829, 
    20.94371, 21.20904, 21.47427, 21.7394, 22.00443, 22.26933, 22.5341, 
    22.79874, 23.06325, 23.32759, 23.59179, 23.85582, 24.11967, 24.38335, 
    24.64684, 24.91013, 25.17323, 25.43611, 25.69877, 25.96122, 26.22342, 
    26.4854, 26.74712, 27.0086, 27.26981, 27.53075, 27.79143, 28.05182, 
    28.31192, 28.57173, 28.83124, 29.09044, 29.34932, 29.60789, 29.86612, 
    30.12402, 30.38158, 30.6388, 30.89566, 31.15216, 31.4083, 31.66407, 
    31.91945, 32.17446, 32.42907, 32.68329, 32.93711, 33.19053, 33.44353, 
    33.69611, 33.94827, 34.2, 34.4513, 34.70216, 34.95257, 35.20254, 
    35.45205, 35.7011, 35.94969, 36.19781, 36.44545, 36.69262, 36.9393, 
    37.1855, 37.43121, 37.67642, 37.92113, 38.16533, 38.40903, 38.65222, 
    38.89489, 39.13703, 39.37866, 39.61975, 39.86032, 40.10035, 40.33984, 
    40.57879, 40.81719, 41.05505, 41.29235, 41.5291, 41.76529, 42.00092, 
    42.23599, 42.47049, 42.70442, 42.93778, 43.17056, 43.40277, 43.6344, 
    43.86544, 44.09591, 44.32578, 44.55507, 44.78376, 45.01187, 45.23938, 
    45.46629, 45.6926, 45.91832, 46.14343, 46.36794, 46.59185, 46.81514, 
    47.03783, 47.25991, 47.48138, 47.70224, 47.92249, 48.14212, 48.36114, 
    48.57954, 48.79732, 49.01449, 49.23104, 49.44696, 49.66227, 49.87696, 
    50.09103, 50.30447, 50.5173, 50.7295, 50.94107, 51.15203, 51.36236, 
    51.57206, 51.78115, 51.98961, 52.19744, 52.40465, 52.61124, 52.8172, 
    53.02254, 53.22726, 53.43135, 53.63482, 53.83767, 54.0399, 54.2415, 
    54.44248, 54.64285, 54.84259, 55.04171, 55.24021, 55.43809, 55.63536, 
    55.832, 56.02804, 56.22345, 56.41825, 56.61244, 56.80602, 56.99898, 
    57.19133, 57.38307, 57.57421, 57.76473, 57.95465, 58.14396, 58.33267,
  -37.5708, -37.43081, -37.29038, -37.14951, -37.00821, -36.86646, -36.72426, 
    -36.58162, -36.43853, -36.29499, -36.151, -36.00656, -35.86165, 
    -35.71629, -35.57047, -35.42418, -35.27744, -35.13022, -34.98253, 
    -34.83437, -34.68575, -34.53664, -34.38706, -34.237, -34.08645, 
    -33.93542, -33.78391, -33.63191, -33.47942, -33.32644, -33.17297, 
    -33.019, -32.86453, -32.70956, -32.55409, -32.39812, -32.24164, 
    -32.08465, -31.92715, -31.76914, -31.61062, -31.45158, -31.29202, 
    -31.13194, -30.97134, -30.81021, -30.64856, -30.48638, -30.32367, 
    -30.16043, -29.99665, -29.83234, -29.66749, -29.5021, -29.33616, 
    -29.16969, -29.00266, -28.83509, -28.66697, -28.4983, -28.32907, 
    -28.15929, -27.98896, -27.81806, -27.6466, -27.47458, -27.302, -27.12885, 
    -26.95513, -26.78084, -26.60598, -26.43054, -26.25453, -26.07795, 
    -25.90078, -25.72304, -25.54471, -25.3658, -25.18631, -25.00623, 
    -24.82556, -24.6443, -24.46244, -24.28, -24.09696, -23.91333, -23.7291, 
    -23.54427, -23.35884, -23.17281, -22.98617, -22.79894, -22.61109, 
    -22.42264, -22.23359, -22.04392, -21.85364, -21.66275, -21.47125, 
    -21.27913, -21.0864, -20.89306, -20.69909, -20.50451, -20.30931, 
    -20.11349, -19.91706, -19.72, -19.52231, -19.32401, -19.12508, -18.92552, 
    -18.72535, -18.52454, -18.32311, -18.12105, -17.91837, -17.71506, 
    -17.51112, -17.30655, -17.10136, -16.89553, -16.68908, -16.48199, 
    -16.27428, -16.06594, -15.85697, -15.64737, -15.43714, -15.22628, 
    -15.01479, -14.80268, -14.58993, -14.37656, -14.16256, -13.94793, 
    -13.73267, -13.51679, -13.30029, -13.08315, -12.8654, -12.64702, 
    -12.42801, -12.20839, -11.98815, -11.76728, -11.5458, -11.3237, 
    -11.10098, -10.87765, -10.65371, -10.42915, -10.20398, -9.978204, 
    -9.75182, -9.524829, -9.297235, -9.069038, -8.840241, -8.610846, 
    -8.380855, -8.150269, -7.91909, -7.687322, -7.454967, -7.222026, 
    -6.988503, -6.754399, -6.519718, -6.284461, -6.048634, -5.812236, 
    -5.575272, -5.337745, -5.099658, -4.861012, -4.621814, -4.382064, 
    -4.141768, -3.900927, -3.659546, -3.417628, -3.175177, -2.932196, 
    -2.68869, -2.444663, -2.200117, -1.955059, -1.70949, -1.463417, 
    -1.216842, -0.9697714, -0.7222083, -0.4741577, -0.225624, 0.02338787, 
    0.2728733, 0.5228274, 0.7732453, 1.024122, 1.275452, 1.527231, 1.779454, 
    2.032114, 2.285207, 2.538728, 2.79267, 3.047028, 3.301797, 3.556971, 
    3.812543, 4.068509, 4.324862, 4.581596, 4.838706, 5.096184, 5.354024, 
    5.612222, 5.87077, 6.129661, 6.388889, 6.648448, 6.908331, 7.168532, 
    7.429043, 7.689859, 7.950971, 8.212374, 8.47406, 8.736022, 8.998254, 
    9.260748, 9.523497, 9.786493, 10.04973, 10.3132, 10.5769, 10.84081, 
    11.10494, 11.36927, 11.63379, 11.89851, 12.1634, 12.42847, 12.6937, 
    12.95909, 13.22464, 13.49032, 13.75614, 14.02208, 14.28815, 14.55432, 
    14.8206, 15.08698, 15.35344, 15.61998, 15.88659, 16.15327, 16.42, 
    16.68678, 16.9536, 17.22045, 17.48732, 17.75421, 18.02111, 18.28801, 
    18.55489, 18.82176, 19.08861, 19.35542, 19.62219, 19.88892, 20.15558, 
    20.42219, 20.68871, 20.95516, 21.22153, 21.48779, 21.75395, 22.01999, 
    22.28592, 22.55172, 22.81738, 23.0829, 23.34826, 23.61347, 23.87851, 
    24.14338, 24.40807, 24.67256, 24.93686, 25.20095, 25.46483, 25.72849, 
    25.99193, 26.25513, 26.51808, 26.78079, 27.04324, 27.30543, 27.56735, 
    27.82899, 28.09035, 28.35142, 28.61219, 28.87265, 29.1328, 29.39263, 
    29.65214, 29.91131, 30.17015, 30.42864, 30.68678, 30.94457, 31.20199, 
    31.45904, 31.71571, 31.97201, 32.22791, 32.48342, 32.73853, 32.99323, 
    33.24753, 33.5014, 33.75486, 34.00788, 34.26047, 34.51263, 34.76434, 
    35.01559, 35.2664, 35.51674, 35.76662, 36.01603, 36.26497, 36.51343, 
    36.7614, 37.00889, 37.25588, 37.50238, 37.74837, 37.99386, 38.23883, 
    38.4833, 38.72725, 38.97066, 39.21356, 39.45593, 39.69777, 39.93906, 
    40.17981, 40.42002, 40.65969, 40.8988, 41.13736, 41.37535, 41.61279, 
    41.84967, 42.08598, 42.32171, 42.55688, 42.79147, 43.02548, 43.25891, 
    43.49176, 43.72402, 43.9557, 44.18678, 44.41727, 44.64717, 44.87647, 
    45.10518, 45.33327, 45.56078, 45.78767, 46.01396, 46.23964, 46.46471, 
    46.68917, 46.91302, 47.13625, 47.35887, 47.58088, 47.80226, 48.02303, 
    48.24317, 48.4627, 48.6816, 48.89988, 49.11754, 49.33458, 49.55098, 
    49.76677, 49.98192, 50.19645, 50.41035, 50.62363, 50.83627, 51.04829, 
    51.25968, 51.47044, 51.68057, 51.89007, 52.09894, 52.30718, 52.51479, 
    52.72178, 52.92813, 53.13386, 53.33895, 53.54342, 53.74726, 53.95047, 
    54.15306, 54.35501, 54.55635, 54.75705, 54.95713, 55.15659, 55.35542, 
    55.55362, 55.75121, 55.94817, 56.14451, 56.34023, 56.53534, 56.72982, 
    56.92368, 57.11693, 57.30956, 57.50158, 57.69299, 57.88378, 58.07396, 
    58.26353, 58.45249,
  -37.70018, -37.5602, -37.41979, -37.27893, -37.13763, -36.9959, -36.85371, 
    -36.71107, -36.56799, -36.42445, -36.28046, -36.13601, -35.9911, 
    -35.84574, -35.69991, -35.55361, -35.40685, -35.25962, -35.11192, 
    -34.96375, -34.8151, -34.66597, -34.51637, -34.36628, -34.21571, 
    -34.06465, -33.91311, -33.76107, -33.60855, -33.45553, -33.30201, 
    -33.148, -32.99348, -32.83847, -32.68295, -32.52692, -32.37039, 
    -32.21334, -32.05578, -31.89771, -31.73912, -31.58001, -31.42038, 
    -31.26023, -31.09955, -30.93835, -30.77662, -30.61435, -30.45155, 
    -30.28822, -30.12435, -29.95994, -29.79499, -29.6295, -29.46346, 
    -29.29688, -29.12975, -28.96206, -28.79382, -28.62503, -28.45568, 
    -28.28577, -28.11531, -27.94428, -27.77268, -27.60052, -27.42779, 
    -27.2545, -27.08063, -26.90618, -26.73116, -26.55557, -26.3794, 
    -26.20264, -26.0253, -25.84739, -25.66888, -25.48979, -25.3101, 
    -25.12983, -24.94897, -24.76751, -24.58545, -24.40281, -24.21956, 
    -24.03571, -23.85126, -23.6662, -23.48055, -23.29428, -23.10741, 
    -22.91994, -22.73185, -22.54315, -22.35384, -22.16391, -21.97337, 
    -21.78222, -21.59044, -21.39805, -21.20504, -21.01141, -20.81716, 
    -20.62228, -20.42678, -20.23066, -20.03391, -19.83653, -19.63853, 
    -19.4399, -19.24064, -19.04076, -18.84024, -18.63909, -18.43731, 
    -18.2349, -18.03185, -17.82818, -17.62387, -17.41893, -17.21335, 
    -17.00714, -16.80029, -16.59281, -16.3847, -16.17595, -15.96657, 
    -15.75655, -15.54589, -15.3346, -15.12268, -14.91012, -14.69693, 
    -14.4831, -14.26864, -14.05355, -13.83782, -13.62147, -13.40448, 
    -13.18686, -12.96861, -12.74973, -12.53022, -12.31009, -12.08933, 
    -11.86794, -11.64593, -11.42329, -11.20004, -10.97616, -10.75166, 
    -10.52654, -10.30081, -10.07446, -9.847501, -9.619926, -9.391743, 
    -9.162951, -8.933552, -8.703548, -8.472943, -8.241736, -8.009933, 
    -7.777532, -7.544538, -7.310952, -7.076777, -6.842017, -6.606672, 
    -6.370747, -6.134243, -5.897164, -5.659512, -5.421291, -5.182503, 
    -4.943152, -4.703241, -4.462774, -4.221752, -3.980181, -3.738064, 
    -3.495403, -3.252204, -3.008469, -2.764203, -2.519409, -2.274091, 
    -2.028255, -1.781902, -1.535039, -1.287669, -1.039797, -0.7914271, 
    -0.5425639, -0.293212, -0.04337627, 0.2069386, 0.4577276, 0.7089859, 
    0.9607084, 1.21289, 1.465526, 1.71861, 1.972137, 2.226103, 2.480501, 
    2.735326, 2.990571, 3.246233, 3.502304, 3.758779, 4.015652, 4.272917, 
    4.530568, 4.788598, 5.047002, 5.305773, 5.564906, 5.824392, 6.084227, 
    6.344403, 6.604913, 6.865752, 7.126913, 7.388388, 7.650171, 7.912254, 
    8.174632, 8.437297, 8.700241, 8.963458, 9.22694, 9.490681, 9.754673, 
    10.01891, 10.28338, 10.54808, 10.813, 11.07814, 11.34348, 11.60902, 
    11.87475, 12.14066, 12.40675, 12.67301, 12.93943, 13.206, 13.47271, 
    13.73956, 14.00654, 14.27364, 14.54085, 14.80817, 15.07558, 15.34308, 
    15.61067, 15.87832, 16.14604, 16.41381, 16.68164, 16.9495, 17.2174, 
    17.48532, 17.75325, 18.02119, 18.28913, 18.55707, 18.82498, 19.09287, 
    19.36073, 19.62855, 19.89631, 20.16402, 20.43167, 20.69924, 20.96672, 
    21.23412, 21.50142, 21.76862, 22.0357, 22.30266, 22.56949, 22.83618, 
    23.10272, 23.36912, 23.63535, 23.90141, 24.1673, 24.433, 24.69851, 
    24.96382, 25.22892, 25.49381, 25.75847, 26.02291, 26.2871, 26.55106, 
    26.81475, 27.0782, 27.34137, 27.60427, 27.86689, 28.12922, 28.39126, 
    28.65299, 28.91442, 29.17553, 29.43632, 29.69678, 29.9569, 30.21668, 
    30.47611, 30.73518, 30.9939, 31.25224, 31.51021, 31.7678, 32.02501, 
    32.28182, 32.53823, 32.79424, 33.04983, 33.30501, 33.55977, 33.8141, 
    34.068, 34.32145, 34.57447, 34.82703, 35.07914, 35.33079, 35.58197, 
    35.83269, 36.08293, 36.33269, 36.58196, 36.83075, 37.07904, 37.32683, 
    37.57412, 37.8209, 38.06718, 38.31293, 38.55817, 38.80288, 39.04706, 
    39.29071, 39.53382, 39.7764, 40.01843, 40.25991, 40.50085, 40.74123, 
    40.98105, 41.22031, 41.45901, 41.69714, 41.9347, 42.17169, 42.4081, 
    42.64394, 42.87919, 43.11386, 43.34794, 43.58143, 43.81433, 44.04664, 
    44.27835, 44.50946, 44.73997, 44.96988, 45.19918, 45.42788, 45.65597, 
    45.88344, 46.11031, 46.33656, 46.56219, 46.78721, 47.01161, 47.23539, 
    47.45855, 47.68109, 47.903, 48.12429, 48.34495, 48.56499, 48.7844, 
    49.00317, 49.22132, 49.43885, 49.65574, 49.87199, 50.08762, 50.30261, 
    50.51697, 50.73069, 50.94379, 51.15624, 51.36807, 51.57925, 51.78981, 
    51.99973, 52.20901, 52.41766, 52.62568, 52.83305, 53.0398, 53.24591, 
    53.45139, 53.65623, 53.86044, 54.06401, 54.26696, 54.46927, 54.67095, 
    54.872, 55.07242, 55.27221, 55.47136, 55.6699, 55.8678, 56.06507, 
    56.26172, 56.45775, 56.65315, 56.84792, 57.04208, 57.23561, 57.42852, 
    57.62082, 57.8125, 58.00355, 58.194, 58.38382, 58.57304,
  -37.8301, -37.69014, -37.54974, -37.4089, -37.26762, -37.12589, -36.98371, 
    -36.84108, -36.698, -36.55447, -36.41048, -36.26603, -36.12112, 
    -35.97575, -35.82992, -35.68362, -35.53685, -35.3896, -35.24189, 
    -35.0937, -34.94503, -34.79589, -34.64626, -34.49615, -34.34556, 
    -34.19447, -34.0429, -33.89083, -33.73827, -33.58522, -33.43166, 
    -33.27761, -33.12305, -32.96799, -32.81242, -32.65635, -32.49976, 
    -32.34266, -32.18504, -32.02691, -31.86825, -31.70908, -31.54938, 
    -31.38916, -31.22841, -31.06713, -30.90532, -30.74297, -30.58009, 
    -30.41667, -30.25271, -30.0882, -29.92316, -29.75757, -29.59142, 
    -29.42474, -29.25749, -29.0897, -28.92134, -28.75243, -28.58296, 
    -28.41293, -28.24234, -28.07117, -27.89945, -27.72715, -27.55428, 
    -27.38083, -27.20682, -27.03222, -26.85705, -26.68129, -26.50496, 
    -26.32804, -26.15053, -25.97243, -25.79375, -25.61448, -25.43461, 
    -25.25415, -25.07309, -24.89144, -24.70918, -24.52632, -24.34286, 
    -24.1588, -23.97414, -23.78886, -23.60298, -23.41648, -23.22938, 
    -23.04166, -22.85333, -22.66438, -22.47482, -22.28464, -22.09384, 
    -21.90241, -21.71037, -21.5177, -21.32441, -21.1305, -20.93596, 
    -20.74079, -20.54499, -20.34856, -20.1515, -19.95382, -19.7555, 
    -19.55654, -19.35695, -19.15673, -18.95588, -18.75438, -18.55226, 
    -18.34949, -18.14609, -17.94205, -17.73737, -17.53205, -17.32609, 
    -17.11949, -16.91226, -16.70438, -16.49586, -16.28671, -16.07691, 
    -15.86647, -15.65539, -15.44367, -15.23131, -15.01831, -14.80467, 
    -14.59039, -14.37547, -14.15991, -13.94372, -13.72688, -13.50941, 
    -13.29131, -13.07256, -12.85318, -12.63317, -12.41252, -12.19124, 
    -11.96933, -11.74679, -11.52362, -11.29982, -11.07539, -10.85034, 
    -10.62466, -10.39836, -10.17144, -9.943896, -9.715737, -9.486961, 
    -9.257571, -9.027569, -8.796955, -8.565732, -8.333903, -8.10147, 
    -7.868433, -7.634798, -7.400565, -7.165736, -6.930315, -6.694304, 
    -6.457705, -6.220523, -5.982759, -5.744415, -5.505497, -5.266005, 
    -5.025944, -4.785316, -4.544127, -4.302377, -4.060071, -3.817212, 
    -3.573805, -3.329853, -3.085359, -2.840328, -2.594763, -2.348668, 
    -2.102048, -1.854907, -1.607249, -1.359079, -1.1104, -0.861218, 
    -0.6115367, -0.3613611, -0.1106959, 0.1404541, 0.3920839, 0.6441885, 
    0.8967628, 1.149802, 1.4033, 1.657252, 1.911653, 2.166498, 2.42178, 
    2.677493, 2.933634, 3.190195, 3.44717, 3.704554, 3.962342, 4.220526, 
    4.4791, 4.738059, 4.997396, 5.257105, 5.517179, 5.777613, 6.038398, 
    6.299529, 6.560999, 6.822802, 7.08493, 7.347377, 7.610135, 7.873198, 
    8.136559, 8.40021, 8.664145, 8.928355, 9.192835, 9.457576, 9.722571, 
    9.987813, 10.25329, 10.51901, 10.78494, 11.0511, 11.31746, 11.58402, 
    11.85078, 12.11772, 12.38484, 12.65214, 12.91959, 13.18719, 13.45495, 
    13.72284, 13.99086, 14.259, 14.52726, 14.79562, 15.06408, 15.33263, 
    15.60127, 15.86997, 16.13874, 16.40757, 16.67645, 16.94537, 17.21432, 
    17.48329, 17.75228, 18.02127, 18.29027, 18.55926, 18.82823, 19.09718, 
    19.36609, 19.63496, 19.90377, 20.17254, 20.44123, 20.70985, 20.97839, 
    21.24683, 21.51518, 21.78342, 22.05155, 22.31955, 22.58742, 22.85515, 
    23.12273, 23.39016, 23.65742, 23.92451, 24.19143, 24.45815, 24.72469, 
    24.99102, 25.25714, 25.52304, 25.78872, 26.05416, 26.31936, 26.58432, 
    26.84902, 27.11346, 27.37762, 27.64151, 27.90512, 28.16843, 28.43145, 
    28.69416, 28.95656, 29.21863, 29.48038, 29.7418, 30.00288, 30.26361, 
    30.52398, 30.784, 31.04365, 31.30293, 31.56183, 31.82034, 32.07846, 
    32.33619, 32.59351, 32.85042, 33.10691, 33.36298, 33.61863, 33.87384, 
    34.12862, 34.38295, 34.63683, 34.89025, 35.14322, 35.39572, 35.64775, 
    35.89931, 36.15038, 36.40097, 36.65107, 36.90067, 37.14977, 37.39837, 
    37.64646, 37.89404, 38.14109, 38.38763, 38.63364, 38.87912, 39.12407, 
    39.36848, 39.61234, 39.85566, 40.09844, 40.34066, 40.58232, 40.82342, 
    41.06396, 41.30393, 41.54333, 41.78215, 42.02041, 42.25808, 42.49517, 
    42.73167, 42.96759, 43.20292, 43.43766, 43.67179, 43.90533, 44.13828, 
    44.37061, 44.60235, 44.83347, 45.06399, 45.2939, 45.52319, 45.75187, 
    45.97993, 46.20737, 46.4342, 46.6604, 46.88598, 47.11093, 47.33526, 
    47.55896, 47.78203, 48.00447, 48.22629, 48.44747, 48.66801, 48.88793, 
    49.1072, 49.32585, 49.54386, 49.76123, 49.97796, 50.19405, 50.40951, 
    50.62433, 50.83851, 51.05205, 51.26495, 51.4772, 51.68882, 51.8998, 
    52.11014, 52.31983, 52.52889, 52.7373, 52.94508, 53.15222, 53.35871, 
    53.56457, 53.76979, 53.97437, 54.17831, 54.38161, 54.58427, 54.7863, 
    54.98769, 55.18845, 55.38857, 55.58805, 55.78691, 55.98513, 56.18272, 
    56.37967, 56.576, 56.7717, 56.96677, 57.16121, 57.35503, 57.54822, 
    57.74079, 57.93274, 58.12406, 58.31476, 58.50485, 58.69431,
  -37.96057, -37.82063, -37.68025, -37.53942, -37.39815, -37.25644, 
    -37.11427, -36.97165, -36.82858, -36.68505, -36.54107, -36.39662, 
    -36.25172, -36.10634, -35.96051, -35.8142, -35.66742, -35.52017, 
    -35.37245, -35.22425, -35.07557, -34.9264, -34.77676, -34.62663, 
    -34.47601, -34.3249, -34.1733, -34.0212, -33.86861, -33.71552, -33.56193, 
    -33.40784, -33.25324, -33.09814, -32.94252, -32.7864, -32.62976, 
    -32.4726, -32.31493, -32.15674, -31.99803, -31.83879, -31.67902, 
    -31.51873, -31.35791, -31.19655, -31.03466, -30.87224, -30.70927, 
    -30.54577, -30.38172, -30.21712, -30.05198, -29.8863, -29.72005, 
    -29.55326, -29.38591, -29.21801, -29.04954, -28.88052, -28.71093, 
    -28.54077, -28.37005, -28.19876, -28.0269, -27.85446, -27.68145, 
    -27.50787, -27.3337, -27.15896, -26.98363, -26.80772, -26.63122, 
    -26.45414, -26.27646, -26.09819, -25.91933, -25.73988, -25.55983, 
    -25.37918, -25.19793, -25.01608, -24.83362, -24.65056, -24.4669, 
    -24.28262, -24.09774, -23.91224, -23.72614, -23.53942, -23.35208, 
    -23.16412, -22.97555, -22.78635, -22.59654, -22.4061, -22.21504, 
    -22.02335, -21.83104, -21.6381, -21.44453, -21.25033, -21.0555, 
    -20.86004, -20.66394, -20.46721, -20.26985, -20.07185, -19.87321, 
    -19.67393, -19.47402, -19.27346, -19.07227, -18.87043, -18.66796, 
    -18.46484, -18.26107, -18.05667, -17.85162, -17.64593, -17.43959, 
    -17.2326, -17.02498, -16.8167, -16.60778, -16.39822, -16.18801, 
    -15.97715, -15.76564, -15.55349, -15.3407, -15.12725, -14.91317, 
    -14.69843, -14.48305, -14.26703, -14.05036, -13.83305, -13.6151, 
    -13.3965, -13.17726, -12.95738, -12.73686, -12.5157, -12.2939, -12.07146, 
    -11.84839, -11.62468, -11.40033, -11.17535, -10.94975, -10.72351, 
    -10.49664, -10.26914, -10.04102, -9.812269, -9.582899, -9.352909, 
    -9.122299, -8.891072, -8.659231, -8.426776, -8.19371, -7.960036, 
    -7.725756, -7.490872, -7.255386, -7.019301, -6.78262, -6.545346, 
    -6.307481, -6.069028, -5.829989, -5.590369, -5.35017, -5.109395, 
    -4.868048, -4.626131, -4.383648, -4.140604, -3.897, -3.652842, -3.408132, 
    -3.162874, -2.917073, -2.670732, -2.423856, -2.176448, -1.928513, 
    -1.680055, -1.431079, -1.181589, -0.9315885, -0.6810836, -0.4300786, 
    -0.1785782, 0.07341266, 0.3258891, 0.5788459, 0.8322782, 1.086181, 
    1.340548, 1.595375, 1.850656, 2.106385, 2.362557, 2.619167, 2.876209, 
    3.133676, 3.391562, 3.649863, 3.908571, 4.167682, 4.427187, 4.687082, 
    4.94736, 5.208014, 5.469038, 5.730425, 5.992169, 6.254263, 6.516701, 
    6.779475, 7.042579, 7.306005, 7.569747, 7.833797, 8.098149, 8.362796, 
    8.627728, 8.892941, 9.158427, 9.424177, 9.690185, 9.956442, 10.22294, 
    10.48968, 10.75664, 11.02382, 11.29121, 11.55881, 11.8266, 12.09458, 
    12.36274, 12.63107, 12.89957, 13.16822, 13.43702, 13.70596, 13.97504, 
    14.24423, 14.51355, 14.78296, 15.05248, 15.32209, 15.59178, 15.86155, 
    16.13138, 16.40127, 16.67121, 16.94119, 17.21121, 17.48125, 17.7513, 
    18.02136, 18.29142, 18.56147, 18.83151, 19.10151, 19.37149, 19.64142, 
    19.9113, 20.18113, 20.45088, 20.72056, 20.99016, 21.25966, 21.52906, 
    21.79836, 22.06753, 22.33659, 22.6055, 22.87428, 23.14291, 23.41138, 
    23.67969, 23.94782, 24.21577, 24.48353, 24.7511, 25.01846, 25.28561, 
    25.55253, 25.81923, 26.08569, 26.35191, 26.61788, 26.88359, 27.14903, 
    27.4142, 27.67909, 27.94369, 28.20799, 28.47199, 28.73569, 28.99906, 
    29.26211, 29.52484, 29.78722, 30.04926, 30.31095, 30.57228, 30.83324, 
    31.09384, 31.35406, 31.61389, 31.87333, 32.13238, 32.39102, 32.64926, 
    32.90708, 33.16448, 33.42145, 33.67799, 33.9341, 34.18975, 34.44497, 
    34.69972, 34.95401, 35.20784, 35.4612, 35.71408, 35.96648, 36.2184, 
    36.46982, 36.72074, 36.97117, 37.22109, 37.4705, 37.71939, 37.96777, 
    38.21562, 38.46294, 38.70974, 38.95599, 39.20171, 39.44688, 39.6915, 
    39.93557, 40.17908, 40.42204, 40.66444, 40.90626, 41.14752, 41.3882, 
    41.62831, 41.86784, 42.10678, 42.34515, 42.58292, 42.8201, 43.05669, 
    43.29268, 43.52806, 43.76286, 43.99704, 44.23062, 44.46359, 44.69595, 
    44.92769, 45.15882, 45.38933, 45.61922, 45.8485, 46.07714, 46.30517, 
    46.53257, 46.75933, 46.98547, 47.21098, 47.43586, 47.66011, 47.88372, 
    48.10669, 48.32903, 48.55072, 48.77178, 48.9922, 49.21198, 49.43112, 
    49.64962, 49.86747, 50.08468, 50.30125, 50.51717, 50.73244, 50.94707, 
    51.16106, 51.3744, 51.58709, 51.79914, 52.01054, 52.2213, 52.43141, 
    52.64087, 52.84969, 53.05787, 53.26539, 53.47227, 53.67851, 53.8841, 
    54.08905, 54.29335, 54.49701, 54.70003, 54.9024, 55.10414, 55.30523, 
    55.50568, 55.7055, 55.90467, 56.10321, 56.30111, 56.49837, 56.695, 
    56.891, 57.08636, 57.28109, 57.47519, 57.66866, 57.8615, 58.05372, 
    58.2453, 58.43627, 58.62661, 58.81632,
  -38.09159, -37.95167, -37.81131, -37.6705, -37.52925, -37.38755, -37.24539, 
    -37.10279, -36.95973, -36.81621, -36.67223, -36.52779, -36.38288, 
    -36.23751, -36.09167, -35.94537, -35.79859, -35.65133, -35.5036, 
    -35.35538, -35.20669, -35.05751, -34.90785, -34.75771, -34.60706, 
    -34.45593, -34.30431, -34.15218, -33.99957, -33.84644, -33.69282, 
    -33.53869, -33.38405, -33.2289, -33.07325, -32.91708, -32.76039, 
    -32.60318, -32.44546, -32.28721, -32.12844, -31.96914, -31.80931, 
    -31.64895, -31.48806, -31.32663, -31.16467, -31.00216, -30.83912, 
    -30.67553, -30.5114, -30.34671, -30.18148, -30.0157, -29.84936, 
    -29.68246, -29.51501, -29.34699, -29.17842, -29.00928, -28.83957, 
    -28.6693, -28.49845, -28.32703, -28.15504, -27.98247, -27.80933, 
    -27.6356, -27.46129, -27.2864, -27.11092, -26.93485, -26.75819, 
    -26.58094, -26.4031, -26.22467, -26.04563, -25.866, -25.68577, -25.50493, 
    -25.32349, -25.14145, -24.95879, -24.77553, -24.59166, -24.40718, 
    -24.22208, -24.03636, -23.85003, -23.66308, -23.47551, -23.28732, 
    -23.09851, -22.90907, -22.719, -22.52831, -22.33699, -22.14504, 
    -21.95246, -21.75925, -21.5654, -21.37092, -21.1758, -20.98005, 
    -20.78365, -20.58662, -20.38895, -20.19064, -19.99168, -19.79208, 
    -19.59184, -19.39095, -19.18942, -18.98724, -18.78442, -18.58094, 
    -18.37682, -18.17205, -17.96664, -17.76057, -17.55385, -17.34648, 
    -17.13846, -16.92979, -16.72047, -16.51049, -16.29987, -16.08859, 
    -15.87666, -15.66408, -15.45084, -15.23696, -15.02242, -14.80723, 
    -14.5914, -14.37491, -14.15777, -13.93998, -13.72154, -13.50245, 
    -13.28271, -13.06233, -12.8413, -12.61962, -12.3973, -12.17434, 
    -11.95073, -11.72648, -11.50159, -11.27606, -11.04989, -10.82309, 
    -10.59565, -10.36757, -10.13887, -9.909531, -9.679564, -9.448971, 
    -9.217752, -8.98591, -8.753447, -8.520364, -8.286663, -8.052348, 
    -7.81742, -7.581882, -7.345736, -7.108985, -6.871631, -6.633677, 
    -6.395125, -6.15598, -5.916243, -5.675918, -5.435007, -5.193514, 
    -4.951442, -4.708795, -4.465576, -4.221788, -3.977435, -3.73252, 
    -3.487048, -3.241023, -2.994447, -2.747326, -2.499663, -2.251462, 
    -2.002728, -1.753465, -1.503677, -1.253369, -1.002546, -0.7512121, 
    -0.499372, -0.2470307, 0.005806944, 0.2591359, 0.5129511, 0.7672474, 
    1.022019, 1.277262, 1.53297, 1.789137, 2.045758, 2.302828, 2.56034, 
    2.818289, 3.076669, 3.335474, 3.594699, 3.854336, 4.114379, 4.374823, 
    4.635661, 4.896886, 5.158494, 5.420475, 5.682824, 5.945535, 6.2086, 
    6.472013, 6.735766, 6.999854, 7.264267, 7.529001, 7.794048, 8.0594, 
    8.325049, 8.590989, 8.857213, 9.123713, 9.39048, 9.657509, 9.92479, 
    10.19232, 10.46008, 10.72808, 10.99629, 11.26473, 11.53336, 11.8022, 
    12.07123, 12.34044, 12.60982, 12.87937, 13.14908, 13.41894, 13.68894, 
    13.95907, 14.22933, 14.49971, 14.77019, 15.04078, 15.31145, 15.58222, 
    15.85305, 16.12395, 16.39492, 16.66593, 16.93698, 17.20807, 17.47918, 
    17.75031, 18.02144, 18.29258, 18.56371, 18.83481, 19.1059, 19.37694, 
    19.64795, 19.9189, 20.18979, 20.46062, 20.73137, 21.00203, 21.2726, 
    21.54307, 21.81343, 22.08367, 22.35378, 22.62376, 22.89359, 23.16328, 
    23.4328, 23.70216, 23.97134, 24.24034, 24.50914, 24.77775, 25.04615, 
    25.31433, 25.58229, 25.85002, 26.11751, 26.38475, 26.65174, 26.91846, 
    27.18492, 27.4511, 27.71699, 27.9826, 28.2479, 28.5129, 28.77758, 
    29.04194, 29.30598, 29.56968, 29.83304, 30.09604, 30.3587, 30.62099, 
    30.88291, 31.14446, 31.40562, 31.6664, 31.92678, 32.18676, 32.44633, 
    32.70549, 32.96423, 33.22254, 33.48042, 33.73787, 33.99487, 34.25142, 
    34.50751, 34.76315, 35.01831, 35.27301, 35.52723, 35.78097, 36.03422, 
    36.28698, 36.53924, 36.791, 37.04226, 37.293, 37.54322, 37.79293, 
    38.04211, 38.29076, 38.53888, 38.78645, 39.03349, 39.27998, 39.52591, 
    39.7713, 40.01612, 40.26039, 40.50409, 40.74722, 40.98977, 41.23175, 
    41.47315, 41.71397, 41.9542, 42.19385, 42.4329, 42.67136, 42.90922, 
    43.14648, 43.38313, 43.61918, 43.85462, 44.08945, 44.32367, 44.55727, 
    44.79026, 45.02262, 45.25437, 45.48549, 45.71598, 45.94585, 46.17509, 
    46.40369, 46.63167, 46.85901, 47.08571, 47.31178, 47.53721, 47.762, 
    47.98615, 48.20965, 48.43251, 48.65473, 48.8763, 49.09723, 49.31751, 
    49.53715, 49.75613, 49.97447, 50.19216, 50.40919, 50.62558, 50.84132, 
    51.0564, 51.27084, 51.48462, 51.69775, 51.91022, 52.12205, 52.33323, 
    52.54375, 52.75362, 52.96284, 53.17141, 53.37933, 53.58659, 53.79321, 
    53.99917, 54.20449, 54.40916, 54.61317, 54.81654, 55.01927, 55.22134, 
    55.42277, 55.62356, 55.8237, 56.02319, 56.22205, 56.42026, 56.61783, 
    56.81476, 57.01105, 57.20671, 57.40172, 57.5961, 57.78985, 57.98296, 
    58.17545, 58.3673, 58.55852, 58.74911, 58.93908,
  -38.22316, -38.08326, -37.94292, -37.80214, -37.6609, -37.51922, -37.37708, 
    -37.23449, -37.09144, -36.94794, -36.80397, -36.65953, -36.51463, 
    -36.36927, -36.22343, -36.07712, -35.93034, -35.78308, -35.63534, 
    -35.48712, -35.33842, -35.18923, -35.03955, -34.88939, -34.73873, 
    -34.58758, -34.43593, -34.28378, -34.13113, -33.97798, -33.82433, 
    -33.67016, -33.51549, -33.36031, -33.20461, -33.04839, -32.89166, 
    -32.7344, -32.57663, -32.41832, -32.25949, -32.10014, -31.94025, 
    -31.77983, -31.61887, -31.45737, -31.29533, -31.13275, -30.96963, 
    -30.80596, -30.64174, -30.47697, -30.31165, -30.14577, -29.97934, 
    -29.81234, -29.64478, -29.47667, -29.30798, -29.13873, -28.96891, 
    -28.79851, -28.62755, -28.456, -28.28388, -28.11118, -27.9379, -27.76403, 
    -27.58958, -27.41454, -27.23891, -27.06269, -26.88588, -26.70847, 
    -26.53046, -26.35186, -26.17265, -25.99284, -25.81243, -25.63141, 
    -25.44978, -25.26755, -25.0847, -24.90123, -24.71716, -24.53246, 
    -24.34715, -24.16122, -23.97467, -23.78749, -23.59969, -23.41127, 
    -23.22221, -23.03253, -22.84222, -22.65127, -22.45969, -22.26748, 
    -22.07463, -21.88115, -21.68703, -21.49226, -21.29686, -21.10081, 
    -20.90412, -20.70679, -20.50881, -20.31019, -20.11092, -19.911, 
    -19.71043, -19.50921, -19.30734, -19.10482, -18.90165, -18.69782, 
    -18.49334, -18.28821, -18.08242, -17.87598, -17.66888, -17.46113, 
    -17.25271, -17.04365, -16.83392, -16.62354, -16.4125, -16.2008, 
    -15.98845, -15.77543, -15.56176, -15.34743, -15.13245, -14.9168, 
    -14.7005, -14.48355, -14.26593, -14.04766, -13.82874, -13.60916, 
    -13.38893, -13.16804, -12.9465, -12.72431, -12.50147, -12.27797, 
    -12.05383, -11.82904, -11.6036, -11.37752, -11.15079, -10.92342, 
    -10.69541, -10.46675, -10.23746, -10.00753, -9.776965, -9.545767, 
    -9.313936, -9.081476, -8.848389, -8.614675, -8.380337, -8.145377, 
    -7.909799, -7.673604, -7.436794, -7.199373, -6.961343, -6.722706, 
    -6.483465, -6.243624, -6.003184, -5.76215, -5.520524, -5.278309, 
    -5.035509, -4.792127, -4.548167, -4.303631, -4.058524, -3.81285, 
    -3.566611, -3.319813, -3.072458, -2.824551, -2.576096, -2.327097, 
    -2.077559, -1.827485, -1.576881, -1.325751, -1.074099, -0.8219298, 
    -0.569249, -0.3160609, -0.06237053, 0.191817, 0.4464966, 0.701663, 
    0.9573111, 1.213435, 1.47003, 1.72709, 1.98461, 2.242584, 2.501005, 
    2.759869, 3.01917, 3.2789, 3.539055, 3.799627, 4.060612, 4.322001, 
    4.58379, 4.845971, 5.108538, 5.371485, 5.634804, 5.898489, 6.162533, 
    6.426929, 6.69167, 6.956749, 7.222159, 7.487894, 7.753944, 8.020304, 
    8.286965, 8.553922, 8.821164, 9.088687, 9.356482, 9.624539, 9.892855, 
    10.16142, 10.43022, 10.69926, 10.96852, 11.238, 11.50769, 11.77758, 
    12.04766, 12.31793, 12.58838, 12.85899, 13.12976, 13.40069, 13.67176, 
    13.94296, 14.21429, 14.48574, 14.7573, 15.02896, 15.30072, 15.57256, 
    15.84448, 16.11646, 16.3885, 16.6606, 16.93273, 17.2049, 17.4771, 
    17.74931, 18.02153, 18.29375, 18.56596, 18.83815, 19.11032, 19.38245, 
    19.65453, 19.92657, 20.19854, 20.47045, 20.74227, 21.01402, 21.28566, 
    21.55721, 21.82864, 22.09995, 22.37113, 22.64218, 22.91308, 23.18383, 
    23.45442, 23.72483, 23.99507, 24.26513, 24.53498, 24.80464, 25.07409, 
    25.34331, 25.61231, 25.88108, 26.1496, 26.41788, 26.6859, 26.95365, 
    27.22113, 27.48833, 27.75524, 28.02185, 28.28816, 28.55416, 28.81985, 
    29.0852, 29.35023, 29.61492, 29.87926, 30.14325, 30.40687, 30.67013, 
    30.93302, 31.19553, 31.45765, 31.71937, 31.9807, 32.24162, 32.50212, 
    32.76221, 33.02188, 33.28111, 33.5399, 33.79825, 34.05616, 34.3136, 
    34.57059, 34.82711, 35.08316, 35.33873, 35.59382, 35.84842, 36.10253, 
    36.35614, 36.60925, 36.86185, 37.11394, 37.36551, 37.61656, 37.86708, 
    38.11707, 38.36652, 38.61543, 38.8638, 39.11162, 39.35889, 39.6056, 
    39.85175, 40.09734, 40.34235, 40.5868, 40.83067, 41.07396, 41.31666, 
    41.55878, 41.80032, 42.04126, 42.2816, 42.52135, 42.76049, 42.99903, 
    43.23697, 43.47429, 43.71101, 43.94711, 44.18259, 44.41745, 44.65168, 
    44.8853, 45.11829, 45.35065, 45.58238, 45.81348, 46.04395, 46.27377, 
    46.50296, 46.73151, 46.95943, 47.1867, 47.41332, 47.63931, 47.86464, 
    48.08933, 48.31337, 48.53676, 48.7595, 48.98159, 49.20303, 49.42381, 
    49.64394, 49.86341, 50.08223, 50.3004, 50.51791, 50.73476, 50.95096, 
    51.1665, 51.38138, 51.5956, 51.80917, 52.02208, 52.23433, 52.44593, 
    52.65686, 52.86714, 53.07676, 53.28572, 53.49403, 53.70168, 53.90868, 
    54.11502, 54.3207, 54.52573, 54.73011, 54.93383, 55.1369, 55.33932, 
    55.54108, 55.7422, 55.94267, 56.14248, 56.34165, 56.54017, 56.73805, 
    56.93528, 57.13187, 57.32781, 57.52311, 57.71777, 57.9118, 58.10518, 
    58.29793, 58.49004, 58.68152, 58.87236, 59.06258,
  -38.35528, -38.21541, -38.0751, -37.93434, -37.79313, -37.65146, -37.50934, 
    -37.36677, -37.22374, -37.08024, -36.93628, -36.79186, -36.64697, 
    -36.50161, -36.35577, -36.20947, -36.06269, -35.91542, -35.76768, 
    -35.61946, -35.47075, -35.32155, -35.17186, -35.02168, -34.87101, 
    -34.71983, -34.56816, -34.416, -34.26332, -34.11015, -33.95646, 
    -33.80227, -33.64756, -33.49234, -33.3366, -33.18034, -33.02357, 
    -32.86626, -32.70844, -32.55009, -32.3912, -32.23179, -32.07184, 
    -31.91136, -31.75033, -31.58877, -31.42666, -31.26401, -31.10081, 
    -30.93706, -30.77276, -30.6079, -30.44249, -30.27653, -30.11, -29.94291, 
    -29.77525, -29.60703, -29.43824, -29.26887, -29.09894, -28.92843, 
    -28.75734, -28.58568, -28.41343, -28.2406, -28.06718, -27.89318, 
    -27.71859, -27.5434, -27.36763, -27.19125, -27.01429, -26.83672, 
    -26.65855, -26.47978, -26.3004, -26.12042, -25.93983, -25.75862, 
    -25.57681, -25.39438, -25.21134, -25.02768, -24.8434, -24.65849, 
    -24.47297, -24.28683, -24.10005, -23.91265, -23.72462, -23.53596, 
    -23.34667, -23.15675, -22.96619, -22.77499, -22.58316, -22.39068, 
    -22.19757, -22.00381, -21.80942, -21.61437, -21.41868, -21.22235, 
    -21.02536, -20.82773, -20.62945, -20.43051, -20.23092, -20.03069, 
    -19.82979, -19.62824, -19.42604, -19.22318, -19.01966, -18.81548, 
    -18.61064, -18.40514, -18.19899, -17.99217, -17.78469, -17.57655, 
    -17.36775, -17.15828, -16.94815, -16.73736, -16.52591, -16.31379, 
    -16.10101, -15.88757, -15.67346, -15.45868, -15.24325, -15.02715, 
    -14.81039, -14.59296, -14.37488, -14.15613, -13.93672, -13.71665, 
    -13.49591, -13.27452, -13.05247, -12.82976, -12.60639, -12.38237, 
    -12.15769, -11.93236, -11.70637, -11.47973, -11.25244, -11.0245, 
    -10.79591, -10.56668, -10.3368, -10.10628, -9.875111, -9.643305, 
    -9.41086, -9.177779, -8.944064, -8.709717, -8.474739, -8.239133, 
    -8.002901, -7.766046, -7.52857, -7.290475, -7.051765, -6.812442, 
    -6.572508, -6.331967, -6.090822, -5.849075, -5.60673, -5.363789, 
    -5.120256, -4.876136, -4.63143, -4.386143, -4.140277, -3.893838, 
    -3.646828, -3.399252, -3.151113, -2.902416, -2.653164, -2.403362, 
    -2.153014, -1.902125, -1.650699, -1.39874, -1.146254, -0.8932445, 
    -0.639717, -0.3856763, -0.1311274, 0.1239248, 0.3794749, 0.6355178, 
    0.8920482, 1.14906, 1.406549, 1.664509, 1.922934, 2.181818, 2.441156, 
    2.700942, 2.961169, 3.221832, 3.482924, 3.74444, 4.006372, 4.268716, 
    4.531463, 4.794607, 5.058143, 5.322062, 5.586359, 5.851026, 6.116057, 
    6.381444, 6.647182, 6.913261, 7.179676, 7.446418, 7.713481, 7.980858, 
    8.24854, 8.516521, 8.784792, 9.053346, 9.322175, 9.591272, 9.86063, 
    10.13024, 10.40009, 10.67018, 10.9405, 11.21103, 11.48178, 11.75274, 
    12.02388, 12.29522, 12.56674, 12.83842, 13.11027, 13.38227, 13.65442, 
    13.9267, 14.19912, 14.47165, 14.74429, 15.01704, 15.28989, 15.56281, 
    15.83582, 16.1089, 16.38203, 16.65522, 16.92845, 17.20171, 17.475, 
    17.7483, 18.02162, 18.29493, 18.56823, 18.84152, 19.11478, 19.388, 
    19.66118, 19.9343, 20.20737, 20.48036, 20.75328, 21.02611, 21.29884, 
    21.57147, 21.84398, 22.11638, 22.38864, 22.66077, 22.93274, 23.20457, 
    23.47622, 23.74771, 24.01902, 24.29014, 24.56106, 24.83177, 25.10228, 
    25.37256, 25.64261, 25.91243, 26.182, 26.45131, 26.72037, 26.98915, 
    27.25766, 27.52589, 27.79382, 28.06146, 28.32878, 28.5958, 28.86249, 
    29.12885, 29.39488, 29.66056, 29.92589, 30.19086, 30.45547, 30.71971, 
    30.98357, 31.24704, 31.51013, 31.77281, 32.03509, 32.29696, 32.5584, 
    32.81943, 33.08002, 33.34018, 33.5999, 33.85917, 34.11798, 34.37633, 
    34.63421, 34.89163, 35.14856, 35.40502, 35.66098, 35.91645, 36.17142, 
    36.4259, 36.67986, 36.9333, 37.18623, 37.43863, 37.69051, 37.94185, 
    38.19265, 38.44291, 38.69263, 38.94179, 39.1904, 39.43845, 39.68594, 
    39.93286, 40.17921, 40.42498, 40.67018, 40.91479, 41.15882, 41.40226, 
    41.6451, 41.88736, 42.12901, 42.37006, 42.6105, 42.85034, 43.08957, 
    43.32818, 43.56618, 43.80355, 44.04031, 44.27644, 44.51195, 44.74683, 
    44.98108, 45.21469, 45.44767, 45.68002, 45.91172, 46.14278, 46.37321, 
    46.60299, 46.83212, 47.0606, 47.28844, 47.51562, 47.74216, 47.96805, 
    48.19328, 48.41785, 48.64177, 48.86503, 49.08764, 49.30959, 49.53087, 
    49.7515, 49.97147, 50.19077, 50.40942, 50.6274, 50.84472, 51.06138, 
    51.27737, 51.4927, 51.70737, 51.92137, 52.13471, 52.34739, 52.5594, 
    52.77075, 52.98144, 53.19146, 53.40082, 53.60952, 53.81755, 54.02493, 
    54.23164, 54.43769, 54.64309, 54.84782, 55.05189, 55.25531, 55.45807, 
    55.66017, 55.86161, 56.0624, 56.26254, 56.46202, 56.66085, 56.85904, 
    57.05656, 57.25345, 57.44968, 57.64527, 57.84021, 58.03451, 58.22816, 
    58.42117, 58.61354, 58.80528, 58.99637, 59.18683,
  -38.48796, -38.34813, -38.20784, -38.0671, -37.92591, -37.78427, -37.64217, 
    -37.49962, -37.3566, -37.21312, -37.06918, -36.92477, -36.77989, 
    -36.63454, -36.48871, -36.34241, -36.19563, -36.04837, -35.90062, 
    -35.7524, -35.60368, -35.45447, -35.30478, -35.15459, -35.0039, 
    -34.85271, -34.70102, -34.54884, -34.39614, -34.24294, -34.08923, 
    -33.935, -33.78026, -33.62501, -33.46923, -33.31294, -33.15612, 
    -32.99878, -32.8409, -32.6825, -32.52357, -32.3641, -32.20409, -32.04355, 
    -31.88246, -31.72083, -31.55866, -31.39593, -31.23266, -31.06883, 
    -30.90445, -30.73952, -30.57402, -30.40796, -30.24134, -30.07416, 
    -29.9064, -29.73808, -29.56919, -29.39972, -29.22967, -29.05905, 
    -28.88784, -28.71605, -28.54368, -28.37072, -28.19718, -28.02304, 
    -27.84831, -27.67298, -27.49706, -27.32054, -27.14342, -26.96569, 
    -26.78736, -26.60843, -26.42888, -26.24872, -26.06796, -25.88657, 
    -25.70457, -25.52196, -25.33872, -25.15486, -24.97038, -24.78528, 
    -24.59954, -24.41318, -24.22619, -24.03857, -23.85031, -23.66142, 
    -23.47189, -23.28173, -23.09092, -22.89948, -22.70739, -22.51465, 
    -22.32128, -22.12725, -21.93258, -21.73726, -21.54128, -21.34466, 
    -21.14738, -20.94945, -20.75086, -20.55161, -20.35172, -20.15116, 
    -19.94994, -19.74806, -19.54552, -19.34231, -19.13844, -18.93392, 
    -18.72872, -18.52286, -18.31634, -18.10915, -17.90129, -17.69276, 
    -17.48357, -17.27371, -17.06318, -16.85198, -16.64011, -16.42757, 
    -16.21436, -16.00049, -15.78594, -15.57072, -15.35484, -15.13828, 
    -14.92106, -14.70317, -14.4846, -14.26537, -14.04548, -13.82491, 
    -13.60368, -13.38178, -13.15922, -12.93599, -12.7121, -12.48754, 
    -12.26233, -12.03645, -11.80991, -11.58272, -11.35486, -11.12635, 
    -10.89719, -10.66737, -10.4369, -10.20578, -9.974009, -9.741593, 
    -9.508533, -9.274829, -9.040483, -8.8055, -8.569879, -8.333623, 
    -8.096735, -7.859217, -7.621071, -7.3823, -7.142907, -6.902894, 
    -6.662263, -6.421019, -6.179164, -5.9367, -5.693632, -5.449962, 
    -5.205693, -4.960829, -4.715374, -4.46933, -4.222702, -3.975493, 
    -3.727708, -3.479349, -3.230421, -2.980928, -2.730875, -2.480264, 
    -2.229102, -1.977392, -1.725138, -1.472346, -1.21902, -0.9651641, 
    -0.7107842, -0.4558849, -0.2004713, 0.05545162, 0.3118786, 0.5688042, 
    0.8262233, 1.08413, 1.342519, 1.601385, 1.860722, 2.120524, 2.380785, 
    2.6415, 2.902661, 3.164264, 3.426302, 3.688768, 3.951656, 4.21496, 
    4.478673, 4.742788, 5.007299, 5.2722, 5.537482, 5.80314, 6.069166, 
    6.335553, 6.602294, 6.869382, 7.13681, 7.40457, 7.672654, 7.941056, 
    8.209767, 8.478782, 8.74809, 9.017685, 9.287559, 9.557704, 9.828113, 
    10.09878, 10.36969, 10.64084, 10.91222, 11.18382, 11.45564, 11.72766, 
    11.99989, 12.2723, 12.5449, 12.81766, 13.0906, 13.36368, 13.63692, 
    13.91029, 14.1838, 14.45743, 14.73117, 15.00501, 15.27895, 15.55298, 
    15.82709, 16.10126, 16.3755, 16.64979, 16.92412, 17.19849, 17.47288, 
    17.74729, 18.0217, 18.29612, 18.57053, 18.84492, 19.11928, 19.3936, 
    19.66788, 19.94211, 20.21628, 20.49037, 20.76439, 21.03831, 21.31214, 
    21.58586, 21.85947, 22.13296, 22.40631, 22.67952, 22.95259, 23.22549, 
    23.49824, 23.7708, 24.04319, 24.31538, 24.58737, 24.85916, 25.13073, 
    25.40207, 25.67318, 25.94406, 26.21468, 26.48505, 26.75515, 27.02498, 
    27.29453, 27.56379, 27.83276, 28.10142, 28.36977, 28.63781, 28.90552, 
    29.17289, 29.43992, 29.70661, 29.97294, 30.23891, 30.50451, 30.76973, 
    31.03457, 31.29902, 31.56307, 31.82672, 32.08996, 32.35278, 32.61518, 
    32.87715, 33.13868, 33.39977, 33.66042, 33.9206, 34.18033, 34.43959, 
    34.69839, 34.9567, 35.21453, 35.47187, 35.72872, 35.98507, 36.24091, 
    36.49624, 36.75106, 37.00536, 37.25913, 37.51237, 37.76508, 38.01724, 
    38.26887, 38.51994, 38.77047, 39.02043, 39.26984, 39.51867, 39.76694, 
    40.01464, 40.26175, 40.50829, 40.75424, 40.9996, 41.24437, 41.48855, 
    41.73212, 41.97509, 42.21746, 42.45922, 42.70037, 42.9409, 43.18082, 
    43.42011, 43.65878, 43.89683, 44.13425, 44.37104, 44.60719, 44.84271, 
    45.07759, 45.31184, 45.54544, 45.7784, 46.01072, 46.24238, 46.4734, 
    46.70377, 46.93348, 47.16254, 47.39095, 47.6187, 47.84579, 48.07222, 
    48.298, 48.52311, 48.74756, 48.97134, 49.19447, 49.41693, 49.63872, 
    49.85984, 50.0803, 50.30009, 50.51922, 50.73767, 50.95546, 51.17258, 
    51.38903, 51.60481, 51.81992, 52.03436, 52.24813, 52.46124, 52.67367, 
    52.88543, 53.09652, 53.30695, 53.5167, 53.72579, 53.93421, 54.14196, 
    54.34905, 54.55547, 54.76122, 54.96631, 55.17074, 55.3745, 55.5776, 
    55.78003, 55.98181, 56.18292, 56.38338, 56.58318, 56.78232, 56.9808, 
    57.17863, 57.3758, 57.57232, 57.7682, 57.96341, 58.15799, 58.35191, 
    58.54519, 58.73782, 58.9298, 59.12115, 59.31185,
  -38.62121, -38.4814, -38.34114, -38.20044, -38.05927, -37.91766, -37.77559, 
    -37.63305, -37.49005, -37.34659, -37.20266, -37.05827, -36.9134, 
    -36.76806, -36.62224, -36.47594, -36.32917, -36.18191, -36.03417, 
    -35.88594, -35.73722, -35.58801, -35.43831, -35.28811, -35.13741, 
    -34.98621, -34.83451, -34.6823, -34.52959, -34.37636, -34.22263, 
    -34.06837, -33.9136, -33.75832, -33.60251, -33.44618, -33.28932, 
    -33.13194, -32.97402, -32.81557, -32.65659, -32.49707, -32.33701, 
    -32.1764, -32.01526, -31.85357, -31.69133, -31.52853, -31.36519, 
    -31.20129, -31.03683, -30.87181, -30.70624, -30.54009, -30.37338, 
    -30.2061, -30.03826, -29.86983, -29.70084, -29.53126, -29.36111, 
    -29.19037, -29.01905, -28.84715, -28.67465, -28.50157, -28.32789, 
    -28.15362, -27.97875, -27.80329, -27.62722, -27.45055, -27.27328, 
    -27.0954, -26.91691, -26.73781, -26.5581, -26.37777, -26.19683, 
    -26.01527, -25.83309, -25.65029, -25.46686, -25.2828, -25.09812, 
    -24.91282, -24.72687, -24.5403, -24.35309, -24.16525, -23.97677, 
    -23.78764, -23.59788, -23.40748, -23.21643, -23.02473, -22.83239, 
    -22.6394, -22.44576, -22.25146, -22.05652, -21.86092, -21.66466, 
    -21.46775, -21.27018, -21.07195, -20.87306, -20.67351, -20.47329, 
    -20.27241, -20.07087, -19.86866, -19.66578, -19.46224, -19.25803, 
    -19.05315, -18.8476, -18.64137, -18.43448, -18.22692, -18.01868, 
    -17.80977, -17.60018, -17.38993, -17.17899, -16.96738, -16.7551, 
    -16.54214, -16.32851, -16.1142, -15.89922, -15.68355, -15.46722, 
    -15.25021, -15.03252, -14.81416, -14.59512, -14.37541, -14.15502, 
    -13.93396, -13.71223, -13.48983, -13.26675, -13.043, -12.81859, -12.5935, 
    -12.36774, -12.14132, -11.91423, -11.68647, -11.45805, -11.22897, 
    -10.99923, -10.76882, -10.53776, -10.30604, -10.07367, -9.840641, 
    -9.606961, -9.372632, -9.137655, -8.902032, -8.665765, -8.428857, 
    -8.191309, -7.953125, -7.714306, -7.474856, -7.234776, -6.99407, 
    -6.752739, -6.510789, -6.26822, -6.025036, -5.781241, -5.536837, 
    -5.291828, -5.046216, -4.800007, -4.553203, -4.305808, -4.057825, 
    -3.809258, -3.560112, -3.31039, -3.060097, -2.809237, -2.557813, 
    -2.305831, -2.053294, -1.800207, -1.546576, -1.292404, -1.037696, 
    -0.7824584, -0.5266945, -0.2704102, -0.01361032, 0.2436997, 0.5015145, 
    0.7598287, 1.018637, 1.277933, 1.537712, 1.797968, 2.058694, 2.319885, 
    2.581536, 2.843639, 3.106189, 3.369179, 3.632603, 3.896455, 4.160727, 
    4.425414, 4.690508, 4.956003, 5.221893, 5.488169, 5.754825, 6.021854, 
    6.28925, 6.557003, 6.825109, 7.093558, 7.362343, 7.631458, 7.900894, 
    8.170644, 8.4407, 8.711055, 8.981699, 9.252626, 9.523829, 9.795298, 
    10.06703, 10.339, 10.61122, 10.88368, 11.15636, 11.42926, 11.70236, 
    11.97567, 12.24917, 12.52286, 12.79672, 13.07074, 13.34493, 13.61926, 
    13.89374, 14.16834, 14.44307, 14.71792, 14.99287, 15.26792, 15.54305, 
    15.81827, 16.09356, 16.36891, 16.64431, 16.91975, 17.19523, 17.47074, 
    17.74626, 18.02179, 18.29732, 18.57284, 18.84835, 19.12382, 19.39926, 
    19.67465, 19.94999, 20.22527, 20.50047, 20.7756, 21.05063, 21.32556, 
    21.60039, 21.8751, 22.14969, 22.42414, 22.69845, 22.97261, 23.24661, 
    23.52045, 23.7941, 24.06757, 24.34085, 24.61393, 24.88679, 25.15944, 
    25.43185, 25.70403, 25.97598, 26.24766, 26.51909, 26.79025, 27.06113, 
    27.33173, 27.60204, 27.87205, 28.14175, 28.41113, 28.6802, 28.94893, 
    29.21732, 29.48537, 29.75307, 30.02041, 30.28738, 30.55398, 30.82019, 
    31.08602, 31.35145, 31.61648, 31.8811, 32.14531, 32.4091, 32.67245, 
    32.93537, 33.19785, 33.45988, 33.72146, 33.98258, 34.24323, 34.50341, 
    34.76311, 35.02234, 35.28107, 35.5393, 35.79704, 36.05426, 36.31099, 
    36.56719, 36.82287, 37.07802, 37.33265, 37.58673, 37.84028, 38.09328, 
    38.34573, 38.59762, 38.84896, 39.09973, 39.34993, 39.59956, 39.84862, 
    40.09709, 40.34498, 40.59228, 40.83899, 41.08511, 41.33062, 41.57554, 
    41.81985, 42.06355, 42.30663, 42.5491, 42.79095, 43.03219, 43.27279, 
    43.51278, 43.75212, 43.99084, 44.22893, 44.46637, 44.70318, 44.93935, 
    45.17487, 45.40974, 45.64397, 45.87754, 46.11047, 46.34274, 46.57436, 
    46.80531, 47.03561, 47.26525, 47.49423, 47.72255, 47.9502, 48.17718, 
    48.4035, 48.62915, 48.85413, 49.07844, 49.30208, 49.52505, 49.74735, 
    49.96898, 50.18993, 50.41021, 50.62981, 50.84874, 51.067, 51.28458, 
    51.50148, 51.71771, 51.93327, 52.14814, 52.36235, 52.57587, 52.78873, 
    53.0009, 53.2124, 53.42323, 53.63338, 53.84286, 54.05166, 54.2598, 
    54.46725, 54.67404, 54.88016, 55.0856, 55.29037, 55.49448, 55.69792, 
    55.90069, 56.10279, 56.30423, 56.505, 56.70512, 56.90456, 57.10335, 
    57.30148, 57.49894, 57.69575, 57.8919, 58.0874, 58.28224, 58.47643, 
    58.66997, 58.86286, 59.0551, 59.24669, 59.43764,
  -38.75502, -38.61524, -38.47502, -38.33434, -38.19321, -38.05162, 
    -37.90957, -37.76706, -37.62408, -37.48064, -37.33673, -37.19236, 
    -37.0475, -36.90218, -36.75637, -36.61008, -36.46332, -36.31607, 
    -36.16833, -36.0201, -35.87138, -35.72217, -35.57246, -35.42225, 
    -35.27155, -35.12033, -34.96862, -34.8164, -34.66367, -34.51042, 
    -34.35666, -34.20238, -34.04759, -33.89228, -33.73643, -33.58007, 
    -33.42318, -33.26575, -33.1078, -32.9493, -32.79027, -32.6307, -32.47059, 
    -32.30993, -32.14873, -31.98698, -31.82467, -31.66181, -31.4984, 
    -31.33443, -31.1699, -31.0048, -30.83914, -30.67291, -30.50612, 
    -30.33875, -30.17081, -30.00229, -29.83319, -29.66352, -29.49325, 
    -29.32241, -29.15098, -28.97895, -28.80634, -28.63313, -28.45933, 
    -28.28493, -28.10993, -27.93432, -27.75812, -27.5813, -27.40388, 
    -27.22585, -27.0472, -26.86794, -26.68806, -26.50757, -26.32645, 
    -26.14472, -25.96235, -25.77937, -25.59575, -25.4115, -25.22663, 
    -25.04111, -24.85497, -24.66818, -24.48076, -24.2927, -24.10399, 
    -23.91464, -23.72464, -23.534, -23.34271, -23.15077, -22.95817, 
    -22.76492, -22.57102, -22.37646, -22.18124, -21.98537, -21.78883, 
    -21.59163, -21.39377, -21.19524, -20.99605, -20.79619, -20.59566, 
    -20.39446, -20.1926, -19.99006, -19.78685, -19.58297, -19.37841, 
    -19.17318, -18.96727, -18.76069, -18.55343, -18.34549, -18.13687, 
    -17.92758, -17.7176, -17.50695, -17.29561, -17.0836, -16.8709, -16.65752, 
    -16.44346, -16.22872, -16.01329, -15.79719, -15.5804, -15.36293, 
    -15.14478, -14.92595, -14.70644, -14.48624, -14.26537, -14.04382, 
    -13.82158, -13.59867, -13.37508, -13.15081, -12.92586, -12.70024, 
    -12.47395, -12.24697, -12.01933, -11.79102, -11.56203, -11.33237, 
    -11.10205, -10.87106, -10.6394, -10.40708, -10.1741, -9.940457, 
    -9.706157, -9.471199, -9.235587, -8.999323, -8.762407, -8.524843, 
    -8.286633, -8.04778, -7.808285, -7.568152, -7.327382, -7.085979, 
    -6.843946, -6.601285, -6.357998, -6.11409, -5.869564, -5.624423, 
    -5.378668, -5.132306, -4.885338, -4.637769, -4.389602, -4.140841, 
    -3.891489, -3.641551, -3.39103, -3.139931, -2.888259, -2.636016, 
    -2.383209, -2.12984, -1.875915, -1.621439, -1.366415, -1.11085, 
    -0.8547477, -0.5981133, -0.3409519, -0.08326896, 0.1749304, 0.4336408, 
    0.6928567, 0.9525726, 1.212783, 1.473481, 1.734663, 1.996321, 2.25845, 
    2.521044, 2.784096, 3.0476, 3.31155, 3.57594, 3.840762, 4.106011, 
    4.371679, 4.63776, 4.904248, 5.171134, 5.438412, 5.706076, 5.974117, 
    6.242528, 6.511303, 6.780434, 7.049913, 7.319734, 7.589887, 7.860366, 
    8.131164, 8.402271, 8.67368, 8.945384, 9.217375, 9.489643, 9.762182, 
    10.03498, 10.30804, 10.58134, 10.85488, 11.12864, 11.40263, 11.67683, 
    11.95123, 12.22583, 12.50061, 12.77557, 13.0507, 13.326, 13.60144, 
    13.87702, 14.15274, 14.42859, 14.70455, 14.98061, 15.25678, 15.53304, 
    15.80937, 16.08578, 16.36225, 16.63877, 16.91534, 17.19195, 17.46858, 
    17.74523, 18.02188, 18.29854, 18.57518, 18.85181, 19.12841, 19.40497, 
    19.68149, 19.95795, 20.23434, 20.51067, 20.78691, 21.06306, 21.33911, 
    21.61506, 21.89088, 22.16658, 22.44214, 22.71756, 22.99283, 23.26793, 
    23.54287, 23.81762, 24.09219, 24.36656, 24.64072, 24.91468, 25.18841, 
    25.46191, 25.73517, 26.00819, 26.28095, 26.55344, 26.82567, 27.09761, 
    27.36927, 27.64063, 27.91169, 28.18244, 28.45287, 28.72297, 28.99274, 
    29.26216, 29.53124, 29.79995, 30.06831, 30.33629, 30.60389, 30.87111, 
    31.13793, 31.40436, 31.67037, 31.93598, 32.20116, 32.46591, 32.73023, 
    32.99411, 33.25755, 33.52053, 33.78305, 34.0451, 34.30668, 34.56779, 
    34.82841, 35.08854, 35.34818, 35.60732, 35.86595, 36.12407, 36.38166, 
    36.63874, 36.89529, 37.15131, 37.40679, 37.66173, 37.91612, 38.16996, 
    38.42324, 38.67595, 38.92811, 39.17969, 39.4307, 39.68113, 39.93097, 
    40.18023, 40.4289, 40.67697, 40.92445, 41.17132, 41.41758, 41.66324, 
    41.90829, 42.15271, 42.39652, 42.63971, 42.88227, 43.12421, 43.36551, 
    43.60618, 43.84621, 44.08561, 44.32436, 44.56247, 44.79993, 45.03674, 
    45.2729, 45.50841, 45.74326, 45.97746, 46.211, 46.44387, 46.67609, 
    46.90764, 47.13853, 47.36874, 47.5983, 47.82718, 48.05539, 48.28292, 
    48.50979, 48.73598, 48.96149, 49.18633, 49.41049, 49.63398, 49.85678, 
    50.07891, 50.30035, 50.52112, 50.74121, 50.96061, 51.17934, 51.39738, 
    51.61474, 51.83142, 52.04742, 52.26273, 52.47737, 52.69132, 52.90459, 
    53.11718, 53.32909, 53.54031, 53.75086, 53.96073, 54.16992, 54.37843, 
    54.58626, 54.79341, 54.99989, 55.20569, 55.41081, 55.61526, 55.81904, 
    56.02214, 56.22458, 56.42633, 56.62743, 56.82785, 57.0276, 57.22669, 
    57.42511, 57.62287, 57.81996, 58.0164, 58.21217, 58.40728, 58.60174, 
    58.79554, 58.98868, 59.18117, 59.37301, 59.5642,
  -38.88939, -38.74966, -38.60947, -38.46882, -38.32772, -38.18616, 
    -38.04414, -37.90166, -37.75871, -37.61529, -37.4714, -37.32704, 
    -37.18221, -37.0369, -36.8911, -36.74483, -36.59807, -36.45083, -36.3031, 
    -36.15487, -36.00616, -35.85694, -35.70723, -35.55702, -35.40631, 
    -35.25509, -35.10336, -34.95113, -34.79838, -34.64512, -34.49134, 
    -34.33704, -34.18222, -34.02688, -33.87101, -33.71462, -33.55769, 
    -33.40023, -33.24223, -33.0837, -32.92462, -32.76501, -32.60484, 
    -32.44413, -32.28288, -32.12107, -31.9587, -31.79578, -31.6323, 
    -31.46826, -31.30366, -31.13848, -30.97275, -30.80644, -30.63956, 
    -30.4721, -30.30407, -30.13546, -29.96626, -29.79648, -29.62612, 
    -29.45517, -29.28362, -29.11149, -28.93876, -28.76542, -28.5915, 
    -28.41697, -28.24183, -28.0661, -27.88975, -27.71279, -27.53522, 
    -27.35704, -27.17824, -26.99882, -26.81878, -26.63812, -26.45683, 
    -26.27492, -26.09238, -25.90921, -25.72541, -25.54097, -25.35589, 
    -25.17018, -24.98383, -24.79684, -24.6092, -24.42092, -24.23199, 
    -24.04242, -23.85219, -23.66131, -23.46977, -23.27759, -23.08474, 
    -22.89124, -22.69707, -22.50225, -22.30676, -22.11061, -21.91379, 
    -21.71631, -21.51815, -21.31933, -21.11984, -20.91967, -20.71883, 
    -20.51732, -20.31513, -20.11227, -19.90872, -19.7045, -19.4996, 
    -19.29402, -19.08776, -18.88081, -18.67318, -18.46487, -18.25588, 
    -18.0462, -17.83583, -17.62478, -17.41304, -17.20062, -16.98751, 
    -16.77371, -16.55922, -16.34405, -16.12819, -15.91164, -15.6944, 
    -15.47647, -15.25786, -15.03855, -14.81856, -14.59789, -14.37652, 
    -14.15447, -13.93174, -13.70832, -13.48421, -13.25942, -13.03394, 
    -12.80779, -12.58095, -12.35343, -12.12523, -11.89635, -11.6668, 
    -11.43657, -11.20566, -10.97408, -10.74183, -10.5089, -10.27531, 
    -10.04105, -9.806128, -9.570539, -9.33429, -9.097381, -8.859814, 
    -8.621592, -8.382716, -8.143191, -7.903017, -7.662197, -7.420734, 
    -7.178632, -6.935891, -6.692515, -6.448508, -6.203873, -5.958611, 
    -5.712728, -5.466225, -5.219107, -4.971376, -4.723038, -4.474094, 
    -4.224549, -3.974408, -3.723673, -3.472348, -3.220439, -2.967949, 
    -2.714883, -2.461245, -2.207038, -1.95227, -1.696943, -1.441062, 
    -1.184633, -0.9276603, -0.6701493, -0.4121049, -0.1535324, 0.1055628, 
    0.3651753, 0.6252995, 0.8859299, 1.147061, 1.408686, 1.6708, 1.933397, 
    2.196471, 2.460015, 2.724023, 2.988489, 3.253407, 3.51877, 3.784571, 
    4.050804, 4.317462, 4.584538, 4.852026, 5.119917, 5.388206, 5.656885, 
    5.925946, 6.195383, 6.465188, 6.735353, 7.005871, 7.276735, 7.547936, 
    7.819468, 8.091321, 8.363489, 8.635963, 8.908735, 9.181798, 9.455143, 
    9.728761, 10.00264, 10.27679, 10.55118, 10.82581, 11.10067, 11.37576, 
    11.65106, 11.92656, 12.20227, 12.47816, 12.75424, 13.03048, 13.30689, 
    13.58345, 13.86015, 14.137, 14.41396, 14.69105, 14.96824, 15.24554, 
    15.52293, 15.80039, 16.07793, 16.35553, 16.63319, 16.91089, 17.18863, 
    17.4664, 17.74418, 18.02197, 18.29976, 18.57754, 18.8553, 19.13304, 
    19.41073, 19.68838, 19.96597, 20.2435, 20.52096, 20.79833, 21.07561, 
    21.35279, 21.62986, 21.90681, 22.18363, 22.46031, 22.73685, 23.01323, 
    23.28945, 23.56549, 23.84136, 24.11703, 24.39251, 24.66777, 24.94283, 
    25.21765, 25.49224, 25.7666, 26.0407, 26.31454, 26.58811, 26.86142, 
    27.13443, 27.40716, 27.67958, 27.9517, 28.22351, 28.49499, 28.76613, 
    29.03694, 29.30741, 29.57751, 29.84726, 30.11664, 30.38564, 30.65426, 
    30.92249, 31.19031, 31.45774, 31.72475, 31.99134, 32.2575, 32.52324, 
    32.78853, 33.05338, 33.31777, 33.5817, 33.84517, 34.10817, 34.37069, 
    34.63273, 34.89428, 35.15533, 35.41588, 35.67593, 35.93546, 36.19447, 
    36.45296, 36.71092, 36.96835, 37.22523, 37.48158, 37.73737, 37.99261, 
    38.24729, 38.5014, 38.75495, 39.00793, 39.26033, 39.51214, 39.76337, 
    40.01402, 40.26406, 40.51351, 40.76236, 41.0106, 41.25824, 41.50526, 
    41.75166, 41.99745, 42.24261, 42.48715, 42.73106, 42.97433, 43.21697, 
    43.45897, 43.70033, 43.94105, 44.18112, 44.42055, 44.65932, 44.89744, 
    45.1349, 45.3717, 45.60785, 45.84333, 46.07815, 46.31231, 46.54579, 
    46.77861, 47.01075, 47.24223, 47.47303, 47.70316, 47.9326, 48.16137, 
    48.38947, 48.61687, 48.84361, 49.06966, 49.29502, 49.51971, 49.7437, 
    49.96702, 50.18964, 50.41159, 50.63284, 50.85341, 51.07329, 51.29248, 
    51.51099, 51.72881, 51.94593, 52.16238, 52.37813, 52.5932, 52.80757, 
    53.02126, 53.23426, 53.44658, 53.65821, 53.86915, 54.07941, 54.28898, 
    54.49787, 54.70607, 54.91359, 55.12043, 55.32658, 55.53206, 55.73685, 
    55.94096, 56.1444, 56.34716, 56.54924, 56.75065, 56.95138, 57.15144, 
    57.35083, 57.54955, 57.74759, 57.94497, 58.14168, 58.33773, 58.53311, 
    58.72783, 58.92189, 59.11529, 59.30803, 59.50011, 59.69155,
  -39.02434, -38.88464, -38.74449, -38.60388, -38.46281, -38.32129, 
    -38.17929, -38.03684, -37.89392, -37.75053, -37.60666, -37.46232, 
    -37.31751, -37.17221, -37.02644, -36.88018, -36.73344, -36.5862, 
    -36.43848, -36.29026, -36.14155, -35.99234, -35.84263, -35.69242, 
    -35.5417, -35.39048, -35.23875, -35.0865, -34.93374, -34.78046, 
    -34.62667, -34.47235, -34.31751, -34.16214, -34.00625, -33.84982, 
    -33.69286, -33.53537, -33.37734, -33.21877, -33.05965, -32.89999, 
    -32.73978, -32.57902, -32.41771, -32.25584, -32.09342, -31.93044, 
    -31.76689, -31.60279, -31.43811, -31.27287, -31.10705, -30.94067, 
    -30.7737, -30.60616, -30.43804, -30.26933, -30.10005, -29.93017, 
    -29.7597, -29.58865, -29.41699, -29.24475, -29.0719, -28.89845, -28.7244, 
    -28.54975, -28.37448, -28.19861, -28.02213, -27.84503, -27.66731, 
    -27.48898, -27.31003, -27.13046, -26.95025, -26.76943, -26.58797, 
    -26.40589, -26.22317, -26.03982, -25.85583, -25.67121, -25.48594, 
    -25.30003, -25.11347, -24.92627, -24.73843, -24.54993, -24.36078, 
    -24.17098, -23.98052, -23.78941, -23.59763, -23.4052, -23.21211, 
    -23.01835, -22.82393, -22.62884, -22.43308, -22.23666, -22.03956, 
    -21.84179, -21.64335, -21.44423, -21.24444, -21.04397, -20.84282, 
    -20.64099, -20.43848, -20.23528, -20.03141, -19.82685, -19.6216, 
    -19.41567, -19.20906, -19.00175, -18.79376, -18.58507, -18.3757, 
    -18.16564, -17.95488, -17.74343, -17.53129, -17.31846, -17.10494, 
    -16.89072, -16.6758, -16.4602, -16.2439, -16.0269, -15.80921, -15.59083, 
    -15.37175, -15.15198, -14.93151, -14.71035, -14.48849, -14.26595, 
    -14.04271, -13.81878, -13.59415, -13.36884, -13.14283, -12.91614, 
    -12.68876, -12.46069, -12.23193, -12.00249, -11.77237, -11.54156, 
    -11.31007, -11.07789, -10.84504, -10.61152, -10.37731, -10.14243, 
    -9.906882, -9.670661, -9.433771, -9.196216, -8.957994, -8.719111, 
    -8.479568, -8.239367, -7.99851, -7.757001, -7.514842, -7.272036, 
    -7.028584, -6.784491, -6.539759, -6.294392, -6.048391, -5.801762, 
    -5.554506, -5.306628, -5.058131, -4.809018, -4.559294, -4.308961, 
    -4.058024, -3.806487, -3.554354, -3.30163, -3.048317, -2.794421, 
    -2.539947, -2.284898, -2.029279, -1.773096, -1.516353, -1.259054, 
    -1.001205, -0.742811, -0.4838772, -0.2244088, 0.03558867, 0.2961098, 
    0.5571491, 0.8187007, 1.080759, 1.343318, 1.606372, 1.869915, 2.13394, 
    2.398443, 2.663414, 2.92885, 3.194743, 3.461087, 3.727875, 3.9951, 
    4.262756, 4.530835, 4.799331, 5.068236, 5.337543, 5.607246, 5.877336, 
    6.147807, 6.41865, 6.689859, 6.961425, 7.233341, 7.5056, 7.778193, 
    8.051112, 8.324349, 8.597898, 8.871748, 9.145892, 9.420322, 9.695029, 
    9.970006, 10.24524, 10.52073, 10.79647, 11.07244, 11.34863, 11.62504, 
    11.90166, 12.17849, 12.4555, 12.7327, 13.01007, 13.2876, 13.56529, 
    13.84313, 14.1211, 14.3992, 14.67743, 14.95576, 15.23419, 15.51272, 
    15.79133, 16.07001, 16.34875, 16.62756, 16.9064, 17.18529, 17.4642, 
    17.74312, 18.02206, 18.301, 18.57992, 18.85883, 19.13771, 19.41655, 
    19.69534, 19.97408, 20.25275, 20.53135, 20.80986, 21.08828, 21.36659, 
    21.6448, 21.92288, 22.20083, 22.47865, 22.75631, 23.03382, 23.31116, 
    23.58833, 23.86531, 24.14211, 24.4187, 24.69507, 24.97123, 25.24717, 
    25.52286, 25.79831, 26.07351, 26.34844, 26.62311, 26.89749, 27.17159, 
    27.44539, 27.71889, 27.99208, 28.26495, 28.53749, 28.80969, 29.08156, 
    29.35307, 29.62422, 29.895, 30.16541, 30.43544, 30.70508, 30.97433, 
    31.24317, 31.5116, 31.77961, 32.0472, 32.31435, 32.58107, 32.84735, 
    33.11317, 33.37853, 33.64343, 33.90786, 34.17181, 34.43527, 34.69825, 
    34.96073, 35.22271, 35.48418, 35.74514, 36.00557, 36.26549, 36.52487, 
    36.78372, 37.04203, 37.29979, 37.557, 37.81366, 38.06975, 38.32528, 
    38.58024, 38.83462, 39.08842, 39.34164, 39.59428, 39.84632, 40.09776, 
    40.3486, 40.59883, 40.84846, 41.09748, 41.34588, 41.59366, 41.84082, 
    42.08735, 42.33325, 42.57851, 42.82315, 43.06714, 43.31049, 43.55319, 
    43.79525, 44.03665, 44.2774, 44.5175, 44.75694, 44.99572, 45.23384, 
    45.47129, 45.70807, 45.94419, 46.17963, 46.4144, 46.6485, 46.88192, 
    47.11467, 47.34673, 47.57811, 47.80882, 48.03883, 48.26817, 48.49681, 
    48.72477, 48.95205, 49.17863, 49.40453, 49.62973, 49.85424, 50.07807, 
    50.3012, 50.52364, 50.74538, 50.96643, 51.18679, 51.40645, 51.62542, 
    51.84369, 52.06127, 52.27816, 52.49435, 52.70985, 52.92465, 53.13876, 
    53.35217, 53.5649, 53.77693, 53.98827, 54.19891, 54.40887, 54.61813, 
    54.82671, 55.03459, 55.24179, 55.4483, 55.65412, 55.85925, 56.06371, 
    56.26747, 56.47056, 56.67296, 56.87468, 57.07572, 57.27608, 57.47577, 
    57.67478, 57.87312, 58.07078, 58.26777, 58.46409, 58.65974, 58.85472, 
    59.04904, 59.24269, 59.43568, 59.62801, 59.81968,
  -39.15986, -39.02021, -38.88009, -38.73952, -38.59849, -38.457, -38.31504, 
    -38.17262, -38.02972, -37.88636, -37.74252, -37.59821, -37.45341, 
    -37.30814, -37.16239, -37.01615, -36.86942, -36.7222, -36.57449, 
    -36.42628, -36.27757, -36.12837, -35.97866, -35.82845, -35.67773, 
    -35.5265, -35.37477, -35.22252, -35.06974, -34.91646, -34.76265, 
    -34.60831, -34.45345, -34.29807, -34.14215, -33.98569, -33.82871, 
    -33.67118, -33.51311, -33.3545, -33.19535, -33.03564, -32.87539, 
    -32.71458, -32.55322, -32.3913, -32.22883, -32.06579, -31.90218, 
    -31.73801, -31.57327, -31.40796, -31.24207, -31.0756, -30.90856, 
    -30.74094, -30.57273, -30.40393, -30.23455, -30.06458, -29.89402, 
    -29.72286, -29.5511, -29.37874, -29.20578, -29.03222, -28.85805, 
    -28.68327, -28.50788, -28.33187, -28.15525, -27.97802, -27.80016, 
    -27.62168, -27.44258, -27.26285, -27.08249, -26.9015, -26.71988, 
    -26.53763, -26.35474, -26.17121, -25.98703, -25.80222, -25.61676, 
    -25.43065, -25.2439, -25.05649, -24.86844, -24.67973, -24.49036, 
    -24.30033, -24.10965, -23.9183, -23.72629, -23.53361, -23.34027, 
    -23.14626, -22.95158, -22.75623, -22.56021, -22.36351, -22.16614, 
    -21.96808, -21.76935, -21.56994, -21.36985, -21.16908, -20.96762, 
    -20.76547, -20.56264, -20.35913, -20.15492, -19.95002, -19.74443, 
    -19.53815, -19.33118, -19.12352, -18.91516, -18.7061, -18.49635, 
    -18.2859, -18.07476, -17.86292, -17.65037, -17.43713, -17.22319, 
    -17.00855, -16.79321, -16.57718, -16.36044, -16.14299, -15.92485, 
    -15.70601, -15.48647, -15.26622, -15.04528, -14.82363, -14.60129, 
    -14.37825, -14.1545, -13.93006, -13.70492, -13.47908, -13.25254, 
    -13.02531, -12.79739, -12.56877, -12.33945, -12.10944, -11.87875, 
    -11.64736, -11.41528, -11.18251, -10.94906, -10.71493, -10.48011, 
    -10.24461, -10.00843, -9.771575, -9.534042, -9.295836, -9.056958, 
    -8.81741, -8.577196, -8.336317, -8.094775, -7.852573, -7.609715, -7.3662, 
    -7.122035, -6.877221, -6.631761, -6.385657, -6.138914, -5.891534, 
    -5.643522, -5.394879, -5.14561, -4.895719, -4.645209, -4.394084, 
    -4.142347, -3.890004, -3.637057, -3.383512, -3.129371, -2.874641, 
    -2.619325, -2.363427, -2.106954, -1.849908, -1.592295, -1.334121, 
    -1.07539, -0.8161067, -0.5562773, -0.2959066, -0.03500031, 0.2264362, 
    0.4883972, 0.750877, 1.01387, 1.27737, 1.541371, 1.805867, 2.070852, 
    2.336319, 2.602262, 2.868675, 3.135552, 3.402884, 3.670667, 3.938892, 
    4.207553, 4.476644, 4.746157, 5.016084, 5.286418, 5.557154, 5.828281, 
    6.099794, 6.371685, 6.643946, 6.91657, 7.189548, 7.462872, 7.736536, 
    8.01053, 8.284847, 8.559478, 8.834415, 9.109652, 9.385177, 9.660983, 
    9.937063, 10.21341, 10.49001, 10.76685, 11.04394, 11.32125, 11.59879, 
    11.87653, 12.15448, 12.43263, 12.71095, 12.98946, 13.26813, 13.54696, 
    13.82594, 14.10506, 14.3843, 14.66367, 14.94315, 15.22274, 15.50241, 
    15.78218, 16.06201, 16.34191, 16.62187, 16.90187, 17.18191, 17.46198, 
    17.74206, 18.02215, 18.30225, 18.58233, 18.86239, 19.14243, 19.42242, 
    19.70237, 19.98226, 20.26208, 20.54183, 20.82149, 21.10106, 21.38053, 
    21.65988, 21.9391, 22.2182, 22.49716, 22.77596, 23.05461, 23.33308, 
    23.61139, 23.8895, 24.16742, 24.44513, 24.72263, 24.99991, 25.27696, 
    25.55376, 25.83032, 26.10663, 26.38266, 26.65843, 26.9339, 27.2091, 
    27.48398, 27.75857, 28.03283, 28.30678, 28.58039, 28.85366, 29.12658, 
    29.39915, 29.67135, 29.94318, 30.21463, 30.4857, 30.75637, 31.02664, 
    31.2965, 31.56595, 31.83497, 32.10357, 32.37172, 32.63943, 32.90669, 
    33.1735, 33.43984, 33.7057, 33.9711, 34.236, 34.50042, 34.76434, 
    35.02776, 35.29068, 35.55307, 35.81495, 36.07631, 36.33713, 36.59742, 
    36.85716, 37.11635, 37.375, 37.63308, 37.89061, 38.14756, 38.40395, 
    38.65975, 38.91497, 39.16961, 39.42366, 39.67711, 39.92996, 40.18221, 
    40.43385, 40.68488, 40.93529, 41.18508, 41.43425, 41.6828, 41.93071, 
    42.17799, 42.42463, 42.67063, 42.91599, 43.1607, 43.40476, 43.64817, 
    43.89093, 44.13303, 44.37447, 44.61524, 44.85535, 45.09479, 45.33356, 
    45.57166, 45.80909, 46.04584, 46.28191, 46.5173, 46.75201, 46.98604, 
    47.21938, 47.45203, 47.68401, 47.91528, 48.14587, 48.37577, 48.60498, 
    48.83349, 49.0613, 49.28843, 49.51485, 49.74058, 49.96561, 50.18994, 
    50.41357, 50.63651, 50.85874, 51.08028, 51.30111, 51.52124, 51.74067, 
    51.9594, 52.17744, 52.39477, 52.6114, 52.82732, 53.04255, 53.25708, 
    53.47091, 53.68404, 53.89647, 54.1082, 54.31924, 54.52958, 54.73922, 
    54.94816, 55.15641, 55.36397, 55.57083, 55.777, 55.98248, 56.18727, 
    56.39137, 56.59477, 56.7975, 56.99953, 57.20088, 57.40155, 57.60153, 
    57.80083, 57.99946, 58.1974, 58.39467, 58.59126, 58.78718, 58.98242, 
    59.17699, 59.3709, 59.56414, 59.75671, 59.94861,
  -39.29596, -39.15635, -39.01628, -38.87575, -38.73476, -38.5933, -38.45138, 
    -38.30899, -38.16613, -38.02279, -37.87899, -37.7347, -37.58993, 
    -37.44468, -37.29895, -37.15273, -37.00602, -36.85881, -36.71111, 
    -36.56292, -36.41422, -36.26503, -36.11533, -35.96512, -35.8144, 
    -35.66317, -35.51143, -35.35918, -35.2064, -35.0531, -34.89928, 
    -34.74493, -34.59006, -34.43465, -34.27871, -34.12223, -33.96522, 
    -33.80766, -33.64957, -33.49092, -33.33173, -33.17199, -33.01169, 
    -32.85084, -32.68943, -32.52747, -32.36493, -32.20184, -32.03817, 
    -31.87394, -31.70913, -31.54375, -31.37779, -31.21125, -31.04414, 
    -30.87643, -30.70814, -30.53926, -30.36979, -30.19972, -30.02906, 
    -29.8578, -29.68594, -29.51348, -29.3404, -29.16673, -28.99244, 
    -28.81754, -28.64202, -28.46589, -28.28914, -28.11176, -27.93377, 
    -27.75515, -27.5759, -27.39602, -27.2155, -27.03435, -26.85257, 
    -26.67014, -26.48708, -26.30337, -26.11902, -25.93402, -25.74837, 
    -25.56207, -25.37512, -25.18751, -24.99924, -24.81032, -24.62073, 
    -24.43049, -24.23957, -24.048, -23.85575, -23.66283, -23.46925, 
    -23.27499, -23.08005, -22.88444, -22.68815, -22.49118, -22.29353, 
    -22.0952, -21.89618, -21.69648, -21.49609, -21.29501, -21.09324, 
    -20.89079, -20.68764, -20.48379, -20.27926, -20.07402, -19.86809, 
    -19.66147, -19.45414, -19.24612, -19.03739, -18.82796, -18.61784, 
    -18.40701, -18.19547, -17.98323, -17.77029, -17.55664, -17.34229, 
    -17.12723, -16.91146, -16.69499, -16.47781, -16.25993, -16.04133, 
    -15.82203, -15.60202, -15.38131, -15.15988, -14.93776, -14.71492, 
    -14.49138, -14.26713, -14.04217, -13.81651, -13.59015, -13.36308, 
    -13.13531, -12.90684, -12.67767, -12.44779, -12.21722, -11.98594, 
    -11.75397, -11.52131, -11.28795, -11.0539, -10.81915, -10.58372, 
    -10.34759, -10.11078, -9.873289, -9.635111, -9.396253, -9.156715, 
    -8.916501, -8.675612, -8.434052, -8.191821, -7.948923, -7.705361, 
    -7.461136, -7.216253, -6.970714, -6.724521, -6.477678, -6.230188, 
    -5.982055, -5.733281, -5.48387, -5.233825, -4.98315, -4.73185, -4.479928, 
    -4.227386, -3.974231, -3.720466, -3.466094, -3.211121, -2.95555, 
    -2.699387, -2.442636, -2.185301, -1.927387, -1.6689, -1.409844, 
    -1.150224, -0.8900453, -0.6293137, -0.3680343, -0.1062126, 0.1561459, 
    0.4190356, 0.6824505, 0.9463848, 1.210833, 1.475788, 1.741244, 2.007196, 
    2.273636, 2.540559, 2.807957, 3.075824, 3.344154, 3.612939, 3.882173, 
    4.151848, 4.421958, 4.692496, 4.963454, 5.234824, 5.5066, 5.778775, 
    6.051339, 6.324286, 6.597609, 6.871299, 7.145348, 7.419748, 7.694491, 
    7.96957, 8.244976, 8.5207, 8.796735, 9.073072, 9.349703, 9.626618, 
    9.903811, 10.18127, 10.45899, 10.73696, 11.01517, 11.29361, 11.57228, 
    11.85116, 12.13025, 12.40953, 12.68901, 12.96866, 13.24848, 13.52846, 
    13.80859, 14.08886, 14.36926, 14.64979, 14.93043, 15.21117, 15.49201, 
    15.77294, 16.05394, 16.335, 16.61612, 16.89729, 17.1785, 17.45973, 
    17.74098, 18.02225, 18.30351, 18.58476, 18.86599, 19.14719, 19.42835, 
    19.70946, 19.99052, 20.27151, 20.55242, 20.83324, 21.11397, 21.39459, 
    21.6751, 21.95548, 22.23573, 22.51584, 22.7958, 23.07559, 23.35521, 
    23.63466, 23.91391, 24.19297, 24.47182, 24.75045, 25.02885, 25.30703, 
    25.58496, 25.86264, 26.14005, 26.4172, 26.69407, 26.97066, 27.24695, 
    27.52294, 27.79861, 28.07397, 28.34899, 28.62368, 28.89803, 29.17202, 
    29.44565, 29.71891, 29.9918, 30.26431, 30.53642, 30.80813, 31.07944, 
    31.35033, 31.6208, 31.89084, 32.16045, 32.42961, 32.69832, 32.96658, 
    33.23437, 33.5017, 33.76854, 34.0349, 34.30078, 34.56616, 34.83103, 
    35.0954, 35.35925, 35.62259, 35.88539, 36.14766, 36.4094, 36.67059, 
    36.93124, 37.19133, 37.45086, 37.70983, 37.96822, 38.22604, 38.48329, 
    38.73995, 38.99602, 39.25149, 39.50637, 39.76065, 40.01432, 40.26738, 
    40.51982, 40.77164, 41.02285, 41.27342, 41.52337, 41.77267, 42.02135, 
    42.26938, 42.51677, 42.76351, 43.0096, 43.25503, 43.49981, 43.74393, 
    43.98739, 44.23018, 44.47231, 44.71376, 44.95454, 45.19465, 45.43408, 
    45.67283, 45.9109, 46.14829, 46.38499, 46.62101, 46.85633, 47.09097, 
    47.32491, 47.55816, 47.79071, 48.02258, 48.25373, 48.4842, 48.71396, 
    48.94303, 49.17139, 49.39905, 49.626, 49.85226, 50.0778, 50.30265, 
    50.52678, 50.75021, 50.97294, 51.19496, 51.41627, 51.63687, 51.85677, 
    52.07596, 52.29444, 52.51221, 52.72928, 52.94564, 53.1613, 53.37624, 
    53.59048, 53.80402, 54.01685, 54.22898, 54.4404, 54.65112, 54.86114, 
    55.07045, 55.27907, 55.48698, 55.6942, 55.90071, 56.10653, 56.31166, 
    56.51608, 56.71982, 56.92286, 57.12521, 57.32686, 57.52783, 57.72812, 
    57.92771, 58.12662, 58.32484, 58.52238, 58.71925, 58.91543, 59.11093, 
    59.30576, 59.49992, 59.69339, 59.8862, 60.07835,
  -39.43264, -39.29307, -39.15305, -39.01256, -38.87161, -38.73019, 
    -38.58831, -38.44596, -38.30313, -38.15983, -38.01606, -37.8718, 
    -37.72706, -37.58184, -37.43613, -37.28992, -37.14323, -36.99605, 
    -36.84837, -36.70019, -36.55151, -36.40232, -36.25263, -36.10243, 
    -35.95172, -35.80049, -35.64875, -35.49649, -35.34371, -35.1904, 
    -35.03657, -34.88221, -34.72733, -34.5719, -34.41594, -34.25945, 
    -34.10241, -33.94483, -33.7867, -33.62803, -33.4688, -33.30902, 
    -33.14869, -32.98779, -32.82634, -32.66432, -32.50174, -32.33859, 
    -32.17487, -32.01058, -31.84571, -31.68026, -31.51424, -31.34763, 
    -31.18043, -31.01265, -30.84428, -30.67531, -30.50576, -30.3356, 
    -30.16484, -29.99349, -29.82152, -29.64895, -29.47578, -29.30199, 
    -29.12758, -28.95256, -28.77693, -28.60067, -28.42379, -28.24628, 
    -28.06814, -27.88938, -27.70998, -27.52995, -27.34929, -27.16798, 
    -26.98603, -26.80344, -26.62021, -26.43633, -26.25179, -26.06661, 
    -25.88077, -25.69428, -25.50713, -25.31932, -25.13085, -24.94172, 
    -24.75192, -24.56145, -24.37031, -24.1785, -23.98602, -23.79287, 
    -23.59904, -23.40453, -23.20934, -23.01347, -22.81692, -22.61968, 
    -22.42175, -22.22314, -22.02384, -21.82384, -21.62316, -21.42178, 
    -21.2197, -21.01693, -20.81347, -20.6093, -20.40443, -20.19886, 
    -19.99259, -19.78562, -19.57794, -19.36956, -19.16047, -18.95067, 
    -18.74017, -18.52895, -18.31703, -18.1044, -17.89105, -17.677, -17.46223, 
    -17.24675, -17.03056, -16.81365, -16.59604, -16.3777, -16.15866, 
    -15.9389, -15.71842, -15.49724, -15.27534, -15.05272, -14.82939, 
    -14.60535, -14.3806, -14.15513, -13.92895, -13.70206, -13.47446, 
    -13.24615, -13.01713, -12.7874, -12.55696, -12.32582, -12.09397, 
    -11.86142, -11.62817, -11.39421, -11.15955, -10.9242, -10.68814, 
    -10.45139, -10.21395, -9.975814, -9.736988, -9.497475, -9.257275, 
    -9.016391, -8.774824, -8.532579, -8.289657, -8.04606, -7.801791, 
    -7.556853, -7.311248, -7.06498, -6.818051, -6.570465, -6.322224, 
    -6.073332, -5.823792, -5.573608, -5.322783, -5.071321, -4.819226, 
    -4.566501, -4.313151, -4.059179, -3.804589, -3.549387, -3.293575, 
    -3.037159, -2.780143, -2.522532, -2.26433, -2.005543, -1.746174, 
    -1.48623, -1.225716, -0.9646354, -0.7029953, -0.4408006, -0.1780567, 
    0.08523062, 0.3490557, 0.6134127, 0.8782957, 1.143699, 1.409616, 1.67604, 
    1.942966, 2.210387, 2.478296, 2.746687, 3.015553, 3.284888, 3.554683, 
    3.824934, 4.095632, 4.36677, 4.638341, 4.910339, 5.182754, 5.45558, 
    5.72881, 6.002435, 6.276448, 6.550841, 6.825606, 7.100735, 7.376221, 
    7.652054, 7.928227, 8.204731, 8.481559, 8.7587, 9.036148, 9.313894, 
    9.591928, 9.870244, 10.14883, 10.42768, 10.70678, 10.98613, 11.26571, 
    11.54552, 11.82555, 12.10579, 12.38622, 12.66685, 12.94766, 13.22864, 
    13.50978, 13.79107, 14.07251, 14.35408, 14.63577, 14.91758, 15.1995, 
    15.48151, 15.76361, 16.04578, 16.32803, 16.61032, 16.89267, 17.17505, 
    17.45747, 17.7399, 18.02234, 18.30478, 18.58721, 18.86962, 19.15199, 
    19.43433, 19.71663, 19.99886, 20.28102, 20.5631, 20.8451, 21.127, 
    21.40879, 21.69047, 21.97202, 22.25344, 22.53471, 22.81582, 23.09677, 
    23.37755, 23.65815, 23.93855, 24.21876, 24.49875, 24.77853, 25.05807, 
    25.33739, 25.61645, 25.89526, 26.1738, 26.45207, 26.73006, 27.00776, 
    27.28516, 27.56225, 27.83903, 28.11548, 28.3916, 28.66738, 28.94281, 
    29.21788, 29.49259, 29.76692, 30.04087, 30.31444, 30.5876, 30.86036, 
    31.13272, 31.40465, 31.67615, 31.94722, 32.21785, 32.48803, 32.75775, 
    33.02701, 33.2958, 33.56411, 33.83195, 34.09929, 34.36614, 34.63248, 
    34.89832, 35.16364, 35.42844, 35.69271, 35.95645, 36.21965, 36.48231, 
    36.74442, 37.00597, 37.26696, 37.52739, 37.78724, 38.04652, 38.30521, 
    38.56332, 38.82084, 39.07776, 39.33408, 39.58979, 39.8449, 40.0994, 
    40.35327, 40.60652, 40.85915, 41.11114, 41.3625, 41.61322, 41.86331, 
    42.11275, 42.36153, 42.60967, 42.85715, 43.10398, 43.35014, 43.59564, 
    43.84047, 44.08464, 44.32813, 44.57094, 44.81308, 45.05454, 45.29531, 
    45.53541, 45.77481, 46.01353, 46.25156, 46.48889, 46.72553, 46.96147, 
    47.19672, 47.43126, 47.66511, 47.89825, 48.1307, 48.36243, 48.59346, 
    48.82379, 49.0534, 49.28231, 49.51051, 49.738, 49.96478, 50.19084, 
    50.41619, 50.64084, 50.86477, 51.08798, 51.31049, 51.53227, 51.75335, 
    51.97371, 52.19336, 52.41229, 52.63051, 52.84801, 53.0648, 53.28088, 
    53.49625, 53.71091, 53.92485, 54.13808, 54.3506, 54.56241, 54.77351, 
    54.98391, 55.19359, 55.40257, 55.61084, 55.81841, 56.02527, 56.23143, 
    56.43689, 56.64164, 56.8457, 57.04905, 57.25172, 57.45368, 57.65495, 
    57.85553, 58.05541, 58.2546, 58.45311, 58.65092, 58.84805, 59.0445, 
    59.24026, 59.43534, 59.62975, 59.82347, 60.01652, 60.20889,
  -39.5699, -39.43039, -39.29041, -39.14996, -39.00906, -38.86769, -38.72584, 
    -38.58353, -38.44074, -38.29748, -38.15373, -38.00951, -37.8648, 
    -37.7196, -37.57392, -37.42775, -37.28108, -37.13392, -36.98626, 
    -36.83809, -36.68943, -36.54025, -36.39057, -36.24038, -36.08968, 
    -35.93845, -35.78672, -35.63446, -35.48167, -35.32837, -35.17453, 
    -35.02016, -34.86526, -34.70982, -34.55385, -34.39734, -34.24028, 
    -34.08267, -33.92452, -33.76582, -33.60656, -33.44674, -33.28637, 
    -33.12544, -32.96395, -32.80188, -32.63926, -32.47606, -32.31228, 
    -32.14793, -31.983, -31.8175, -31.6514, -31.48472, -31.31746, -31.1496, 
    -30.98115, -30.81211, -30.64246, -30.47222, -30.30137, -30.12992, 
    -29.95786, -29.78518, -29.6119, -29.438, -29.26349, -29.08835, -28.91259, 
    -28.73621, -28.5592, -28.38156, -28.20329, -28.02439, -27.84485, 
    -27.66467, -27.48385, -27.30239, -27.12028, -26.93753, -26.75413, 
    -26.57007, -26.38536, -26.2, -26.01398, -25.82729, -25.63995, -25.45194, 
    -25.26327, -25.07392, -24.88391, -24.69323, -24.50187, -24.30983, 
    -24.11712, -23.92373, -23.72965, -23.5349, -23.33945, -23.14333, 
    -22.94651, -22.749, -22.5508, -22.35191, -22.15233, -21.95205, -21.75106, 
    -21.54939, -21.34701, -21.14392, -20.94014, -20.73565, -20.53045, 
    -20.32455, -20.11794, -19.91062, -19.70259, -19.49385, -19.2844, 
    -19.07423, -18.86335, -18.65175, -18.43944, -18.22642, -18.01267, 
    -17.79821, -17.58303, -17.36713, -17.15051, -16.93317, -16.71511, 
    -16.49634, -16.27684, -16.05662, -15.83568, -15.61402, -15.39164, 
    -15.16854, -14.94472, -14.72018, -14.49492, -14.26894, -14.04224, 
    -13.81482, -13.58668, -13.35783, -13.12826, -12.89798, -12.66698, 
    -12.43527, -12.20284, -11.9697, -11.73586, -11.5013, -11.26604, 
    -11.03007, -10.79339, -10.55602, -10.31794, -10.07916, -9.839684, 
    -9.599512, -9.358646, -9.117089, -8.874844, -8.63191, -8.388293, 
    -8.143993, -7.899015, -7.653359, -7.40703, -7.160029, -6.91236, 
    -6.664026, -6.41503, -6.165376, -5.915067, -5.664105, -5.412496, 
    -5.160242, -4.907347, -4.653815, -4.39965, -4.144856, -3.889438, 
    -3.633399, -3.376743, -3.119476, -2.861602, -2.603125, -2.344051, 
    -2.084383, -1.824128, -1.56329, -1.301874, -1.039886, -0.7773309, 
    -0.5142142, -0.2505415, 0.01368151, 0.278449, 0.5437552, 0.809594, 
    1.075959, 1.342845, 1.610245, 1.878153, 2.146562, 2.415466, 2.684858, 
    2.954731, 3.225079, 3.495894, 3.767169, 4.038898, 4.311073, 4.583687, 
    4.856732, 5.130201, 5.404086, 5.67838, 5.953075, 6.228163, 6.503636, 
    6.779486, 7.055705, 7.332285, 7.609218, 7.886494, 8.164107, 8.442047, 
    8.720306, 8.998876, 9.277746, 9.556911, 9.836358, 10.11608, 10.39607, 
    10.67632, 10.95681, 11.23755, 11.51851, 11.7997, 12.08109, 12.36269, 
    12.64448, 12.92646, 13.2086, 13.49092, 13.77339, 14.056, 14.33875, 
    14.62162, 14.90461, 15.18771, 15.47091, 15.75419, 16.03755, 16.32098, 
    16.60447, 16.888, 17.17158, 17.45518, 17.7388, 18.02243, 18.30606, 
    18.58968, 18.87328, 19.15685, 19.44038, 19.72386, 20.00727, 20.29062, 
    20.57389, 20.85707, 21.14016, 21.42313, 21.70599, 21.98872, 22.27131, 
    22.55375, 22.83604, 23.11816, 23.40011, 23.68187, 23.96343, 24.2448, 
    24.52595, 24.80688, 25.08757, 25.36803, 25.64824, 25.92818, 26.20786, 
    26.48727, 26.76639, 27.04521, 27.32373, 27.60194, 27.87983, 28.15739, 
    28.43461, 28.71149, 28.98801, 29.26417, 29.53996, 29.81538, 30.0904, 
    30.36504, 30.63927, 30.91309, 31.18649, 31.45947, 31.73201, 32.00412, 
    32.27577, 32.54697, 32.81772, 33.08799, 33.35779, 33.6271, 33.89593, 
    34.16426, 34.43209, 34.69941, 34.96621, 35.23249, 35.49825, 35.76347, 
    36.02815, 36.29229, 36.55587, 36.8189, 37.08137, 37.34327, 37.60459, 
    37.86533, 38.1255, 38.38507, 38.64405, 38.90244, 39.16021, 39.41738, 
    39.67394, 39.92988, 40.1852, 40.4399, 40.69396, 40.94739, 41.20019, 
    41.45234, 41.70385, 41.9547, 42.20491, 42.45446, 42.70335, 42.95158, 
    43.19915, 43.44604, 43.69226, 43.93781, 44.18268, 44.42688, 44.67038, 
    44.91321, 45.15535, 45.39679, 45.63755, 45.87761, 46.11698, 46.35564, 
    46.59361, 46.83088, 47.06744, 47.3033, 47.53845, 47.7729, 48.00663, 
    48.23965, 48.47197, 48.70357, 48.93445, 49.16462, 49.39408, 49.62282, 
    49.85084, 50.07814, 50.30473, 50.5306, 50.75574, 50.98017, 51.20388, 
    51.42686, 51.64913, 51.87068, 52.0915, 52.31161, 52.53099, 52.74966, 
    52.9676, 53.18482, 53.40133, 53.61712, 53.83218, 54.04653, 54.26016, 
    54.47308, 54.68527, 54.89676, 55.10752, 55.31758, 55.52692, 55.73555, 
    55.94346, 56.15067, 56.35717, 56.56296, 56.76804, 56.97242, 57.17609, 
    57.37907, 57.58133, 57.7829, 57.98377, 58.18394, 58.38342, 58.5822, 
    58.78029, 58.97769, 59.1744, 59.37041, 59.56575, 59.7604, 59.95436, 
    60.14765, 60.34025,
  -39.70775, -39.56829, -39.42836, -39.28796, -39.14711, -39.00578, 
    -38.86398, -38.72171, -38.57896, -38.43573, -38.29203, -38.14783, 
    -38.00316, -37.858, -37.71235, -37.5662, -37.41956, -37.27242, -37.12477, 
    -36.97663, -36.82798, -36.67883, -36.52916, -36.37898, -36.22829, 
    -36.07708, -35.92534, -35.77308, -35.6203, -35.46699, -35.31315, 
    -35.15878, -35.00387, -34.84842, -34.69244, -34.5359, -34.37883, 
    -34.2212, -34.06303, -33.9043, -33.74501, -33.58517, -33.42476, 
    -33.26379, -33.10226, -32.94016, -32.77748, -32.61423, -32.45041, 
    -32.28601, -32.12102, -31.95545, -31.7893, -31.62255, -31.45522, 
    -31.28729, -31.11876, -30.94964, -30.77991, -30.60958, -30.43864, 
    -30.2671, -30.09494, -29.92217, -29.74879, -29.57478, -29.40015, 
    -29.22491, -29.04903, -28.87253, -28.69539, -28.51762, -28.33922, 
    -28.16018, -27.9805, -27.80017, -27.61921, -27.43759, -27.25533, 
    -27.07241, -26.88884, -26.70462, -26.51974, -26.33419, -26.14799, 
    -25.96112, -25.77358, -25.58537, -25.3965, -25.20695, -25.01673, 
    -24.82582, -24.63424, -24.44198, -24.24904, -24.05541, -23.8611, 
    -23.6661, -23.4704, -23.27402, -23.07694, -22.87917, -22.6807, -22.48153, 
    -22.28166, -22.08109, -21.87982, -21.67784, -21.47516, -21.27176, 
    -21.06766, -20.86285, -20.65733, -20.4511, -20.24415, -20.03648, 
    -19.8281, -19.619, -19.40919, -19.19865, -18.98739, -18.77542, -18.56272, 
    -18.3493, -18.13515, -17.92028, -17.70469, -17.48837, -17.27133, 
    -17.05355, -16.83506, -16.61584, -16.39588, -16.17521, -15.9538, 
    -15.73167, -15.50881, -15.28522, -15.06091, -14.83586, -14.6101, 
    -14.3836, -14.15638, -13.92844, -13.69976, -13.47037, -13.24025, 
    -13.00941, -12.77785, -12.54556, -12.31256, -12.07884, -11.84439, 
    -11.60924, -11.37337, -11.13678, -10.89948, -10.66148, -10.42276, 
    -10.18334, -9.943206, -9.702374, -9.460841, -9.218609, -8.975679, 
    -8.732056, -8.48774, -8.242735, -7.997042, -7.750666, -7.503607, 
    -7.255871, -7.007458, -6.758373, -6.508618, -6.258197, -6.007114, 
    -5.755371, -5.502972, -5.249921, -4.996222, -4.741878, -4.486894, 
    -4.231273, -3.97502, -3.718139, -3.460635, -3.202511, -2.943773, 
    -2.684425, -2.424472, -2.163919, -1.902771, -1.641032, -1.378709, 
    -1.115806, -0.8523296, -0.5882842, -0.3236758, -0.05851023, 0.2072068, 
    0.4734693, 0.7402712, 1.007607, 1.275469, 1.543852, 1.812749, 2.082155, 
    2.352061, 2.622462, 2.89335, 3.164719, 3.436561, 3.70887, 3.981639, 
    4.254859, 4.528524, 4.802626, 5.077158, 5.352111, 5.627479, 5.903253, 
    6.179425, 6.455987, 6.732932, 7.01025, 7.287934, 7.565976, 7.844367, 
    8.123098, 8.402161, 8.681547, 8.961248, 9.241255, 9.521559, 9.80215, 
    10.08302, 10.36416, 10.64556, 10.92721, 11.20911, 11.49124, 11.77359, 
    12.05616, 12.33893, 12.6219, 12.90505, 13.18838, 13.47188, 13.75553, 
    14.03933, 14.32327, 14.60734, 14.89152, 15.17581, 15.4602, 15.74468, 
    16.02924, 16.31387, 16.59856, 16.88329, 17.16807, 17.45287, 17.7377, 
    18.02253, 18.30736, 18.59218, 18.87698, 19.16175, 19.44648, 19.73116, 
    20.01577, 20.30032, 20.58479, 20.86917, 21.15344, 21.43761, 21.72165, 
    22.00557, 22.28935, 22.57298, 22.85645, 23.13975, 23.42288, 23.70581, 
    23.98855, 24.27109, 24.5534, 24.8355, 25.11735, 25.39897, 25.68033, 
    25.96143, 26.24225, 26.5228, 26.80306, 27.08302, 27.36267, 27.642, 
    27.92101, 28.19969, 28.47803, 28.75601, 29.03364, 29.3109, 29.58779, 
    29.86429, 30.1404, 30.41611, 30.69141, 30.9663, 31.24076, 31.51479, 
    31.78839, 32.06154, 32.33424, 32.60647, 32.87824, 33.14953, 33.42035, 
    33.69067, 33.96049, 34.22982, 34.49863, 34.76694, 35.03472, 35.30197, 
    35.56868, 35.83486, 36.10049, 36.36557, 36.63009, 36.89405, 37.15743, 
    37.42024, 37.68247, 37.94412, 38.20517, 38.46563, 38.72549, 38.98474, 
    39.24338, 39.50141, 39.75882, 40.0156, 40.27175, 40.52727, 40.78215, 
    41.0364, 41.28999, 41.54294, 41.79523, 42.04688, 42.29786, 42.54817, 
    42.79782, 43.0468, 43.2951, 43.54273, 43.78968, 44.03595, 44.28154, 
    44.52643, 44.77064, 45.01415, 45.25697, 45.49909, 45.74052, 45.98124, 
    46.22126, 46.46057, 46.69917, 46.93707, 47.17425, 47.41072, 47.64648, 
    47.88153, 48.11585, 48.34946, 48.58235, 48.81452, 49.04597, 49.2767, 
    49.5067, 49.73598, 49.96454, 50.19237, 50.41948, 50.64586, 50.87151, 
    51.09644, 51.32064, 51.54411, 51.76685, 51.98887, 52.21016, 52.43073, 
    52.65056, 52.86967, 53.08805, 53.30571, 53.52264, 53.73884, 53.95432, 
    54.16908, 54.38311, 54.59641, 54.809, 55.02086, 55.232, 55.44242, 
    55.65213, 55.86111, 56.06938, 56.27693, 56.48376, 56.68989, 56.8953, 
    57.1, 57.30399, 57.50726, 57.70984, 57.91171, 58.11287, 58.31332, 
    58.51308, 58.71214, 58.9105, 59.10816, 59.30513, 59.5014, 59.69699, 
    59.89188, 60.08609, 60.27961, 60.47244,
  -39.84619, -39.70678, -39.5669, -39.42656, -39.28575, -39.14447, -39.00272, 
    -38.86049, -38.71778, -38.5746, -38.43093, -38.28679, -38.14214, 
    -37.99702, -37.85139, -37.70528, -37.55867, -37.41155, -37.26394, 
    -37.11581, -36.96719, -36.81805, -36.6684, -36.51823, -36.36755, 
    -36.21635, -36.06462, -35.91238, -35.7596, -35.60629, -35.45245, 
    -35.29807, -35.14316, -34.9877, -34.8317, -34.67516, -34.51807, 
    -34.36042, -34.20223, -34.04348, -33.88417, -33.72429, -33.56386, 
    -33.40285, -33.24128, -33.07914, -32.91642, -32.75313, -32.58926, 
    -32.4248, -32.25977, -32.09414, -31.92793, -31.76112, -31.59372, 
    -31.42572, -31.25712, -31.08792, -30.91811, -30.7477, -30.57668, 
    -30.40504, -30.23279, -30.05992, -29.88644, -29.71233, -29.53759, 
    -29.36223, -29.18624, -29.00962, -28.83236, -28.65447, -28.47593, 
    -28.29676, -28.11694, -27.93647, -27.75536, -27.57359, -27.39117, 
    -27.2081, -27.02437, -26.83997, -26.65492, -26.4692, -26.28281, 
    -26.09576, -25.90803, -25.71963, -25.53055, -25.3408, -25.15037, 
    -24.95925, -24.76745, -24.57497, -24.3818, -24.18793, -23.99338, 
    -23.79814, -23.6022, -23.40556, -23.20822, -23.01018, -22.81144, -22.612, 
    -22.41185, -22.21099, -22.00943, -21.80715, -21.60417, -21.40047, 
    -21.19605, -20.99092, -20.78507, -20.5785, -20.37122, -20.16321, 
    -19.95448, -19.74502, -19.53484, -19.32394, -19.11231, -18.89995, 
    -18.68686, -18.47305, -18.2585, -18.04323, -17.82722, -17.61049, 
    -17.39301, -17.17481, -16.95588, -16.73621, -16.5158, -16.29467, 
    -16.07279, -15.85019, -15.62685, -15.40277, -15.17797, -14.95242, 
    -14.72615, -14.49914, -14.27139, -14.04292, -13.81371, -13.58377, 
    -13.3531, -13.1217, -12.88958, -12.65672, -12.42313, -12.18882, 
    -11.95379, -11.71803, -11.48155, -11.24434, -11.00642, -10.76778, 
    -10.52842, -10.28835, -10.04757, -9.806071, -9.563868, -9.320957, 
    -9.077342, -8.833024, -8.588007, -8.342293, -8.095883, -7.848783, 
    -7.600992, -7.352515, -7.103355, -6.853515, -6.602997, -6.351806, 
    -6.099944, -5.847414, -5.594222, -5.34037, -5.085861, -4.830701, 
    -4.574892, -4.318439, -4.061347, -3.803619, -3.54526, -3.286274, 
    -3.026667, -2.766442, -2.505604, -2.244159, -1.982111, -1.719466, 
    -1.456229, -1.192406, -0.9280005, -0.6630197, -0.3974688, -0.1313536, 
    0.13532, 0.402546, 0.6703184, 0.938631, 1.207477, 1.476851, 1.746746, 
    2.017155, 2.288072, 2.55949, 2.831402, 3.1038, 3.376679, 3.65003, 
    3.923847, 4.198121, 4.472846, 4.748014, 5.023618, 5.299648, 5.576099, 
    5.852961, 6.130227, 6.407888, 6.685937, 6.964365, 7.243163, 7.522324, 
    7.801838, 8.081698, 8.361895, 8.642418, 8.923261, 9.204413, 9.485868, 
    9.767612, 10.04964, 10.33194, 10.61451, 10.89733, 11.1804, 11.4637, 
    11.74723, 12.03098, 12.31494, 12.59909, 12.88344, 13.16796, 13.45265, 
    13.7375, 14.0225, 14.30764, 14.59291, 14.8783, 15.1638, 15.4494, 
    15.73508, 16.02085, 16.30669, 16.59259, 16.87854, 17.16452, 17.45054, 
    17.73658, 18.02262, 18.30867, 18.5947, 18.88072, 19.1667, 19.45264, 
    19.73853, 20.02436, 20.31011, 20.59579, 20.88137, 21.16685, 21.45222, 
    21.73747, 22.02259, 22.30757, 22.5924, 22.87706, 23.16155, 23.44587, 
    23.72999, 24.01392, 24.29763, 24.58113, 24.86439, 25.14742, 25.4302, 
    25.71273, 25.99499, 26.27697, 26.55867, 26.84008, 27.12119, 27.40198, 
    27.68245, 27.96259, 28.2424, 28.52186, 28.80096, 29.0797, 29.35807, 
    29.63606, 29.91366, 30.19086, 30.46766, 30.74404, 31.02001, 31.29554, 
    31.57064, 31.84529, 32.1195, 32.39324, 32.66652, 32.93932, 33.21164, 
    33.48348, 33.75481, 34.02565, 34.29598, 34.56579, 34.83508, 35.10385, 
    35.37207, 35.63976, 35.9069, 36.17348, 36.43951, 36.70498, 36.96986, 
    37.23418, 37.49791, 37.76105, 38.0236, 38.28556, 38.54691, 38.80764, 
    39.06777, 39.32728, 39.58617, 39.84443, 40.10206, 40.35905, 40.6154, 
    40.87111, 41.12616, 41.38057, 41.63432, 41.88741, 42.13983, 42.39159, 
    42.64267, 42.89308, 43.14281, 43.39186, 43.64024, 43.88792, 44.13491, 
    44.38121, 44.62681, 44.87172, 45.11592, 45.35943, 45.60223, 45.84432, 
    46.0857, 46.32637, 46.56633, 46.80558, 47.04411, 47.28191, 47.519, 
    47.75537, 47.99102, 48.22594, 48.46013, 48.6936, 48.92634, 49.15836, 
    49.38964, 49.62019, 49.85002, 50.07911, 50.30747, 50.5351, 50.76199, 
    50.98815, 51.21358, 51.43827, 51.66223, 51.88545, 52.10794, 52.3297, 
    52.55072, 52.771, 52.99056, 53.20938, 53.42746, 53.64482, 53.86144, 
    54.07733, 54.29249, 54.50692, 54.72062, 54.93359, 55.14583, 55.35735, 
    55.56814, 55.7782, 55.98754, 56.19616, 56.40405, 56.61123, 56.81768, 
    57.02341, 57.22843, 57.43274, 57.63632, 57.8392, 58.04136, 58.24281, 
    58.44356, 58.6436, 58.84293, 59.04156, 59.23948, 59.43671, 59.63324, 
    59.82907, 60.0242, 60.21865, 60.4124, 60.60546,
  -39.98523, -39.84587, -39.70605, -39.56576, -39.425, -39.28377, -39.14207, 
    -38.99989, -38.85723, -38.71409, -38.57047, -38.42635, -38.28175, 
    -38.13666, -37.99107, -37.84499, -37.69841, -37.55133, -37.40374, 
    -37.25565, -37.10704, -36.95792, -36.80829, -36.65815, -36.50748, 
    -36.35629, -36.20457, -36.05233, -35.89956, -35.74626, -35.59242, 
    -35.43805, -35.28313, -35.12767, -34.97166, -34.81511, -34.658, 
    -34.50034, -34.34213, -34.18336, -34.02402, -33.86413, -33.70366, 
    -33.54263, -33.38102, -33.21885, -33.05609, -32.89275, -32.72884, 
    -32.56433, -32.39924, -32.23356, -32.06729, -31.90042, -31.73296, 
    -31.56489, -31.39622, -31.22695, -31.05707, -30.88657, -30.71547, 
    -30.54374, -30.3714, -30.19844, -30.02486, -29.85065, -29.67581, 
    -29.50034, -29.32424, -29.1475, -28.97012, -28.7921, -28.61344, 
    -28.43413, -28.25418, -28.07357, -27.89231, -27.7104, -27.52783, 
    -27.34459, -27.1607, -26.97614, -26.79092, -26.60502, -26.41846, 
    -26.23122, -26.0433, -25.85471, -25.66544, -25.47548, -25.28484, 
    -25.09352, -24.9015, -24.70879, -24.5154, -24.3213, -24.12651, -23.93103, 
    -23.73484, -23.53795, -23.34035, -23.14205, -22.94304, -22.74333, 
    -22.5429, -22.34176, -22.1399, -21.93733, -21.73404, -21.53003, -21.3253, 
    -21.11985, -20.91368, -20.70678, -20.49916, -20.29081, -20.08173, 
    -19.87192, -19.66138, -19.45011, -19.2381, -19.02536, -18.81189, 
    -18.59768, -18.38274, -18.16706, -17.95064, -17.73348, -17.51559, 
    -17.29695, -17.07758, -16.85746, -16.63661, -16.41501, -16.19267, 
    -15.96959, -15.74577, -15.52121, -15.29591, -15.06986, -14.84308, 
    -14.61555, -14.38729, -14.15828, -13.92854, -13.69805, -13.46683, 
    -13.23487, -13.00218, -12.76875, -12.53458, -12.29968, -12.06405, 
    -11.82768, -11.59059, -11.35277, -11.11422, -10.87494, -10.63494, 
    -10.39422, -10.15278, -9.910615, -9.667738, -9.424146, -9.179841, 
    -8.934827, -8.689106, -8.442678, -8.195549, -7.94772, -7.699194, 
    -7.449974, -7.200062, -6.949462, -6.698177, -6.446211, -6.193566, 
    -5.940247, -5.686256, -5.431597, -5.176275, -4.920293, -4.663655, 
    -4.406365, -4.148428, -3.889848, -3.630629, -3.370775, -3.110292, 
    -2.849184, -2.587456, -2.325113, -2.06216, -1.798602, -1.534445, 
    -1.269693, -1.004353, -0.73843, -0.4719296, -0.2048578, 0.06277964, 
    0.3309765, 0.5997268, 0.8690242, 1.138862, 1.409235, 1.680135, 1.951556, 
    2.223492, 2.495935, 2.768878, 3.042315, 3.316238, 3.59064, 3.865514, 
    4.140851, 4.416646, 4.692889, 4.969573, 5.24669, 5.524233, 5.802193, 
    6.080562, 6.359332, 6.638495, 6.918042, 7.197965, 7.478255, 7.758903, 
    8.039902, 8.321241, 8.602913, 8.884909, 9.167217, 9.449832, 9.732742, 
    10.01594, 10.29941, 10.58316, 10.86716, 11.15141, 11.4359, 11.72062, 
    12.00556, 12.29072, 12.57607, 12.86161, 13.14734, 13.43324, 13.71929, 
    14.0055, 14.29186, 14.57834, 14.86495, 15.15166, 15.43848, 15.72539, 
    16.01238, 16.29944, 16.58656, 16.87373, 17.16095, 17.44819, 17.73545, 
    18.02272, 18.30999, 18.59725, 18.88449, 19.1717, 19.45886, 19.74597, 
    20.03302, 20.32, 20.6069, 20.8937, 21.1804, 21.46699, 21.75345, 22.03978, 
    22.32597, 22.612, 22.89787, 23.18357, 23.46908, 23.7544, 24.03952, 
    24.32443, 24.60912, 24.89357, 25.17778, 25.46174, 25.74544, 26.02888, 
    26.31203, 26.59489, 26.87746, 27.15972, 27.44166, 27.72328, 28.00457, 
    28.28551, 28.56611, 28.84634, 29.1262, 29.40569, 29.68479, 29.9635, 
    30.2418, 30.5197, 30.79717, 31.07422, 31.35084, 31.62701, 31.90273, 
    32.178, 32.4528, 32.72712, 33.00097, 33.27433, 33.5472, 33.81956, 
    34.09141, 34.36275, 34.63357, 34.90386, 35.17361, 35.44282, 35.71148, 
    35.9796, 36.24714, 36.51412, 36.78053, 37.04636, 37.31161, 37.57627, 
    37.84033, 38.10379, 38.36665, 38.6289, 38.89053, 39.15154, 39.41192, 
    39.67168, 39.93079, 40.18927, 40.44711, 40.7043, 40.96083, 41.21671, 
    41.47192, 41.72648, 41.98036, 42.23357, 42.48611, 42.73797, 42.98915, 
    43.23964, 43.48944, 43.73855, 43.98697, 44.23469, 44.4817, 44.72802, 
    44.97363, 45.21853, 45.46273, 45.7062, 45.94897, 46.19102, 46.43235, 
    46.67295, 46.91284, 47.152, 47.39043, 47.62814, 47.86512, 48.10137, 
    48.33688, 48.57167, 48.80572, 49.03904, 49.27161, 49.50346, 49.73456, 
    49.96493, 50.19456, 50.42344, 50.65159, 50.879, 51.10567, 51.3316, 
    51.55678, 51.78123, 52.00493, 52.22789, 52.45011, 52.67159, 52.89233, 
    53.11233, 53.33158, 53.55011, 53.76788, 53.98492, 54.20123, 54.41679, 
    54.63162, 54.84571, 55.05907, 55.27169, 55.48357, 55.69473, 55.90516, 
    56.11485, 56.32381, 56.53205, 56.73956, 56.94634, 57.1524, 57.35774, 
    57.56235, 57.76625, 57.96942, 58.17188, 58.37362, 58.57465, 58.77497, 
    58.97457, 59.17347, 59.37165, 59.56914, 59.76592, 59.96199, 60.15737, 
    60.35205, 60.54604, 60.73932,
  -40.12486, -39.98556, -39.84579, -39.70556, -39.56486, -39.42368, 
    -39.28203, -39.1399, -38.99729, -38.8542, -38.71062, -38.56655, 
    -38.42199, -38.27694, -38.13139, -37.98534, -37.83879, -37.69175, 
    -37.54419, -37.39612, -37.24754, -37.09845, -36.94884, -36.79872, 
    -36.64807, -36.49689, -36.3452, -36.19297, -36.0402, -35.88691, 
    -35.73307, -35.5787, -35.42378, -35.26832, -35.11231, -34.95575, 
    -34.79863, -34.64096, -34.48273, -34.32395, -34.16459, -34.00467, 
    -33.84418, -33.68312, -33.52148, -33.35927, -33.19648, -33.0331, 
    -32.86914, -32.7046, -32.53946, -32.37373, -32.2074, -32.04047, 
    -31.87295, -31.70482, -31.53608, -31.36674, -31.19678, -31.02621, 
    -30.85502, -30.68322, -30.51079, -30.33773, -30.16405, -29.98975, 
    -29.81481, -29.63923, -29.46302, -29.28616, -29.10867, -28.93053, 
    -28.75174, -28.57231, -28.39222, -28.21147, -28.03007, -27.84801, 
    -27.66529, -27.48191, -27.29785, -27.11313, -26.92774, -26.74167, 
    -26.55493, -26.36751, -26.17941, -25.99063, -25.80116, -25.611, 
    -25.42016, -25.22862, -25.03639, -24.84347, -24.64985, -24.45552, 
    -24.2605, -24.06477, -23.86834, -23.6712, -23.47334, -23.27478, 
    -23.07551, -22.87552, -22.67481, -22.47339, -22.27125, -22.06838, 
    -21.86479, -21.66048, -21.45544, -21.24967, -21.04317, -20.83594, 
    -20.62798, -20.41929, -20.20986, -19.9997, -19.7888, -19.57716, 
    -19.36478, -19.15167, -18.93781, -18.72321, -18.50787, -18.29178, 
    -18.07495, -17.85737, -17.63905, -17.41998, -17.20017, -16.97961, 
    -16.7583, -16.53625, -16.31344, -16.08989, -15.86559, -15.64054, 
    -15.41474, -15.18819, -14.9609, -14.73286, -14.50407, -14.27453, 
    -14.04425, -13.81322, -13.58144, -13.34892, -13.11566, -12.88165, 
    -12.6469, -12.41141, -12.17518, -11.93821, -11.7005, -11.46206, 
    -11.22288, -10.98297, -10.74232, -10.50095, -10.25884, -10.01601, 
    -9.772461, -9.528185, -9.283189, -9.037475, -8.791045, -8.543902, 
    -8.29605, -8.047489, -7.798223, -7.548255, -7.297588, -7.046226, 
    -6.794169, -6.541424, -6.287992, -6.033877, -5.779084, -5.523614, 
    -5.267474, -5.010665, -4.753193, -4.495061, -4.236274, -3.976835, 
    -3.71675, -3.456023, -3.194659, -2.932662, -2.670038, -2.40679, 
    -2.142926, -1.878449, -1.613364, -1.347679, -1.081397, -0.8145246, 
    -0.5470677, -0.2790321, -0.01042361, 0.2587515, 0.5284872, 0.798777, 
    1.069615, 1.340994, 1.612907, 1.885348, 2.158311, 2.431787, 2.705771, 
    2.980255, 3.255231, 3.530693, 3.806632, 4.083042, 4.359914, 4.637241, 
    4.915016, 5.193229, 5.471874, 5.750941, 6.030424, 6.310312, 6.590599, 
    6.871275, 7.152332, 7.433762, 7.715555, 7.997703, 8.280196, 8.563026, 
    8.846185, 9.129662, 9.413447, 9.697535, 9.981912, 10.26657, 10.5515, 
    10.83669, 11.12214, 11.40783, 11.69375, 11.9799, 12.26625, 12.55282, 
    12.83957, 13.12652, 13.41363, 13.70091, 13.98834, 14.27592, 14.56363, 
    14.85146, 15.13941, 15.42746, 15.7156, 16.00382, 16.29212, 16.58047, 
    16.86888, 17.15733, 17.44581, 17.73431, 18.02282, 18.31133, 18.59982, 
    18.8883, 19.17674, 19.46514, 19.75349, 20.04177, 20.32999, 20.61811, 
    20.90615, 21.19408, 21.48189, 21.76958, 22.05713, 22.34454, 22.6318, 
    22.91888, 23.2058, 23.49253, 23.77906, 24.06538, 24.35149, 24.63738, 
    24.92303, 25.20844, 25.49359, 25.77848, 26.06309, 26.34742, 26.63146, 
    26.9152, 27.19863, 27.48174, 27.76451, 28.04695, 28.32904, 28.61078, 
    28.89215, 29.17315, 29.45376, 29.73399, 30.01381, 30.29323, 30.57223, 
    30.85081, 31.12895, 31.40666, 31.68391, 31.96071, 32.23705, 32.51291, 
    32.7883, 33.0632, 33.3376, 33.61151, 33.8849, 34.15778, 34.43014, 
    34.70197, 34.97326, 35.24401, 35.51422, 35.78386, 36.05295, 36.32147, 
    36.58941, 36.85678, 37.12356, 37.38974, 37.65534, 37.92033, 38.1847, 
    38.44847, 38.71162, 38.97415, 39.23605, 39.49731, 39.75793, 40.01792, 
    40.27725, 40.53594, 40.79396, 41.05133, 41.30804, 41.56407, 41.81943, 
    42.07412, 42.32812, 42.58145, 42.83409, 43.08603, 43.33729, 43.58784, 
    43.8377, 44.08685, 44.3353, 44.58304, 44.83007, 45.07639, 45.32199, 
    45.56687, 45.81104, 46.05447, 46.29719, 46.53918, 46.78044, 47.02097, 
    47.26076, 47.49982, 47.73815, 47.97575, 48.2126, 48.44871, 48.68409, 
    48.91872, 49.15261, 49.38575, 49.61816, 49.84982, 50.08073, 50.31089, 
    50.54031, 50.76898, 50.99691, 51.22408, 51.45051, 51.67619, 51.90112, 
    52.1253, 52.34874, 52.57142, 52.79336, 53.01455, 53.23499, 53.45469, 
    53.67364, 53.89184, 54.1093, 54.32601, 54.54198, 54.75721, 54.97169, 
    55.18543, 55.39843, 55.61069, 55.82221, 56.03299, 56.24304, 56.45235, 
    56.66093, 56.86877, 57.07589, 57.28226, 57.48792, 57.69284, 57.89704, 
    58.10052, 58.30327, 58.5053, 58.70661, 58.9072, 59.10708, 59.30624, 
    59.50469, 59.70243, 59.89946, 60.09578, 60.29139, 60.48631, 60.68052, 
    60.87403,
  -40.26508, -40.12585, -39.98615, -39.84597, -39.70533, -39.56421, 
    -39.42261, -39.28053, -39.13797, -38.99493, -38.8514, -38.70737, 
    -38.56286, -38.41785, -38.27235, -38.12634, -37.97983, -37.83281, 
    -37.68529, -37.53725, -37.3887, -37.23964, -37.09006, -36.93995, 
    -36.78933, -36.63817, -36.48649, -36.33427, -36.18152, -36.02824, 
    -35.87441, -35.72004, -35.56513, -35.40967, -35.25365, -35.09709, 
    -34.93997, -34.78229, -34.62405, -34.46524, -34.30587, -34.14594, 
    -33.98542, -33.82434, -33.66267, -33.50043, -33.3376, -33.17419, 
    -33.01019, -32.8456, -32.68042, -32.51464, -32.34826, -32.18128, 
    -32.01369, -31.8455, -31.6767, -31.50729, -31.33726, -31.16662, 
    -30.99535, -30.82346, -30.65095, -30.47781, -30.30404, -30.12963, 
    -29.95459, -29.77891, -29.60259, -29.42563, -29.24802, -29.06976, 
    -28.89085, -28.71129, -28.53107, -28.35019, -28.16865, -27.98645, 
    -27.80358, -27.62004, -27.43583, -27.25095, -27.06539, -26.87916, 
    -26.69224, -26.50464, -26.31636, -26.12739, -25.93772, -25.74737, 
    -25.55632, -25.36458, -25.17214, -24.979, -24.78515, -24.5906, -24.39534, 
    -24.19938, -24.0027, -23.80531, -23.60721, -23.40839, -23.20885, 
    -23.00859, -22.80761, -22.6059, -22.40347, -22.20031, -21.99642, 
    -21.79181, -21.58645, -21.38037, -21.17355, -20.96599, -20.7577, 
    -20.54867, -20.33889, -20.12838, -19.91712, -19.70511, -19.49236, 
    -19.27887, -19.06462, -18.84963, -18.63389, -18.4174, -18.20016, 
    -17.98217, -17.76342, -17.54392, -17.32367, -17.10266, -16.8809, 
    -16.65838, -16.43511, -16.21109, -15.98631, -15.76077, -15.53448, 
    -15.30743, -15.07962, -14.85106, -14.62175, -14.39168, -14.16086, 
    -13.92928, -13.69695, -13.46387, -13.23004, -12.99545, -12.76012, 
    -12.52403, -12.2872, -12.04962, -11.8113, -11.57223, -11.33242, 
    -11.09187, -10.85058, -10.60855, -10.36578, -10.12228, -9.878048, 
    -9.633085, -9.387394, -9.140977, -8.893837, -8.645975, -8.397395, 
    -8.1481, -7.898091, -7.647372, -7.395946, -7.143816, -6.890984, 
    -6.637455, -6.383232, -6.128318, -5.872717, -5.616432, -5.359468, 
    -5.101828, -4.843516, -4.584537, -4.324893, -4.064592, -3.803636, 
    -3.54203, -3.279778, -3.016887, -2.75336, -2.489202, -2.224419, 
    -1.959016, -1.692999, -1.426372, -1.159142, -0.8913131, -0.6228927, 
    -0.353886, -0.08429916, 0.1858617, 0.4565903, 0.7278803, 0.9997252, 
    1.272118, 1.545053, 1.818523, 2.092521, 2.367039, 2.642072, 2.917611, 
    3.193649, 3.470179, 3.747194, 4.024684, 4.302644, 4.581065, 4.85994, 
    5.139259, 5.419015, 5.6992, 5.979805, 6.260822, 6.542243, 6.824059, 
    7.10626, 7.38884, 7.671787, 7.955095, 8.238753, 8.522753, 8.807085, 
    9.09174, 9.376709, 9.661983, 9.947551, 10.2334, 10.51953, 10.80593, 
    11.09258, 11.37948, 11.66661, 11.95397, 12.24155, 12.52934, 12.81732, 
    13.10549, 13.39383, 13.68234, 13.97101, 14.25982, 14.54877, 14.83785, 
    15.12703, 15.41633, 15.70571, 15.99518, 16.28472, 16.57433, 16.86399, 
    17.15368, 17.44341, 17.73316, 18.02292, 18.31268, 18.60242, 18.89215, 
    19.18184, 19.47149, 19.76108, 20.05061, 20.34007, 20.62944, 20.91872, 
    21.20789, 21.49694, 21.78587, 22.07466, 22.3633, 22.65179, 22.94011, 
    23.22825, 23.5162, 23.80395, 24.0915, 24.37882, 24.66592, 24.95278, 
    25.23939, 25.52575, 25.81183, 26.09764, 26.38316, 26.66839, 26.95331, 
    27.23791, 27.52219, 27.80614, 28.08974, 28.37299, 28.65588, 28.9384, 
    29.22055, 29.5023, 29.78366, 30.06461, 30.34515, 30.62527, 30.90495, 
    31.1842, 31.46301, 31.74136, 32.01924, 32.29666, 32.5736, 32.85005, 
    33.12601, 33.40147, 33.67642, 33.95086, 34.22477, 34.49816, 34.77101, 
    35.04331, 35.31507, 35.58627, 35.85691, 36.12698, 36.39648, 36.66539, 
    36.93372, 37.20145, 37.46859, 37.73512, 38.00104, 38.26635, 38.53103, 
    38.79509, 39.05851, 39.3213, 39.58345, 39.84496, 40.10581, 40.36601, 
    40.62555, 40.88442, 41.14263, 41.40016, 41.65702, 41.91319, 42.16869, 
    42.42349, 42.6776, 42.93102, 43.18375, 43.43576, 43.68708, 43.93769, 
    44.18758, 44.43676, 44.68523, 44.93298, 45.18, 45.42631, 45.67188, 
    45.91673, 46.16085, 46.40423, 46.64688, 46.88879, 47.12997, 47.3704, 
    47.6101, 47.84905, 48.08725, 48.32471, 48.56143, 48.79739, 49.03261, 
    49.26707, 49.50079, 49.73375, 49.96597, 50.19742, 50.42812, 50.65807, 
    50.88727, 51.11571, 51.34339, 51.57032, 51.79649, 52.02191, 52.24657, 
    52.47048, 52.69363, 52.91603, 53.13767, 53.35856, 53.57869, 53.79807, 
    54.0167, 54.23457, 54.4517, 54.66807, 54.88369, 55.09856, 55.31269, 
    55.52607, 55.7387, 55.95058, 56.16172, 56.37212, 56.58178, 56.7907, 
    56.99887, 57.20631, 57.41302, 57.61898, 57.82422, 58.02872, 58.23249, 
    58.43554, 58.63786, 58.83945, 59.04031, 59.24046, 59.43988, 59.63859, 
    59.83658, 60.03386, 60.23042, 60.42628, 60.62142, 60.81586, 61.00959,
  -40.40591, -40.26674, -40.1271, -39.98699, -39.84641, -39.70535, -39.56381, 
    -39.42179, -39.27928, -39.13629, -38.99281, -38.84883, -38.70437, 
    -38.55941, -38.41394, -38.26797, -38.12151, -37.97453, -37.82704, 
    -37.67904, -37.53053, -37.38149, -37.23193, -37.08186, -36.93126, 
    -36.78012, -36.62846, -36.47626, -36.32353, -36.17025, -36.01644, 
    -35.86208, -35.70717, -35.55171, -35.3957, -35.23914, -35.08201, 
    -34.92432, -34.76608, -34.60726, -34.44788, -34.28792, -34.12739, 
    -33.96628, -33.80459, -33.64232, -33.47946, -33.31602, -33.15198, 
    -32.98735, -32.82212, -32.6563, -32.48987, -32.32284, -32.1552, 
    -31.98695, -31.81809, -31.64861, -31.47851, -31.3078, -31.13646, 
    -30.96449, -30.79189, -30.61867, -30.44481, -30.27031, -30.09517, 
    -29.91939, -29.74297, -29.5659, -29.38817, -29.2098, -29.03077, 
    -28.85108, -28.67073, -28.48973, -28.30805, -28.12571, -27.94269, 
    -27.759, -27.57464, -27.3896, -27.20388, -27.01748, -26.83039, -26.64262, 
    -26.45415, -26.26499, -26.07514, -25.88459, -25.69335, -25.5014, 
    -25.30874, -25.11539, -24.92132, -24.72655, -24.53106, -24.33486, 
    -24.13794, -23.9403, -23.74195, -23.54287, -23.34307, -23.14254, 
    -22.94128, -22.7393, -22.53658, -22.33313, -22.12895, -21.92402, 
    -21.71837, -21.51197, -21.30483, -21.09694, -20.88832, -20.67894, 
    -20.46882, -20.25796, -20.04634, -19.83397, -19.62085, -19.40698, 
    -19.19235, -18.97697, -18.76083, -18.54393, -18.32628, -18.10787, 
    -17.8887, -17.66877, -17.44808, -17.22663, -17.00441, -16.78144, 
    -16.5577, -16.3332, -16.10793, -15.88191, -15.65512, -15.42757, 
    -15.19926, -14.97018, -14.74034, -14.50974, -14.27838, -14.04625, 
    -13.81337, -13.57972, -13.34532, -13.11015, -12.87423, -12.63755, 
    -12.40012, -12.16193, -11.92299, -11.6833, -11.44285, -11.20166, 
    -10.95972, -10.71703, -10.4736, -10.22942, -9.98451, -9.738857, 
    -9.492469, -9.245346, -8.997491, -8.748907, -8.499597, -8.249562, 
    -7.998807, -7.747334, -7.495144, -7.242243, -6.988632, -6.734315, 
    -6.479297, -6.223578, -5.967165, -5.71006, -5.452268, -5.193791, 
    -4.934635, -4.674802, -4.414299, -4.153129, -3.891295, -3.628804, 
    -3.36566, -3.101868, -2.837432, -2.572358, -2.306651, -2.040315, 
    -1.773358, -1.505783, -1.237597, -0.9688055, -0.6994143, -0.4294293, 
    -0.1588566, 0.1122975, 0.3840267, 0.6563247, 0.9291849, 1.202601, 
    1.476565, 1.751071, 2.026113, 2.301682, 2.577772, 2.854375, 3.131484, 
    3.409092, 3.68719, 3.965771, 4.244828, 4.524353, 4.804336, 5.08477, 
    5.365648, 5.64696, 5.928698, 6.210854, 6.493419, 6.776384, 7.059741, 
    7.343481, 7.627594, 7.912072, 8.196906, 8.482086, 8.767603, 9.053447, 
    9.33961, 9.626081, 9.912851, 10.19991, 10.48725, 10.77486, 11.06273, 
    11.35085, 11.63921, 11.9278, 12.21661, 12.50563, 12.79484, 13.08425, 
    13.37384, 13.6636, 13.95351, 14.24357, 14.53377, 14.82409, 15.11454, 
    15.40508, 15.69573, 15.98645, 16.27725, 16.56812, 16.85904, 17.15, 
    17.44099, 17.732, 18.02302, 18.31404, 18.60505, 18.89603, 19.18699, 
    19.47789, 19.76875, 20.05954, 20.35025, 20.64088, 20.93141, 21.22184, 
    21.51214, 21.80232, 22.09236, 22.38225, 22.67198, 22.96154, 23.25092, 
    23.54011, 23.82909, 24.11787, 24.40642, 24.69474, 24.98282, 25.27065, 
    25.55822, 25.84552, 26.13253, 26.41925, 26.70568, 26.99179, 27.27758, 
    27.56305, 27.84817, 28.13295, 28.41737, 28.70143, 28.98511, 29.2684, 
    29.55131, 29.83381, 30.1159, 30.39757, 30.67881, 30.95962, 31.23998, 
    31.51989, 31.79935, 32.07833, 32.35683, 32.63485, 32.91238, 33.18941, 
    33.46593, 33.74194, 34.01743, 34.29239, 34.56681, 34.84069, 35.11401, 
    35.38679, 35.65899, 35.93063, 36.20169, 36.47218, 36.74207, 37.01136, 
    37.28006, 37.54815, 37.81563, 38.08249, 38.34872, 38.61433, 38.8793, 
    39.14364, 39.40733, 39.67037, 39.93276, 40.19448, 40.45555, 40.71595, 
    40.97567, 41.23472, 41.49309, 41.75077, 42.00777, 42.26408, 42.51968, 
    42.77459, 43.0288, 43.2823, 43.53508, 43.78716, 44.03852, 44.28916, 
    44.53908, 44.78828, 45.03675, 45.28448, 45.53149, 45.77776, 46.0233, 
    46.2681, 46.51215, 46.75547, 46.99804, 47.23986, 47.48094, 47.72126, 
    47.96084, 48.19966, 48.43773, 48.67504, 48.9116, 49.1474, 49.38245, 
    49.61673, 49.85025, 50.08302, 50.31503, 50.54627, 50.77675, 51.00647, 
    51.23542, 51.46362, 51.69105, 51.91771, 52.14362, 52.36876, 52.59314, 
    52.81676, 53.03961, 53.26171, 53.48304, 53.70361, 53.92342, 54.14247, 
    54.36076, 54.57829, 54.79507, 55.01109, 55.22635, 55.44086, 55.65461, 
    55.86761, 56.07986, 56.29136, 56.50211, 56.71211, 56.92137, 57.12988, 
    57.33764, 57.54467, 57.75095, 57.95649, 58.16129, 58.36536, 58.5687, 
    58.7713, 58.97317, 59.17431, 59.37472, 59.57441, 59.77337, 59.97161, 
    60.16914, 60.36594, 60.56203, 60.7574, 60.95207, 61.14602,
  -40.54735, -40.40825, -40.26867, -40.12863, -39.98811, -39.84711, 
    -39.70563, -39.56367, -39.42122, -39.27828, -39.13485, -38.99094, 
    -38.84652, -38.7016, -38.55619, -38.41026, -38.26384, -38.1169, 
    -37.96945, -37.82149, -37.67301, -37.52401, -37.37449, -37.22443, 
    -37.07386, -36.92275, -36.77111, -36.61893, -36.46622, -36.31296, 
    -36.15916, -36.00481, -35.84991, -35.69446, -35.53845, -35.38189, 
    -35.22477, -35.06707, -34.90882, -34.75, -34.5906, -34.43063, -34.27008, 
    -34.10896, -33.94724, -33.78495, -33.62206, -33.45859, -33.29452, 
    -33.12985, -32.96458, -32.79872, -32.63224, -32.46516, -32.29747, 
    -32.12917, -31.96024, -31.7907, -31.62054, -31.44976, -31.27835, 
    -31.1063, -30.93363, -30.76032, -30.58637, -30.41178, -30.23655, 
    -30.06067, -29.88415, -29.70697, -29.52914, -29.35065, -29.17151, 
    -28.9917, -28.81123, -28.63008, -28.44828, -28.26579, -28.08264, 
    -27.89881, -27.71429, -27.5291, -27.34322, -27.15665, -26.96939, 
    -26.78144, -26.5928, -26.40346, -26.21342, -26.02268, -25.83123, 
    -25.63908, -25.44622, -25.25265, -25.05837, -24.86337, -24.66765, 
    -24.47122, -24.27406, -24.07618, -23.87757, -23.67824, -23.47818, 
    -23.27738, -23.07586, -22.87359, -22.67059, -22.46685, -22.26237, 
    -22.05715, -21.85118, -21.64447, -21.43701, -21.2288, -21.01984, 
    -20.81013, -20.59967, -20.38845, -20.17647, -19.96374, -19.75025, 
    -19.536, -19.32099, -19.10522, -18.88868, -18.67138, -18.45332, 
    -18.23449, -18.0149, -17.79454, -17.57341, -17.35151, -17.12885, 
    -16.90541, -16.68121, -16.45623, -16.23049, -16.00397, -15.77669, 
    -15.54864, -15.31981, -15.09021, -14.85985, -14.62871, -14.39681, 
    -14.16414, -13.9307, -13.69649, -13.46151, -13.22577, -12.98926, 
    -12.75198, -12.51395, -12.27515, -12.03559, -11.79526, -11.55418, 
    -11.31235, -11.06975, -10.82641, -10.58231, -10.33746, -10.09186, 
    -9.845512, -9.598423, -9.350591, -9.102019, -8.85271, -8.602666, 
    -8.35189, -8.100384, -7.848151, -7.595195, -7.341518, -7.087124, 
    -6.832016, -6.576197, -6.31967, -6.06244, -5.80451, -5.545884, -5.286566, 
    -5.02656, -4.76587, -4.5045, -4.242455, -3.97974, -3.716358, -3.452315, 
    -3.187616, -2.922265, -2.656268, -2.38963, -2.122356, -1.854451, 
    -1.585922, -1.316773, -1.047012, -0.7766424, -0.5056717, -0.2341058, 
    0.03804918, 0.3107868, 0.5841006, 0.857984, 1.13243, 1.407433, 1.682984, 
    1.959077, 2.235706, 2.512862, 2.790538, 3.068727, 3.347421, 3.626613, 
    3.906294, 4.186458, 4.467094, 4.748197, 5.029757, 5.311765, 5.594214, 
    5.877096, 6.160401, 6.44412, 6.728246, 7.012769, 7.297679, 7.582969, 
    7.868628, 8.154648, 8.441019, 8.727733, 9.014777, 9.302145, 9.589827, 
    9.87781, 10.16609, 10.45465, 10.74348, 11.03258, 11.32194, 11.61153, 
    11.90136, 12.19141, 12.48168, 12.77215, 13.06281, 13.35365, 13.64466, 
    13.93583, 14.22715, 14.51861, 14.8102, 15.10191, 15.39373, 15.68564, 
    15.97764, 16.26971, 16.56185, 16.85404, 17.14627, 17.43854, 17.73082, 
    18.02312, 18.31541, 18.6077, 18.89996, 19.19218, 19.48437, 19.77649, 
    20.06856, 20.36054, 20.65244, 20.94424, 21.23593, 21.5275, 21.81894, 
    22.11024, 22.40139, 22.69237, 22.98318, 23.27382, 23.56425, 23.85448, 
    24.1445, 24.43429, 24.72385, 25.01316, 25.30222, 25.59101, 25.87953, 
    26.16776, 26.4557, 26.74333, 27.03065, 27.31764, 27.6043, 27.89062, 
    28.17658, 28.46218, 28.74741, 29.03226, 29.31672, 29.60079, 29.88444, 
    30.16768, 30.45049, 30.73287, 31.01481, 31.2963, 31.57733, 31.85789, 
    32.13798, 32.41758, 32.6967, 32.97531, 33.25342, 33.53101, 33.80809, 
    34.08463, 34.36064, 34.6361, 34.91102, 35.18538, 35.45917, 35.7324, 
    36.00504, 36.2771, 36.54858, 36.81945, 37.08973, 37.35939, 37.62844, 
    37.89687, 38.16468, 38.43185, 38.69839, 38.96428, 39.22953, 39.49413, 
    39.75806, 40.02134, 40.28395, 40.54589, 40.80715, 41.06773, 41.32763, 
    41.58684, 41.84536, 42.10318, 42.36029, 42.61671, 42.87242, 43.12741, 
    43.38169, 43.63526, 43.8881, 44.14022, 44.39161, 44.64227, 44.8922, 
    45.14139, 45.38984, 45.63756, 45.88453, 46.13076, 46.37624, 46.62097, 
    46.86495, 47.10818, 47.35065, 47.59237, 47.83333, 48.07353, 48.31297, 
    48.55165, 48.78957, 49.02672, 49.26311, 49.49873, 49.73359, 49.96767, 
    50.20099, 50.43354, 50.66533, 50.89634, 51.12658, 51.35606, 51.58476, 
    51.81269, 52.03986, 52.26625, 52.49187, 52.71672, 52.9408, 53.16412, 
    53.38666, 53.60844, 53.82944, 54.04969, 54.26916, 54.48787, 54.70581, 
    54.92299, 55.1394, 55.35505, 55.56994, 55.78407, 55.99744, 56.21006, 
    56.42191, 56.63301, 56.84335, 57.05294, 57.26179, 57.46988, 57.67722, 
    57.88381, 58.08966, 58.29477, 58.49913, 58.70275, 58.90564, 59.10778, 
    59.30919, 59.50987, 59.70982, 59.90904, 60.10753, 60.30529, 60.50234, 
    60.69866, 60.89426, 61.08915, 61.28332,
  -40.6894, -40.55037, -40.41086, -40.27088, -40.13043, -39.98949, -39.84808, 
    -39.70618, -39.56379, -39.42091, -39.27754, -39.13367, -38.98931, 
    -38.84444, -38.69908, -38.5532, -38.40682, -38.25993, -38.11252, 
    -37.9646, -37.81616, -37.66719, -37.5177, -37.36769, -37.21714, 
    -37.06606, -36.91445, -36.76229, -36.6096, -36.45636, -36.30258, 
    -36.14824, -35.99335, -35.83791, -35.68192, -35.52536, -35.36823, 
    -35.21054, -35.05229, -34.89346, -34.73405, -34.57407, -34.41351, 
    -34.25237, -34.09064, -33.92832, -33.76541, -33.60191, -33.43781, 
    -33.27311, -33.1078, -32.94189, -32.77538, -32.60825, -32.44051, 
    -32.27216, -32.10318, -31.93358, -31.76336, -31.5925, -31.42102, 
    -31.24891, -31.07616, -30.90277, -30.72874, -30.55406, -30.37874, 
    -30.20277, -30.02614, -29.84886, -29.67093, -29.49233, -29.31307, 
    -29.13314, -28.95255, -28.77128, -28.58934, -28.40672, -28.22342, 
    -28.03945, -27.85479, -27.66944, -27.4834, -27.29667, -27.10925, 
    -26.92113, -26.73231, -26.54279, -26.35256, -26.16163, -25.96999, 
    -25.77764, -25.58457, -25.39079, -25.19629, -25.00107, -24.80513, 
    -24.60846, -24.41107, -24.21295, -24.01409, -23.81451, -23.61419, 
    -23.41313, -23.21133, -23.00879, -22.80551, -22.60148, -22.3967, 
    -22.19118, -21.98491, -21.77789, -21.57011, -21.36157, -21.15228, 
    -20.94224, -20.73143, -20.51986, -20.30753, -20.09444, -19.88058, 
    -19.66595, -19.45056, -19.2344, -19.01747, -18.79977, -18.58129, 
    -18.36205, -18.14203, -17.92124, -17.69967, -17.47733, -17.25421, 
    -17.03032, -16.80565, -16.5802, -16.35397, -16.12697, -15.89919, 
    -15.67063, -15.4413, -15.21118, -14.98029, -14.74862, -14.51617, 
    -14.28295, -14.04895, -13.81418, -13.57863, -13.3423, -13.1052, 
    -12.86733, -12.62869, -12.38928, -12.1491, -11.90815, -11.66643, 
    -11.42394, -11.1807, -10.93669, -10.69192, -10.44639, -10.2001, 
    -9.953062, -9.705269, -9.456725, -9.207433, -8.957395, -8.706613, 
    -8.455091, -8.202831, -7.949836, -7.696109, -7.441653, -7.186471, 
    -6.930567, -6.673943, -6.416604, -6.158553, -5.899793, -5.640328, 
    -5.380164, -5.119303, -4.857749, -4.595508, -4.332583, -4.06898, 
    -3.804701, -3.539754, -3.274142, -3.007869, -2.740943, -2.473367, 
    -2.205148, -1.93629, -1.666799, -1.396681, -1.125942, -0.8545872, 
    -0.5826234, -0.3100566, -0.03689307, 0.2368608, 0.5111984, 0.7861131, 
    1.061598, 1.337647, 1.614252, 1.891406, 2.169102, 2.447333, 2.726092, 
    3.00537, 3.28516, 3.565454, 3.846245, 4.127524, 4.409283, 4.691514, 
    4.974209, 5.257359, 5.540956, 5.824991, 6.109455, 6.39434, 6.679636, 
    6.965335, 7.251428, 7.537905, 7.824757, 8.111974, 8.399548, 8.687468, 
    8.975725, 9.26431, 9.553211, 9.842422, 10.13193, 10.42172, 10.7118, 
    11.00214, 11.29273, 11.58358, 11.87466, 12.16597, 12.45749, 12.74922, 
    13.04114, 13.33325, 13.62553, 13.91797, 14.21057, 14.50331, 14.79618, 
    15.08916, 15.38226, 15.67545, 15.96873, 16.26209, 16.55552, 16.84899, 
    17.14251, 17.43606, 17.72964, 18.02322, 18.3168, 18.61037, 18.90392, 
    19.19744, 19.4909, 19.78432, 20.07766, 20.37093, 20.66411, 20.95719, 
    21.25016, 21.54301, 21.83572, 22.1283, 22.42072, 22.71297, 23.00505, 
    23.29694, 23.58864, 23.88013, 24.1714, 24.46244, 24.75325, 25.04381, 
    25.33411, 25.62414, 25.91389, 26.20335, 26.49251, 26.78136, 27.06989, 
    27.3581, 27.64597, 27.93348, 28.22064, 28.50744, 28.79385, 29.07988, 
    29.36552, 29.65075, 29.93557, 30.21997, 30.50393, 30.78746, 31.07054, 
    31.35316, 31.63532, 31.917, 32.1982, 32.47892, 32.75913, 33.03884, 
    33.31804, 33.59671, 33.87486, 34.15247, 34.42954, 34.70606, 34.98202, 
    35.25741, 35.53223, 35.80648, 36.08014, 36.35321, 36.62568, 36.89755, 
    37.16881, 37.43945, 37.70947, 37.97886, 38.24762, 38.51574, 38.78321, 
    39.05003, 39.3162, 39.58171, 39.84655, 40.11072, 40.37422, 40.63704, 
    40.89917, 41.16061, 41.42136, 41.68142, 41.94077, 42.19942, 42.45736, 
    42.71458, 42.9711, 43.22689, 43.48195, 43.73629, 43.98991, 44.24278, 
    44.49493, 44.74633, 44.99699, 45.24692, 45.49609, 45.74451, 45.99219, 
    46.23911, 46.48528, 46.73069, 46.97534, 47.21923, 47.46235, 47.70472, 
    47.94631, 48.18714, 48.4272, 48.66649, 48.90501, 49.14276, 49.37974, 
    49.61594, 49.85137, 50.08602, 50.3199, 50.55299, 50.78532, 51.01686, 
    51.24763, 51.47762, 51.70684, 51.93527, 52.16293, 52.38981, 52.61591, 
    52.84124, 53.06578, 53.28956, 53.51255, 53.73477, 53.95621, 54.17688, 
    54.39678, 54.61591, 54.83426, 55.05183, 55.26864, 55.48468, 55.69995, 
    55.91446, 56.1282, 56.34117, 56.55338, 56.76483, 56.97551, 57.18544, 
    57.39461, 57.60302, 57.81068, 58.01759, 58.22374, 58.42915, 58.6338, 
    58.83771, 59.04087, 59.2433, 59.44498, 59.64592, 59.84613, 60.0456, 
    60.24434, 60.44234, 60.63962, 60.83617, 61.032, 61.22711, 61.42149,
  -40.83205, -40.6931, -40.55367, -40.41376, -40.27337, -40.1325, -39.99115, 
    -39.84932, -39.70699, -39.56417, -39.42086, -39.27706, -39.13275, 
    -38.98794, -38.84262, -38.6968, -38.55047, -38.40362, -38.25626, 
    -38.10838, -37.95998, -37.81105, -37.66161, -37.51162, -37.36111, 
    -37.21006, -37.05848, -36.90635, -36.75368, -36.60046, -36.4467, 
    -36.29238, -36.13751, -35.98208, -35.82609, -35.66954, -35.51242, 
    -35.35474, -35.19648, -35.03765, -34.87824, -34.71825, -34.55768, 
    -34.39652, -34.23478, -34.07244, -33.90951, -33.74598, -33.58186, 
    -33.41713, -33.25179, -33.08584, -32.91929, -32.75212, -32.58433, 
    -32.41592, -32.24689, -32.07724, -31.90696, -31.73604, -31.5645, 
    -31.39231, -31.21949, -31.04602, -30.87191, -30.69715, -30.52174, 
    -30.34568, -30.16896, -29.99158, -29.81354, -29.63483, -29.45546, 
    -29.27542, -29.0947, -28.91331, -28.73124, -28.54849, -28.36506, 
    -28.18094, -27.99614, -27.81064, -27.62444, -27.43756, -27.24997, 
    -27.06168, -26.87269, -26.68299, -26.49258, -26.30146, -26.10962, 
    -25.91708, -25.72381, -25.52982, -25.33511, -25.13967, -24.9435, 
    -24.74661, -24.54898, -24.35061, -24.15152, -23.95168, -23.7511, 
    -23.54978, -23.34771, -23.1449, -22.94133, -22.73702, -22.53196, 
    -22.32614, -22.11956, -21.91222, -21.70413, -21.49528, -21.28566, 
    -21.07527, -20.86412, -20.65221, -20.43952, -20.22607, -20.01184, 
    -19.79684, -19.58107, -19.36452, -19.14719, -18.92909, -18.71021, 
    -18.49055, -18.2701, -18.04888, -17.82688, -17.60409, -17.38052, 
    -17.15617, -16.93103, -16.70511, -16.4784, -16.25091, -16.02263, 
    -15.79357, -15.56372, -15.33309, -15.10167, -14.86947, -14.63648, 
    -14.4027, -14.16815, -13.93281, -13.69668, -13.45977, -13.22209, 
    -12.98362, -12.74437, -12.50434, -12.26353, -12.02195, -11.77959, 
    -11.53646, -11.29256, -11.04788, -10.80244, -10.55623, -10.30926, 
    -10.06152, -9.813017, -9.563758, -9.313742, -9.062972, -8.81145, 
    -8.559178, -8.306161, -8.052401, -7.797898, -7.542659, -7.286685, 
    -7.02998, -6.772548, -6.514391, -6.255514, -5.995919, -5.735612, 
    -5.474596, -5.212874, -4.950452, -4.687334, -4.423523, -4.159026, 
    -3.893845, -3.627987, -3.361456, -3.094256, -2.826394, -2.557874, 
    -2.288702, -2.018884, -1.748425, -1.47733, -1.205606, -0.933259, 
    -0.6602946, -0.3867193, -0.1125394, 0.1622386, 0.4376082, 0.7135624, 
    0.9900946, 1.267198, 1.544865, 1.823089, 2.101862, 2.381177, 2.661026, 
    2.941403, 3.222298, 3.503705, 3.785614, 4.068018, 4.35091, 4.63428, 
    4.91812, 5.202422, 5.487176, 5.772375, 6.05801, 6.34407, 6.630548, 
    6.917434, 7.20472, 7.492395, 7.78045, 8.068876, 8.357664, 8.646803, 
    8.936284, 9.226096, 9.516232, 9.806678, 10.09743, 10.38847, 10.67979, 
    10.97138, 11.26324, 11.55534, 11.84769, 12.14026, 12.43306, 12.72606, 
    13.01926, 13.31265, 13.60621, 13.89994, 14.19382, 14.48785, 14.782, 
    15.07628, 15.37067, 15.66516, 15.95974, 16.2544, 16.54912, 16.84389, 
    17.13871, 17.43357, 17.72844, 18.02332, 18.31821, 18.61308, 18.90792, 
    19.20274, 19.49751, 19.79222, 20.08686, 20.38143, 20.6759, 20.97027, 
    21.26454, 21.55867, 21.85268, 22.14654, 22.44024, 22.73377, 23.02713, 
    23.3203, 23.61327, 23.90603, 24.19857, 24.49088, 24.78295, 25.07476, 
    25.36631, 25.65759, 25.94858, 26.23929, 26.52968, 26.81977, 27.10953, 
    27.39896, 27.68804, 27.97677, 28.26514, 28.55314, 28.84075, 29.12797, 
    29.41479, 29.70121, 29.9872, 30.27277, 30.5579, 30.84258, 31.12681, 
    31.41058, 31.69387, 31.97669, 32.25901, 32.54084, 32.82217, 33.10298, 
    33.38328, 33.66304, 33.94227, 34.22096, 34.4991, 34.77667, 35.05369, 
    35.33013, 35.60599, 35.88127, 36.15595, 36.43003, 36.70351, 36.97638, 
    37.24863, 37.52026, 37.79125, 38.06161, 38.33133, 38.60039, 38.86881, 
    39.13657, 39.40366, 39.67009, 39.93584, 40.20091, 40.4653, 40.729, 
    40.99201, 41.25432, 41.51593, 41.77684, 42.03703, 42.29651, 42.55527, 
    42.81332, 43.07064, 43.32722, 43.58308, 43.83821, 44.09259, 44.34623, 
    44.59913, 44.85129, 45.10269, 45.35334, 45.60324, 45.85238, 46.10076, 
    46.34837, 46.59523, 46.84132, 47.08664, 47.33119, 47.57497, 47.81798, 
    48.06022, 48.30168, 48.54236, 48.78226, 49.02139, 49.25974, 49.4973, 
    49.73409, 49.97009, 50.2053, 50.43974, 50.67339, 50.90625, 51.13833, 
    51.36963, 51.60014, 51.82986, 52.0588, 52.28695, 52.51432, 52.7409, 
    52.9667, 53.19171, 53.41594, 53.63939, 53.86205, 54.08393, 54.30503, 
    54.52534, 54.74488, 54.96364, 55.18162, 55.39882, 55.61525, 55.8309, 
    56.04578, 56.25988, 56.47322, 56.68578, 56.89758, 57.1086, 57.31887, 
    57.52836, 57.7371, 57.94507, 58.15229, 58.35874, 58.56444, 58.76939, 
    58.97358, 59.17703, 59.37972, 59.58167, 59.78288, 59.98334, 60.18306, 
    60.38204, 60.58029, 60.7778, 60.97458, 61.17063, 61.36596, 61.56055,
  -40.97533, -40.83644, -40.69709, -40.55725, -40.41694, -40.27615, 
    -40.13486, -39.9931, -39.85084, -39.70808, -39.56483, -39.42109, 
    -39.27684, -39.13209, -38.98683, -38.84106, -38.69478, -38.54798, 
    -38.40067, -38.25283, -38.10448, -37.9556, -37.80619, -37.65624, 
    -37.50576, -37.35475, -37.2032, -37.0511, -36.89846, -36.74527, 
    -36.59153, -36.43723, -36.28238, -36.12696, -35.97099, -35.81445, 
    -35.65734, -35.49966, -35.34141, -35.18258, -35.02317, -34.86317, 
    -34.70259, -34.54143, -34.37967, -34.21732, -34.05437, -33.89082, 
    -33.72667, -33.56191, -33.39654, -33.23056, -33.06397, -32.89676, 
    -32.72893, -32.56048, -32.3914, -32.22169, -32.05135, -31.88038, 
    -31.70877, -31.53652, -31.36362, -31.19008, -31.0159, -30.84105, 
    -30.66556, -30.48941, -30.3126, -30.13512, -29.95698, -29.77817, 
    -29.59869, -29.41853, -29.2377, -29.05619, -28.874, -28.69112, -28.50755, 
    -28.32329, -28.13834, -27.9527, -27.76635, -27.57931, -27.39156, 
    -27.20311, -27.01394, -26.82407, -26.63348, -26.44217, -26.25015, 
    -26.0574, -25.86394, -25.66974, -25.47482, -25.27916, -25.08278, 
    -24.88565, -24.68779, -24.48919, -24.28985, -24.08976, -23.88893, 
    -23.68735, -23.48501, -23.28193, -23.07808, -22.87349, -22.66813, 
    -22.46202, -22.25514, -22.04749, -21.83909, -21.62991, -21.41996, 
    -21.20925, -20.99776, -20.7855, -20.57246, -20.35864, -20.14405, 
    -19.92867, -19.71252, -19.49558, -19.27786, -19.05936, -18.84007, 
    -18.61999, -18.39913, -18.17748, -17.95504, -17.73181, -17.50778, 
    -17.28297, -17.05737, -16.83097, -16.60378, -16.3758, -16.14703, 
    -15.91746, -15.6871, -15.45595, -15.224, -14.99127, -14.75773, -14.52341, 
    -14.28829, -14.05238, -13.81568, -13.57819, -13.33991, -13.10084, 
    -12.86098, -12.62034, -12.37891, -12.13669, -11.89369, -11.64991, 
    -11.40535, -11.16001, -10.91389, -10.667, -10.41933, -10.17089, 
    -9.921679, -9.671702, -9.420959, -9.169454, -8.917188, -8.664165, 
    -8.410385, -8.155854, -7.900574, -7.644547, -7.387777, -7.130268, 
    -6.872022, -6.613043, -6.353335, -6.092901, -5.831746, -5.569873, 
    -5.307286, -5.04399, -4.779989, -4.515287, -4.24989, -3.983801, 
    -3.717026, -3.449569, -3.181436, -2.912632, -2.643162, -2.373031, 
    -2.102245, -1.83081, -1.558732, -1.286016, -1.012668, -0.7386957, 
    -0.4641041, -0.1889, 0.0869102, 0.3633197, 0.6403218, 0.9179096, 
    1.196076, 1.474814, 1.754116, 2.033975, 2.314383, 2.595333, 2.876817, 
    3.158827, 3.441355, 3.724393, 4.007934, 4.291967, 4.576486, 4.861482, 
    5.146945, 5.432868, 5.719241, 6.006056, 6.293303, 6.580974, 6.869059, 
    7.157547, 7.446432, 7.735703, 8.025349, 8.315362, 8.605731, 8.896447, 
    9.1875, 9.47888, 9.770576, 10.06258, 10.35488, 10.64746, 10.94032, 
    11.23345, 11.52682, 11.82045, 12.1143, 12.40838, 12.70267, 12.99716, 
    13.29184, 13.58669, 13.88172, 14.1769, 14.47223, 14.76769, 15.06327, 
    15.35897, 15.65477, 15.95065, 16.24662, 16.54265, 16.83874, 17.13487, 
    17.43104, 17.72723, 18.02343, 18.31962, 18.61581, 18.91197, 19.2081, 
    19.50418, 19.8002, 20.09616, 20.39203, 20.68781, 20.98349, 21.27906, 
    21.5745, 21.8698, 22.16496, 22.45996, 22.75479, 23.04944, 23.3439, 
    23.63815, 23.9322, 24.22602, 24.5196, 24.81294, 25.10602, 25.39884, 
    25.69138, 25.98363, 26.27559, 26.56723, 26.85856, 27.14956, 27.44022, 
    27.73054, 28.02049, 28.31008, 28.59929, 28.88811, 29.17654, 29.46456, 
    29.75216, 30.03934, 30.32609, 30.61239, 30.89824, 31.18363, 31.46855, 
    31.75299, 32.03695, 32.32041, 32.60337, 32.88582, 33.16774, 33.44915, 
    33.73001, 34.01033, 34.2901, 34.56932, 34.84797, 35.12604, 35.40353, 
    35.68044, 35.95676, 36.23247, 36.50758, 36.78207, 37.05595, 37.3292, 
    37.60181, 37.87379, 38.14512, 38.41581, 38.68583, 38.9552, 39.2239, 
    39.49192, 39.75927, 40.02594, 40.29192, 40.55721, 40.8218, 41.08569, 
    41.34887, 41.61134, 41.8731, 42.13414, 42.39447, 42.65406, 42.91292, 
    43.17105, 43.42844, 43.6851, 43.94101, 44.19617, 44.45058, 44.70424, 
    44.95714, 45.20929, 45.46067, 45.7113, 45.96115, 46.21024, 46.45856, 
    46.7061, 46.95287, 47.19887, 47.44409, 47.68853, 47.93218, 48.17506, 
    48.41715, 48.65846, 48.89898, 49.13871, 49.37766, 49.61581, 49.85318, 
    50.08975, 50.32553, 50.56053, 50.79473, 51.02813, 51.26075, 51.49257, 
    51.72359, 51.95383, 52.18327, 52.41192, 52.63977, 52.86684, 53.09311, 
    53.31859, 53.54327, 53.76717, 53.99028, 54.21259, 54.43412, 54.65486, 
    54.87481, 55.09398, 55.31236, 55.52995, 55.74676, 55.9628, 56.17804, 
    56.39251, 56.60621, 56.81912, 57.03127, 57.24263, 57.45322, 57.66305, 
    57.8721, 58.08039, 58.28791, 58.49467, 58.70067, 58.9059, 59.11038, 
    59.3141, 59.51707, 59.71928, 59.92075, 60.12146, 60.32143, 60.52066, 
    60.71914, 60.91688, 61.11389, 61.31016, 61.5057, 61.70051,
  -41.11922, -40.98042, -40.84114, -40.70138, -40.56115, -40.42042, 
    -40.27921, -40.13752, -39.99532, -39.85264, -39.70945, -39.56577, 
    -39.42159, -39.27689, -39.13169, -38.98598, -38.83976, -38.69301, 
    -38.54575, -38.39797, -38.24966, -38.10082, -37.95145, -37.80155, 
    -37.65111, -37.50014, -37.34862, -37.19655, -37.04394, -36.89078, 
    -36.73706, -36.58279, -36.42796, -36.27257, -36.11661, -35.96008, 
    -35.80299, -35.64532, -35.48707, -35.32824, -35.16883, -35.00884, 
    -34.84826, -34.68708, -34.52531, -34.36295, -34.19999, -34.03642, 
    -33.87225, -33.70746, -33.54207, -33.37606, -33.20944, -33.04219, 
    -32.87432, -32.70583, -32.5367, -32.36694, -32.19655, -32.02552, 
    -31.85385, -31.68154, -31.50858, -31.33496, -31.1607, -30.98578, 
    -30.81021, -30.63397, -30.45707, -30.2795, -30.10126, -29.92235, 
    -29.74276, -29.5625, -29.38155, -29.19992, -29.0176, -28.8346, -28.6509, 
    -28.46651, -28.28142, -28.09563, -27.90914, -27.72194, -27.53403, 
    -27.34541, -27.15608, -26.96603, -26.77527, -26.58378, -26.39157, 
    -26.19863, -26.00496, -25.81056, -25.61543, -25.41957, -25.22296, 
    -25.02561, -24.82752, -24.62868, -24.4291, -24.22877, -24.02768, 
    -23.82584, -23.62324, -23.41989, -23.21577, -23.01089, -22.80525, 
    -22.59883, -22.39166, -22.18371, -21.97499, -21.76549, -21.55522, 
    -21.34417, -21.13234, -20.91973, -20.70634, -20.49217, -20.27721, 
    -20.06146, -19.84493, -19.62761, -19.40949, -19.19059, -18.97089, 
    -18.7504, -18.52912, -18.30703, -18.08416, -17.86048, -17.63601, 
    -17.41074, -17.18467, -16.9578, -16.73013, -16.50166, -16.27239, 
    -16.04232, -15.81145, -15.57978, -15.3473, -15.11403, -14.87995, 
    -14.64507, -14.40939, -14.17292, -13.93564, -13.69756, -13.45869, 
    -13.21902, -12.97855, -12.73729, -12.49523, -12.25238, -12.00874, 
    -11.76431, -11.51908, -11.27307, -11.02628, -10.7787, -10.53033, 
    -10.28119, -10.03127, -9.780569, -9.529097, -9.276853, -9.023839, 
    -8.770059, -8.515515, -8.26021, -8.004148, -7.747329, -7.489759, 
    -7.231441, -6.972377, -6.712572, -6.452028, -6.19075, -5.928741, 
    -5.666007, -5.402549, -5.138374, -4.873485, -4.607886, -4.341583, 
    -4.07458, -3.806882, -3.538494, -3.26942, -2.999667, -2.72924, -2.458143, 
    -2.186383, -1.913966, -1.640896, -1.367181, -1.092826, -0.8178374, 
    -0.5422217, -0.2659853, 0.01086509, 0.2883229, 0.5663811, 0.8450329, 
    1.124271, 1.404089, 1.684478, 1.965432, 2.246942, 2.529002, 2.811603, 
    3.094737, 3.378397, 3.662574, 3.947259, 4.232445, 4.518124, 4.804285, 
    5.090921, 5.378023, 5.665581, 5.953587, 6.242032, 6.530906, 6.8202, 
    7.109905, 7.40001, 7.690507, 7.981385, 8.272635, 8.564247, 8.856211, 
    9.148516, 9.441152, 9.73411, 10.02738, 10.32095, 10.61481, 10.90894, 
    11.20335, 11.49801, 11.79293, 12.08807, 12.38345, 12.67904, 12.97483, 
    13.27081, 13.56698, 13.86331, 14.15981, 14.45645, 14.75323, 15.05013, 
    15.34715, 15.64427, 15.94148, 16.23877, 16.53612, 16.83354, 17.131, 
    17.42849, 17.72601, 18.02353, 18.32106, 18.61857, 18.91606, 19.21351, 
    19.51092, 19.80827, 20.10554, 20.40274, 20.69984, 20.99684, 21.29373, 
    21.59048, 21.8871, 22.18357, 22.47988, 22.77602, 23.07198, 23.36773, 
    23.66329, 23.95863, 24.25374, 24.54861, 24.84324, 25.1376, 25.4317, 
    25.72551, 26.01903, 26.31225, 26.60516, 26.89775, 27.19, 27.4819, 
    27.77346, 28.06465, 28.35547, 28.64591, 28.93595, 29.22559, 29.51482, 
    29.80362, 30.092, 30.37994, 30.66742, 30.95445, 31.24101, 31.5271, 
    31.8127, 32.09781, 32.38241, 32.66651, 32.95008, 33.23314, 33.51565, 
    33.79763, 34.07905, 34.35991, 34.64021, 34.91994, 35.19909, 35.47764, 
    35.75561, 36.03297, 36.30972, 36.58586, 36.86138, 37.13626, 37.41052, 
    37.68414, 37.9571, 38.22942, 38.50107, 38.77206, 39.04238, 39.31203, 
    39.58099, 39.84927, 40.11686, 40.38375, 40.64995, 40.91543, 41.18021, 
    41.44427, 41.70761, 41.97023, 42.23213, 42.49329, 42.75372, 43.0134, 
    43.27235, 43.53055, 43.788, 44.0447, 44.30065, 44.55583, 44.81025, 
    45.06391, 45.3168, 45.56893, 45.82028, 46.07085, 46.32065, 46.56967, 
    46.81791, 47.06537, 47.31204, 47.55793, 47.80302, 48.04733, 48.29085, 
    48.53357, 48.77551, 49.01664, 49.25698, 49.49653, 49.73528, 49.97322, 
    50.21038, 50.44673, 50.68228, 50.91703, 51.15098, 51.38413, 51.61647, 
    51.84802, 52.07877, 52.30871, 52.53786, 52.7662, 52.99374, 53.22049, 
    53.44643, 53.67157, 53.89592, 54.11946, 54.34222, 54.56417, 54.78533, 
    55.0057, 55.22527, 55.44405, 55.66204, 55.87923, 56.09564, 56.31126, 
    56.5261, 56.74015, 56.95341, 57.1659, 57.37761, 57.58853, 57.79868, 
    58.00805, 58.21665, 58.42448, 58.63154, 58.83783, 59.04335, 59.24811, 
    59.4521, 59.65534, 59.85782, 60.05954, 60.26051, 60.46072, 60.66019, 
    60.85891, 61.05688, 61.25411, 61.4506, 61.64635, 61.84137,
  -41.26373, -41.12502, -40.98582, -40.84614, -40.70598, -40.56533, -40.4242, 
    -40.28257, -40.14046, -39.99784, -39.85473, -39.71111, -39.56699, 
    -39.42236, -39.27722, -39.13157, -38.9854, -38.83872, -38.69151, 
    -38.54378, -38.39552, -38.24673, -38.09741, -37.94755, -37.79716, 
    -37.64622, -37.49474, -37.34271, -37.19014, -37.037, -36.88332, 
    -36.72907, -36.57427, -36.4189, -36.26296, -36.10645, -35.94937, 
    -35.79171, -35.63347, -35.47465, -35.31525, -35.15526, -34.99467, 
    -34.8335, -34.67172, -34.50935, -34.34637, -34.18279, -34.0186, -33.8538, 
    -33.68838, -33.52235, -33.35569, -33.18841, -33.0205, -32.85197, 
    -32.6828, -32.513, -32.34256, -32.17147, -31.99975, -31.82737, -31.65435, 
    -31.48067, -31.30633, -31.13134, -30.95568, -30.77936, -30.60238, 
    -30.42472, -30.24638, -30.06737, -29.88768, -29.70731, -29.52626, 
    -29.34451, -29.16208, -28.97895, -28.79512, -28.6106, -28.42537, 
    -28.23944, -28.0528, -27.86545, -27.67739, -27.48861, -27.29911, 
    -27.10889, -26.91795, -26.72629, -26.53389, -26.34076, -26.1469, 
    -25.9523, -25.75696, -25.56088, -25.36406, -25.16649, -24.96817, 
    -24.7691, -24.56928, -24.3687, -24.16736, -23.96527, -23.76241, 
    -23.55878, -23.35439, -23.14923, -22.9433, -22.7366, -22.52912, 
    -22.32087, -22.11184, -21.90202, -21.69143, -21.48005, -21.26788, 
    -21.05493, -20.84119, -20.62666, -20.41133, -20.19522, -19.9783, 
    -19.7606, -19.54209, -19.32279, -19.10268, -18.88178, -18.66007, 
    -18.43756, -18.21425, -17.99014, -17.76521, -17.53948, -17.31295, 
    -17.08561, -16.85745, -16.6285, -16.39873, -16.16815, -15.93677, 
    -15.70457, -15.47157, -15.23776, -15.00314, -14.76771, -14.53147, 
    -14.29442, -14.05657, -13.81791, -13.57844, -13.33816, -13.09708, 
    -12.8552, -12.61252, -12.36903, -12.12474, -11.87965, -11.63377, 
    -11.38709, -11.13961, -10.89134, -10.64228, -10.39243, -10.14179, 
    -9.89037, -9.638165, -9.385179, -9.131414, -8.876875, -8.621563, 
    -8.36548, -8.108631, -7.851017, -7.592643, -7.333511, -7.073625, 
    -6.812988, -6.551605, -6.289477, -6.026611, -5.763009, -5.498676, 
    -5.233616, -4.967833, -4.701332, -4.434117, -4.166194, -3.897567, 
    -3.628241, -3.358221, -3.087512, -2.816121, -2.544051, -2.27131, 
    -1.997903, -1.723835, -1.449113, -1.173742, -0.8977303, -0.6210827, 
    -0.3438061, -0.06590726, 0.2126071, 0.49173, 0.7714545, 1.051773, 
    1.332679, 1.614165, 1.896222, 2.178845, 2.462023, 2.745751, 3.03002, 
    3.314821, 3.600146, 3.885987, 4.172336, 4.459184, 4.746521, 5.03434, 
    5.322631, 5.611386, 5.900595, 6.190248, 6.480337, 6.770852, 7.061783, 
    7.353121, 7.644856, 7.936978, 8.229477, 8.522343, 8.815566, 9.109135, 
    9.403041, 9.697272, 9.991819, 10.28667, 10.58182, 10.87724, 11.17295, 
    11.46891, 11.76512, 12.06158, 12.35826, 12.65516, 12.95227, 13.24957, 
    13.54706, 13.84472, 14.14254, 14.44051, 14.73862, 15.03685, 15.3352, 
    15.63366, 15.9322, 16.23083, 16.52953, 16.82828, 17.12708, 17.42591, 
    17.72477, 18.02364, 18.3225, 18.62136, 18.92019, 19.21898, 19.51773, 
    19.81641, 20.11503, 20.41356, 20.712, 21.01033, 21.30855, 21.60664, 
    21.90458, 22.20238, 22.50001, 22.79747, 23.09474, 23.39182, 23.68868, 
    23.98533, 24.28175, 24.57792, 24.87385, 25.1695, 25.46489, 25.75999, 
    26.05479, 26.34929, 26.64347, 26.93732, 27.23084, 27.52401, 27.81682, 
    28.10926, 28.40132, 28.69299, 28.98426, 29.27513, 29.56558, 29.8556, 
    30.14518, 30.43432, 30.723, 31.01122, 31.29896, 31.58622, 31.87299, 
    32.15926, 32.44502, 32.73027, 33.01498, 33.29917, 33.58281, 33.8659, 
    34.14843, 34.4304, 34.7118, 34.99261, 35.27283, 35.55246, 35.83149, 
    36.10991, 36.38771, 36.66489, 36.94143, 37.21735, 37.49261, 37.76723, 
    38.04119, 38.3145, 38.58713, 38.8591, 39.13038, 39.40098, 39.67089, 
    39.94011, 40.20862, 40.47643, 40.74353, 41.00992, 41.27559, 41.54054, 
    41.80476, 42.06824, 42.33099, 42.593, 42.85427, 43.11478, 43.37455, 
    43.63356, 43.89182, 44.14931, 44.40604, 44.662, 44.91719, 45.17161, 
    45.42525, 45.67811, 45.93019, 46.18149, 46.43201, 46.68173, 46.93067, 
    47.17881, 47.42616, 47.67272, 47.91848, 48.16344, 48.4076, 48.65096, 
    48.89352, 49.13527, 49.37622, 49.61637, 49.85571, 50.09425, 50.33197, 
    50.56889, 50.805, 51.04031, 51.2748, 51.50848, 51.74136, 51.97342, 
    52.20468, 52.43513, 52.66477, 52.8936, 53.12162, 53.34883, 53.57524, 
    53.80085, 54.02564, 54.24963, 54.47282, 54.6952, 54.91678, 55.13755, 
    55.35753, 55.57671, 55.79509, 56.01267, 56.22945, 56.44545, 56.66064, 
    56.87505, 57.08867, 57.30149, 57.51354, 57.72479, 57.93526, 58.14495, 
    58.35386, 58.562, 58.76935, 58.97593, 59.18174, 59.38678, 59.59105, 
    59.79455, 59.99729, 60.19926, 60.40048, 60.60094, 60.80064, 60.99959, 
    61.19779, 61.39524, 61.59195, 61.78791, 61.98313,
  -41.40887, -41.27024, -41.13113, -40.99153, -40.85146, -40.71089, 
    -40.56983, -40.42828, -40.28624, -40.1437, -40.00066, -39.85711, 
    -39.71305, -39.56849, -39.42342, -39.27783, -39.13173, -38.9851, 
    -38.83795, -38.69027, -38.54207, -38.39333, -38.24406, -38.09425, 
    -37.9439, -37.79301, -37.64157, -37.48958, -37.33704, -37.18394, 
    -37.03029, -36.87608, -36.7213, -36.56595, -36.41004, -36.25355, 
    -36.09649, -35.93885, -35.78062, -35.62181, -35.46242, -35.30243, 
    -35.14185, -34.98067, -34.8189, -34.65652, -34.49353, -34.32994, 
    -34.16573, -34.00091, -33.83548, -33.66942, -33.50274, -33.33543, 
    -33.16749, -32.99892, -32.82971, -32.65986, -32.48937, -32.31824, 
    -32.14646, -31.97403, -31.80094, -31.6272, -31.4528, -31.27773, -31.102, 
    -30.9256, -30.74853, -30.57078, -30.39236, -30.21325, -30.03346, 
    -29.85299, -29.67183, -29.48997, -29.30742, -29.12417, -28.94022, 
    -28.75556, -28.5702, -28.38413, -28.19735, -28.00985, -27.82164, 
    -27.6327, -27.44304, -27.25266, -27.06154, -26.8697, -26.67712, -26.4838, 
    -26.28975, -26.09495, -25.89941, -25.70312, -25.50609, -25.3083, 
    -25.10975, -24.91045, -24.71039, -24.50957, -24.30799, -24.10564, 
    -23.90252, -23.69863, -23.49397, -23.28853, -23.08232, -22.87532, 
    -22.66755, -22.45899, -22.24965, -22.03952, -21.8286, -21.61689, 
    -21.40439, -21.1911, -20.97701, -20.76212, -20.54643, -20.32995, 
    -20.11266, -19.89457, -19.67567, -19.45597, -19.23546, -19.01414, 
    -18.79202, -18.56908, -18.34533, -18.12077, -17.8954, -17.66921, 
    -17.44221, -17.2144, -16.98576, -16.75632, -16.52605, -16.29497, 
    -16.06307, -15.83036, -15.59683, -15.36248, -15.12731, -14.89133, 
    -14.65453, -14.41691, -14.17848, -13.93923, -13.69916, -13.45829, 
    -13.21659, -12.97409, -12.73077, -12.48665, -12.24171, -11.99597, 
    -11.74942, -11.50206, -11.25391, -11.00494, -10.75518, -10.50462, 
    -10.25327, -10.00112, -9.748178, -9.494446, -9.239927, -8.984625, 
    -8.72854, -8.471677, -8.214037, -7.955624, -7.696441, -7.436491, 
    -7.175778, -6.914306, -6.652077, -6.389096, -6.125366, -5.860892, 
    -5.595678, -5.329728, -5.063046, -4.795636, -4.527504, -4.258655, 
    -3.989092, -3.718822, -3.447848, -3.176178, -2.903816, -2.630767, 
    -2.357037, -2.082633, -1.807559, -1.531823, -1.255429, -0.9783857, 
    -0.7006981, -0.4223732, -0.1434176, 0.1361617, 0.4163578, 0.6971637, 
    0.978572, 1.260575, 1.543166, 1.826337, 2.11008, 2.394388, 2.679252, 
    2.964664, 3.250617, 3.537101, 3.824108, 4.111629, 4.399657, 4.688182, 
    4.977195, 5.266686, 5.556648, 5.847071, 6.137944, 6.429259, 6.721006, 
    7.013176, 7.305758, 7.598743, 7.89212, 8.185881, 8.480013, 8.774508, 
    9.069353, 9.36454, 9.660058, 9.955896, 10.25204, 10.54849, 10.84522, 
    11.14223, 11.43951, 11.73704, 12.03481, 12.33282, 12.63104, 12.92948, 
    13.22811, 13.52693, 13.82593, 14.12509, 14.4244, 14.72385, 15.02343, 
    15.32313, 15.62294, 15.92283, 16.22281, 16.52286, 16.82297, 17.12312, 
    17.42331, 17.72352, 18.02374, 18.32397, 18.62418, 18.92436, 19.22451, 
    19.52461, 19.82465, 20.12461, 20.4245, 20.72428, 21.02396, 21.32352, 
    21.62296, 21.92225, 22.22138, 22.52035, 22.81914, 23.11774, 23.41615, 
    23.71434, 24.01231, 24.31004, 24.60753, 24.90477, 25.20173, 25.49842, 
    25.79482, 26.09092, 26.38671, 26.68217, 26.97731, 27.2721, 27.56654, 
    27.86061, 28.15431, 28.44763, 28.74055, 29.03307, 29.32517, 29.61685, 
    29.9081, 30.1989, 30.48925, 30.77914, 31.06855, 31.35749, 31.64594, 
    31.93389, 32.22132, 32.50825, 32.79465, 33.08052, 33.36584, 33.65062, 
    33.93484, 34.21849, 34.50158, 34.78407, 35.06598, 35.34729, 35.62801, 
    35.9081, 36.18758, 36.46644, 36.74467, 37.02225, 37.29919, 37.57548, 
    37.85112, 38.12608, 38.40038, 38.674, 38.94695, 39.2192, 39.49076, 
    39.76162, 40.03178, 40.30123, 40.56997, 40.83798, 41.10528, 41.37185, 
    41.63768, 41.90278, 42.16713, 42.43074, 42.69361, 42.95572, 43.21707, 
    43.47766, 43.73749, 43.99655, 44.25484, 44.51236, 44.7691, 45.02506, 
    45.28024, 45.53463, 45.78824, 46.04106, 46.29308, 46.54431, 46.79475, 
    47.04438, 47.29321, 47.54124, 47.78848, 48.0349, 48.28051, 48.52532, 
    48.76932, 49.0125, 49.25488, 49.49644, 49.73719, 49.97713, 50.21625, 
    50.45455, 50.69204, 50.92871, 51.16457, 51.3996, 51.63382, 51.86723, 
    52.09981, 52.33158, 52.56253, 52.79267, 53.02198, 53.25049, 53.47817, 
    53.70505, 53.9311, 54.15635, 54.38078, 54.6044, 54.82721, 55.04921, 
    55.27039, 55.49078, 55.71035, 55.92912, 56.14708, 56.36424, 56.5806, 
    56.79617, 57.01093, 57.22489, 57.43806, 57.65044, 57.86202, 58.07281, 
    58.28281, 58.49203, 58.70047, 58.90812, 59.11499, 59.32108, 59.52639, 
    59.73093, 59.9347, 60.1377, 60.33993, 60.54139, 60.74209, 60.94203, 
    61.14121, 61.33963, 61.5373, 61.73422, 61.93039, 62.12582,
  -41.55465, -41.4161, -41.27707, -41.13756, -40.99757, -40.85709, -40.71611, 
    -40.57464, -40.43267, -40.29021, -40.14724, -40.00377, -39.85979, 
    -39.7153, -39.57029, -39.42477, -39.27873, -39.13216, -38.98507, 
    -38.83746, -38.68931, -38.54063, -38.39141, -38.24165, -38.09135, 
    -37.94051, -37.78911, -37.63717, -37.48466, -37.33161, -37.17799, 
    -37.02381, -36.86906, -36.71375, -36.55786, -36.40139, -36.24435, 
    -36.08673, -35.92852, -35.76973, -35.61034, -35.45037, -35.28979, 
    -35.12862, -34.96684, -34.80446, -34.64147, -34.47787, -34.31365, 
    -34.14882, -33.98336, -33.81728, -33.65058, -33.48324, -33.31527, 
    -33.14667, -32.97742, -32.80754, -32.63701, -32.46583, -32.294, 
    -32.12151, -31.94837, -31.77456, -31.6001, -31.42496, -31.24916, 
    -31.07269, -30.89553, -30.7177, -30.53919, -30.35999, -30.18011, 
    -29.99953, -29.81827, -29.6363, -29.45364, -29.27027, -29.0862, 
    -28.90142, -28.71593, -28.52972, -28.3428, -28.15515, -27.96679, 
    -27.7777, -27.58788, -27.39733, -27.20605, -27.01403, -26.82127, 
    -26.62777, -26.43353, -26.23853, -26.04279, -25.8463, -25.64905, 
    -25.45104, -25.25228, -25.05275, -24.85246, -24.65139, -24.44956, 
    -24.24696, -24.04358, -23.83943, -23.6345, -23.42879, -23.22229, 
    -23.01501, -22.80694, -22.59808, -22.38843, -22.17799, -21.96675, 
    -21.75471, -21.54188, -21.32825, -21.11381, -20.89857, -20.68252, 
    -20.46566, -20.248, -20.02952, -19.81024, -19.59014, -19.36923, -19.1475, 
    -18.92495, -18.70159, -18.47741, -18.25241, -18.02658, -17.79994, 
    -17.57247, -17.34418, -17.11507, -16.88514, -16.65437, -16.42279, 
    -16.19038, -15.95714, -15.72308, -15.48819, -15.25248, -15.01594, 
    -14.77858, -14.54039, -14.30138, -14.06154, -13.82088, -13.5794, 
    -13.33709, -13.09396, -12.85002, -12.60525, -12.35967, -12.11327, 
    -11.86605, -11.61802, -11.36917, -11.11952, -10.86905, -10.61778, 
    -10.36571, -10.11283, -9.859145, -9.604666, -9.34939, -9.09332, -8.83646, 
    -8.578811, -8.320376, -8.06116, -7.801165, -7.540393, -7.278849, 
    -7.016536, -6.753458, -6.489618, -6.22502, -5.959669, -5.693567, 
    -5.426721, -5.159134, -4.89081, -4.621755, -4.351973, -4.081469, 
    -3.810248, -3.538316, -3.265676, -2.992336, -2.718301, -2.443576, 
    -2.168167, -1.89208, -1.615322, -1.337898, -1.059815, -0.7810791, 
    -0.5016977, -0.221677, 0.05897582, 0.3402538, 0.6221499, 0.9046566, 
    1.187767, 1.471472, 1.755766, 2.04064, 2.326086, 2.612096, 2.898662, 
    3.185776, 3.473429, 3.761612, 4.050317, 4.339536, 4.629258, 4.919476, 
    5.210179, 5.501359, 5.793006, 6.085111, 6.377664, 6.670655, 6.964075, 
    7.257914, 7.55216, 7.846806, 8.141839, 8.43725, 8.733028, 9.029163, 
    9.325645, 9.622462, 9.919603, 10.21706, 10.51482, 10.81287, 11.1112, 
    11.4098, 11.70866, 12.00776, 12.30711, 12.60667, 12.90645, 13.20643, 
    13.5066, 13.80694, 14.10746, 14.40812, 14.70894, 15.00988, 15.31094, 
    15.6121, 15.91336, 16.21471, 16.51612, 16.8176, 17.11912, 17.42068, 
    17.72226, 18.02385, 18.32545, 18.62702, 18.92858, 19.23009, 19.53156, 
    19.83296, 20.1343, 20.43554, 20.73669, 21.03773, 21.33866, 21.63944, 
    21.94009, 22.24058, 22.5409, 22.84104, 23.14098, 23.44073, 23.74026, 
    24.03957, 24.33863, 24.63745, 24.93601, 25.2343, 25.5323, 25.83001, 
    26.12742, 26.42451, 26.72128, 27.0177, 27.31378, 27.6095, 27.90486, 
    28.19983, 28.49441, 28.7886, 29.08237, 29.37572, 29.66864, 29.96112, 
    30.25316, 30.54473, 30.83584, 31.12646, 31.4166, 31.70625, 31.99539, 
    32.28401, 32.57211, 32.85968, 33.14671, 33.43318, 33.7191, 34.00446, 
    34.28924, 34.57344, 34.85706, 35.14007, 35.42248, 35.70428, 35.98546, 
    36.26601, 36.54593, 36.82521, 37.10385, 37.38182, 37.65915, 37.9358, 
    38.21178, 38.48708, 38.7617, 39.03562, 39.30885, 39.58138, 39.8532, 
    40.12431, 40.3947, 40.66436, 40.9333, 41.20151, 41.46898, 41.73571, 
    42.00169, 42.26693, 42.5314, 42.79512, 43.05808, 43.32027, 43.5817, 
    43.84234, 44.10221, 44.36131, 44.61962, 44.87714, 45.13388, 45.38982, 
    45.64497, 45.89933, 46.15288, 46.40563, 46.65758, 46.90873, 47.15906, 
    47.40859, 47.65731, 47.90521, 48.15229, 48.39857, 48.64402, 48.88866, 
    49.13248, 49.37547, 49.61765, 49.859, 50.09953, 50.33924, 50.57812, 
    50.81618, 51.05341, 51.28982, 51.5254, 51.76016, 51.99409, 52.2272, 
    52.45948, 52.69093, 52.92156, 53.15137, 53.38035, 53.60851, 53.83585, 
    54.06236, 54.28805, 54.51292, 54.73698, 54.96021, 55.18262, 55.40422, 
    55.62501, 55.84498, 56.06414, 56.28248, 56.50002, 56.71675, 56.93267, 
    57.14778, 57.36209, 57.5756, 57.78831, 58.00022, 58.21133, 58.42165, 
    58.63117, 58.8399, 59.04785, 59.25501, 59.46138, 59.66697, 59.87178, 
    60.07581, 60.27906, 60.48154, 60.68325, 60.88419, 61.08436, 61.28377, 
    61.48241, 61.6803, 61.87743, 62.0738, 62.26943,
  -41.70105, -41.56259, -41.42366, -41.28423, -41.14433, -41.00393, 
    -40.86304, -40.72165, -40.57977, -40.43738, -40.29449, -40.1511, 
    -40.00719, -39.86277, -39.71784, -39.57238, -39.42641, -39.27991, 
    -39.13289, -38.98533, -38.83725, -38.68863, -38.53946, -38.38976, 
    -38.23951, -38.08871, -37.93737, -37.78547, -37.63301, -37.48, -37.32642, 
    -37.17228, -37.01756, -36.86228, -36.70642, -36.54998, -36.39297, 
    -36.23537, -36.07718, -35.9184, -35.75903, -35.59907, -35.4385, 
    -35.27734, -35.11556, -34.95318, -34.79019, -34.62658, -34.46236, 
    -34.29752, -34.13205, -33.96595, -33.79922, -33.63187, -33.46387, 
    -33.29524, -33.12596, -32.95604, -32.78547, -32.61424, -32.44237, 
    -32.26983, -32.09663, -31.92277, -31.74824, -31.57304, -31.39717, 
    -31.22062, -31.0434, -30.86548, -30.68689, -30.5076, -30.32763, 
    -30.14695, -29.96558, -29.78351, -29.60074, -29.41726, -29.23307, 
    -29.04816, -28.86254, -28.6762, -28.48915, -28.30136, -28.11285, 
    -27.92361, -27.73363, -27.54292, -27.35147, -27.15928, -26.96635, 
    -26.77267, -26.57823, -26.38305, -26.18711, -25.99041, -25.79296, 
    -25.59473, -25.39575, -25.19599, -24.99547, -24.79417, -24.5921, 
    -24.38925, -24.18562, -23.9812, -23.776, -23.57001, -23.36324, -23.15567, 
    -22.94731, -22.73815, -22.5282, -22.31744, -22.10588, -21.89352, 
    -21.68036, -21.46638, -21.2516, -21.03601, -20.8196, -20.60238, 
    -20.38434, -20.16548, -19.94581, -19.72531, -19.50399, -19.28185, 
    -19.05889, -18.8351, -18.61049, -18.38504, -18.15877, -17.93167, 
    -17.70374, -17.47498, -17.24539, -17.01496, -16.7837, -16.55161, 
    -16.31869, -16.08493, -15.85034, -15.61492, -15.37866, -15.14156, 
    -14.90364, -14.66488, -14.42528, -14.18486, -13.9436, -13.70151, 
    -13.45859, -13.21484, -12.97026, -12.72485, -12.47861, -12.23155, 
    -11.98366, -11.73496, -11.48542, -11.23507, -10.9839, -10.73192, 
    -10.47912, -10.2255, -9.971082, -9.715851, -9.459814, -9.202974, 
    -8.945334, -8.686896, -8.427664, -8.16764, -7.906827, -7.645229, 
    -7.38285, -7.119692, -6.855759, -6.591055, -6.325584, -6.05935, 
    -5.792357, -5.524609, -5.256112, -4.986868, -4.716884, -4.446163, 
    -4.174711, -3.902533, -3.629634, -3.356019, -3.081695, -2.806666, 
    -2.530938, -2.254517, -1.97741, -1.699622, -1.421159, -1.142029, 
    -0.8622371, -0.5817907, -0.3006966, -0.01896166, 0.263407, 0.5464021, 
    0.8300163, 1.114242, 1.399072, 1.684498, 1.970512, 2.257106, 2.544272, 
    2.832002, 3.120288, 3.40912, 3.69849, 3.988389, 4.27881, 4.569741, 
    4.861174, 5.1531, 5.44551, 5.738393, 6.031741, 6.325544, 6.619791, 
    6.914473, 7.209579, 7.5051, 7.801025, 8.097344, 8.394047, 8.691122, 
    8.98856, 9.286348, 9.584476, 9.882936, 10.18171, 10.4808, 10.78018, 
    11.07984, 11.37978, 11.67998, 11.98044, 12.28113, 12.58205, 12.88318, 
    13.18452, 13.48605, 13.78776, 14.08964, 14.39168, 14.69386, 14.99618, 
    15.29861, 15.60116, 15.9038, 16.20652, 16.50932, 16.81218, 17.11508, 
    17.41802, 17.72099, 18.02396, 18.32694, 18.6299, 18.93283, 19.23573, 
    19.53858, 19.84137, 20.14408, 20.44671, 20.74924, 21.05165, 21.35395, 
    21.65611, 21.95812, 22.25997, 22.56166, 22.86316, 23.16447, 23.46557, 
    23.76645, 24.06711, 24.36752, 24.66768, 24.96758, 25.2672, 25.56653, 
    25.86557, 26.1643, 26.4627, 26.76078, 27.05851, 27.35589, 27.65291, 
    27.94955, 28.24581, 28.54167, 28.83713, 29.13217, 29.42678, 29.72096, 
    30.01469, 30.30797, 30.60078, 30.89311, 31.18496, 31.47631, 31.76716, 
    32.0575, 32.34732, 32.6366, 32.92535, 33.21355, 33.50119, 33.78827, 
    34.07477, 34.36069, 34.64602, 34.93076, 35.21489, 35.49841, 35.7813, 
    36.06357, 36.3452, 36.6262, 36.90654, 37.18623, 37.46525, 37.74361, 
    38.02129, 38.29829, 38.5746, 38.85022, 39.12513, 39.39935, 39.67285, 
    39.94564, 40.2177, 40.48904, 40.75964, 41.02951, 41.29863, 41.56701, 
    41.83464, 42.10151, 42.36763, 42.63298, 42.89756, 43.16137, 43.4244, 
    43.68666, 43.94814, 44.20882, 44.46872, 44.72783, 44.98614, 45.24366, 
    45.50037, 45.75628, 46.01138, 46.26567, 46.51916, 46.77183, 47.02369, 
    47.27473, 47.52495, 47.77435, 48.02293, 48.27069, 48.51762, 48.76372, 
    49.009, 49.25345, 49.49707, 49.73986, 49.98182, 50.22295, 50.46324, 
    50.7027, 50.94133, 51.17912, 51.41608, 51.65221, 51.8875, 52.12196, 
    52.35559, 52.58838, 52.82034, 53.05147, 53.28176, 53.51122, 53.73985, 
    53.96765, 54.19462, 54.42076, 54.64607, 54.87056, 55.09422, 55.31705, 
    55.53906, 55.76025, 55.98061, 56.20015, 56.41888, 56.63679, 56.85388, 
    57.07016, 57.28563, 57.50028, 57.71413, 57.92717, 58.1394, 58.35083, 
    58.56146, 58.77129, 58.98032, 59.18856, 59.396, 59.60265, 59.80851, 
    60.01359, 60.21788, 60.42139, 60.62411, 60.82607, 61.02724, 61.22764, 
    61.42728, 61.62614, 61.82424, 62.02158, 62.21815, 62.41397,
  -41.84808, -41.70972, -41.57088, -41.43155, -41.29173, -41.15142, 
    -41.01062, -40.86932, -40.72752, -40.58522, -40.44241, -40.2991, 
    -40.15527, -40.01093, -39.86607, -39.72068, -39.57478, -39.42835, 
    -39.28139, -39.13391, -38.98588, -38.83732, -38.68822, -38.53857, 
    -38.38838, -38.23764, -38.08635, -37.93449, -37.78209, -37.62912, 
    -37.47558, -37.32148, -37.1668, -37.01155, -36.85573, -36.69933, 
    -36.54234, -36.38476, -36.2266, -36.06784, -35.90849, -35.74854, 
    -35.58799, -35.42683, -35.26507, -35.10269, -34.9397, -34.77609, 
    -34.61187, -34.44701, -34.28153, -34.11543, -33.94868, -33.7813, 
    -33.61329, -33.44463, -33.27532, -33.10536, -32.93476, -32.76349, 
    -32.59157, -32.41899, -32.24574, -32.07183, -31.89724, -31.72198, 
    -31.54604, -31.36942, -31.19212, -31.01414, -30.83546, -30.65609, 
    -30.47602, -30.29525, -30.11379, -29.93161, -29.74873, -29.56514, 
    -29.38083, -29.19581, -29.01007, -28.8236, -28.6364, -28.44848, 
    -28.25983, -28.07044, -27.88031, -27.68944, -27.49783, -27.30547, 
    -27.11236, -26.9185, -26.72388, -26.52851, -26.33237, -26.13548, 
    -25.93781, -25.73938, -25.54018, -25.3402, -25.13945, -24.93791, 
    -24.7356, -24.5325, -24.32862, -24.12395, -23.91848, -23.71222, 
    -23.50517, -23.29732, -23.08867, -22.87921, -22.66895, -22.45789, 
    -22.24601, -22.03333, -21.81983, -21.60552, -21.39039, -21.17445, 
    -20.95768, -20.74009, -20.52168, -20.30245, -20.08238, -19.8615, 
    -19.63978, -19.41723, -19.19385, -18.96963, -18.74458, -18.5187, 
    -18.29198, -18.06442, -17.83603, -17.6068, -17.37672, -17.14581, 
    -16.91405, -16.68146, -16.44802, -16.21375, -15.97862, -15.74266, 
    -15.50585, -15.26821, -15.02971, -14.79038, -14.55021, -14.30919, 
    -14.06733, -13.82464, -13.5811, -13.33672, -13.09151, -12.84545, 
    -12.59857, -12.35084, -12.10228, -11.85289, -11.60267, -11.35162, 
    -11.09975, -10.84704, -10.59352, -10.33917, -10.084, -9.828013, 
    -9.571212, -9.313599, -9.055176, -8.795945, -8.535911, -8.275075, 
    -8.013441, -7.751013, -7.487793, -7.223785, -6.958993, -6.69342, 
    -6.427071, -6.159949, -5.892059, -5.623404, -5.35399, -5.083821, 
    -4.812901, -4.541235, -4.26883, -3.995688, -3.721816, -3.447219, 
    -3.171903, -2.895873, -2.619136, -2.341696, -2.06356, -1.784734, 
    -1.505226, -1.22504, -0.9441836, -0.662664, -0.3804878, -0.09766206, 
    0.1858061, 0.4699093, 0.7546402, 1.039991, 1.325954, 1.612522, 1.899686, 
    2.187438, 2.475771, 2.764675, 3.054143, 3.344165, 3.634732, 3.925837, 
    4.217469, 4.50962, 4.80228, 5.095441, 5.389091, 5.683223, 5.977826, 
    6.27289, 6.568405, 6.864361, 7.160748, 7.457555, 7.754773, 8.05239, 
    8.350397, 8.648782, 8.947534, 9.246642, 9.546097, 9.845885, 10.146, 
    10.44642, 10.74715, 11.04816, 11.34945, 11.65101, 11.95282, 12.25488, 
    12.55716, 12.85967, 13.16238, 13.46529, 13.76838, 14.07164, 14.37506, 
    14.67863, 14.98233, 15.28616, 15.59009, 15.89413, 16.19825, 16.50244, 
    16.8067, 17.111, 17.41534, 17.7197, 18.02407, 18.32845, 18.63281, 
    18.93714, 19.24144, 19.54568, 19.84986, 20.15397, 20.45799, 20.76191, 
    21.06572, 21.3694, 21.67294, 21.97634, 22.27958, 22.58264, 22.88552, 
    23.1882, 23.49067, 23.79292, 24.09494, 24.39671, 24.69823, 24.99947, 
    25.30044, 25.60112, 25.9015, 26.20156, 26.5013, 26.8007, 27.09975, 
    27.39844, 27.69677, 27.99471, 28.29227, 28.58942, 28.88616, 29.18248, 
    29.47837, 29.77382, 30.06881, 30.36333, 30.65739, 30.95097, 31.24405, 
    31.53663, 31.8287, 32.12025, 32.41127, 32.70175, 32.99168, 33.28106, 
    33.56988, 33.85812, 34.14578, 34.43285, 34.71932, 35.00519, 35.29044, 
    35.57507, 35.85908, 36.14244, 36.42517, 36.70724, 36.98866, 37.26941, 
    37.54948, 37.82888, 38.1076, 38.38563, 38.66296, 38.93958, 39.2155, 
    39.4907, 39.76519, 40.03894, 40.31197, 40.58426, 40.8558, 41.12661, 
    41.39666, 41.66595, 41.93449, 42.20226, 42.46925, 42.73548, 43.00093, 
    43.2656, 43.52948, 43.79258, 44.05488, 44.31639, 44.5771, 44.83701, 
    45.09611, 45.3544, 45.61189, 45.86856, 46.12442, 46.37946, 46.63367, 
    46.88707, 47.13964, 47.39139, 47.64231, 47.8924, 48.14166, 48.39008, 
    48.63767, 48.88443, 49.13035, 49.37543, 49.61968, 49.86308, 50.10565, 
    50.34737, 50.58825, 50.8283, 51.0675, 51.30585, 51.54337, 51.78004, 
    52.01587, 52.25086, 52.485, 52.71831, 52.95077, 53.18239, 53.41317, 
    53.64311, 53.87222, 54.10048, 54.3279, 54.55449, 54.78024, 55.00515, 
    55.22924, 55.45249, 55.6749, 55.89649, 56.11725, 56.33718, 56.55629, 
    56.77457, 56.99202, 57.20866, 57.42448, 57.63948, 57.85366, 58.06703, 
    58.27958, 58.49133, 58.70227, 58.9124, 59.12172, 59.33025, 59.53798, 
    59.7449, 59.95103, 60.15637, 60.36092, 60.56468, 60.76765, 60.96984, 
    61.17125, 61.37188, 61.57174, 61.77082, 61.96913, 62.16667, 62.36345, 
    62.55946,
  -41.99575, -41.85749, -41.71875, -41.57951, -41.43979, -41.29958, 
    -41.15886, -41.01765, -40.87594, -40.73373, -40.591, -40.44777, 
    -40.30402, -40.15976, -40.01498, -39.86967, -39.72384, -39.57749, 
    -39.4306, -39.28318, -39.13522, -38.98673, -38.83769, -38.6881, 
    -38.53797, -38.38729, -38.23605, -38.08425, -37.93189, -37.77897, 
    -37.62548, -37.47142, -37.31679, -37.16158, -37.00579, -36.84942, 
    -36.69247, -36.53492, -36.37679, -36.21805, -36.05872, -35.89879, 
    -35.73825, -35.57711, -35.41536, -35.25299, -35.09, -34.9264, -34.76217, 
    -34.59731, -34.43183, -34.26571, -34.09895, -33.93156, -33.76352, 
    -33.59484, -33.42551, -33.25552, -33.08488, -32.91358, -32.74162, 
    -32.569, -32.3957, -32.22174, -32.0471, -31.87178, -31.69578, -31.51909, 
    -31.34172, -31.16366, -30.9849, -30.80545, -30.6253, -30.44444, 
    -30.26288, -30.08061, -29.89762, -29.71392, -29.5295, -29.34436, 
    -29.1585, -28.97191, -28.78458, -28.59652, -28.40773, -28.21819, 
    -28.02791, -27.83689, -27.64512, -27.45259, -27.25931, -27.06528, 
    -26.87048, -26.67492, -26.47859, -26.2815, -26.08363, -25.88499, 
    -25.68557, -25.48537, -25.2844, -25.08263, -24.88008, -24.67674, 
    -24.4726, -24.26767, -24.06195, -23.85542, -23.64809, -23.43996, 
    -23.23102, -23.02127, -22.81071, -22.59934, -22.38715, -22.17414, 
    -21.96032, -21.74567, -21.5302, -21.3139, -21.09678, -20.87883, 
    -20.66005, -20.44043, -20.21999, -19.9987, -19.77658, -19.55363, 
    -19.32983, -19.10519, -18.87971, -18.65339, -18.42622, -18.19821, 
    -17.96935, -17.73964, -17.50909, -17.27769, -17.04544, -16.81234, 
    -16.57839, -16.34359, -16.10794, -15.87144, -15.63408, -15.39588, 
    -15.15682, -14.91692, -14.67616, -14.43455, -14.19209, -13.94879, 
    -13.70463, -13.45963, -13.21378, -12.96708, -12.71954, -12.47115, 
    -12.22192, -11.97185, -11.72093, -11.46918, -11.2166, -10.96317, 
    -10.70892, -10.45383, -10.19791, -9.941167, -9.683599, -9.425208, 
    -9.165998, -8.905972, -8.64513, -8.383479, -8.12102, -7.857757, 
    -7.593692, -7.32883, -7.063173, -6.796727, -6.529494, -6.261479, 
    -5.992686, -5.723119, -5.452783, -5.181682, -4.909821, -4.637204, 
    -4.363838, -4.089726, -3.814875, -3.539289, -3.262974, -2.985936, 
    -2.708181, -2.429714, -2.150543, -1.870672, -1.590109, -1.308859, 
    -1.02693, -0.7443292, -0.4610623, -0.1771369, 0.1074397, 0.3926601, 
    0.6785169, 0.9650023, 1.252109, 1.539828, 1.828152, 2.117073, 2.406582, 
    2.69667, 2.98733, 3.278553, 3.570328, 3.862649, 4.155505, 4.448887, 
    4.742786, 5.037192, 5.332095, 5.627487, 5.923356, 6.219693, 6.516489, 
    6.813731, 7.111411, 7.409518, 7.708041, 8.006969, 8.306293, 8.606, 
    8.90608, 9.206522, 9.507316, 9.808448, 10.10991, 10.41168, 10.71377, 
    11.01614, 11.3188, 11.62173, 11.92492, 12.22835, 12.53202, 12.83591, 
    13.14001, 13.4443, 13.74879, 14.05345, 14.35827, 14.66324, 14.96834, 
    15.27357, 15.57892, 15.88436, 16.18989, 16.49549, 16.80116, 17.10687, 
    17.41262, 17.7184, 18.02419, 18.32997, 18.63574, 18.94149, 19.2472, 
    19.55285, 19.85845, 20.16396, 20.46939, 20.77472, 21.07993, 21.38501, 
    21.68996, 21.99475, 22.29939, 22.60384, 22.90811, 23.21218, 23.51604, 
    23.81967, 24.12306, 24.42621, 24.72909, 25.03171, 25.33404, 25.63607, 
    25.9378, 26.23921, 26.54029, 26.84103, 27.14141, 27.44143, 27.74108, 
    28.04034, 28.33921, 28.63766, 28.93571, 29.23332, 29.53049, 29.82721, 
    30.12348, 30.41927, 30.71459, 31.00941, 31.30374, 31.59756, 31.89086, 
    32.18363, 32.47586, 32.76755, 33.05869, 33.34925, 33.63925, 33.92867, 
    34.21749, 34.50573, 34.79335, 35.08036, 35.36674, 35.6525, 35.93762, 
    36.22209, 36.50591, 36.78908, 37.07157, 37.35339, 37.63454, 37.91499, 
    38.19475, 38.47381, 38.75216, 39.02981, 39.30673, 39.58293, 39.8584, 
    40.13314, 40.40713, 40.68038, 40.95287, 41.22462, 41.4956, 41.76581, 
    42.03526, 42.30392, 42.57182, 42.83893, 43.10525, 43.37078, 43.63552, 
    43.89945, 44.16259, 44.42492, 44.68644, 44.94716, 45.20705, 45.46614, 
    45.7244, 45.98183, 46.23845, 46.49423, 46.74919, 47.00331, 47.25661, 
    47.50906, 47.76068, 48.01146, 48.2614, 48.51049, 48.75875, 49.00616, 
    49.25272, 49.49844, 49.74331, 49.98733, 50.2305, 50.47283, 50.7143, 
    50.95492, 51.19469, 51.43362, 51.67168, 51.9089, 52.14527, 52.38079, 
    52.61545, 52.84927, 53.08223, 53.31435, 53.54562, 53.77604, 54.00561, 
    54.23433, 54.46221, 54.68924, 54.91543, 55.14078, 55.36528, 55.58895, 
    55.81178, 56.03376, 56.25491, 56.47523, 56.69471, 56.91336, 57.13118, 
    57.34817, 57.56434, 57.77968, 57.99419, 58.20789, 58.42077, 58.63283, 
    58.84407, 59.0545, 59.26412, 59.47293, 59.68094, 59.88814, 60.09454, 
    60.30014, 60.50494, 60.70895, 60.91217, 61.1146, 61.31624, 61.51709, 
    61.71717, 61.91646, 62.11498, 62.31273, 62.5097, 62.70591,
  -42.14407, -42.00591, -41.86726, -41.72813, -41.5885, -41.44838, -41.30777, 
    -41.16665, -41.02503, -40.8829, -40.74026, -40.59711, -40.45345, 
    -40.30927, -40.16457, -40.01935, -39.8736, -39.72732, -39.58051, 
    -39.43316, -39.28527, -39.13684, -38.98787, -38.83835, -38.68828, 
    -38.53766, -38.38647, -38.23473, -38.08243, -37.92956, -37.77612, 
    -37.62211, -37.46752, -37.31236, -37.15661, -37.00028, -36.84336, 
    -36.68584, -36.52774, -36.36903, -36.20973, -36.04982, -35.88931, 
    -35.72818, -35.56644, -35.40408, -35.24111, -35.07751, -34.91328, 
    -34.74843, -34.58294, -34.41681, -34.25005, -34.08264, -33.91459, 
    -33.74588, -33.57653, -33.40652, -33.23585, -33.06452, -32.89252, 
    -32.71986, -32.54652, -32.37251, -32.19781, -32.02244, -31.84638, 
    -31.66964, -31.4922, -31.31407, -31.13523, -30.9557, -30.77547, 
    -30.59453, -30.41287, -30.2305, -30.04742, -29.86362, -29.67909, 
    -29.49384, -29.30785, -29.12114, -28.93369, -28.74549, -28.55656, 
    -28.36688, -28.17646, -27.98528, -27.79335, -27.60067, -27.40722, 
    -27.21301, -27.01803, -26.82229, -26.62577, -26.42849, -26.23042, 
    -26.03157, -25.83194, -25.63153, -25.43032, -25.22833, -25.02554, 
    -24.82196, -24.61758, -24.4124, -24.20641, -23.99962, -23.79202, 
    -23.5836, -23.37438, -23.16434, -22.95348, -22.7418, -22.5293, -22.31597, 
    -22.10182, -21.88684, -21.67103, -21.45438, -21.23691, -21.01859, 
    -20.79944, -20.57945, -20.35862, -20.13694, -19.91442, -19.69106, 
    -19.46685, -19.24179, -19.01587, -18.78911, -18.5615, -18.33303, 
    -18.10371, -17.87354, -17.6425, -17.41061, -17.17787, -16.94426, 
    -16.7098, -16.47448, -16.2383, -16.00126, -15.76336, -15.52459, 
    -15.28497, -15.04449, -14.80315, -14.56095, -14.3179, -14.07398, 
    -13.8292, -13.58357, -13.33708, -13.08974, -12.84154, -12.59249, 
    -12.34258, -12.09182, -11.84022, -11.58776, -11.33446, -11.08032, 
    -10.82533, -10.5695, -10.31283, -10.05532, -9.796985, -9.537814, 
    -9.277813, -9.016987, -8.755336, -8.492865, -8.229576, -7.965473, 
    -7.700559, -7.434838, -7.168313, -6.900988, -6.632866, -6.363953, 
    -6.094252, -5.823767, -5.552502, -5.280464, -5.007655, -4.734082, 
    -4.459748, -4.18466, -3.908822, -3.63224, -3.35492, -3.076867, -2.798087, 
    -2.518586, -2.238371, -1.957447, -1.675821, -1.3935, -1.11049, 
    -0.8267982, -0.5424319, -0.257398, 0.02829606, 0.3146429, 0.601635, 
    0.8892645, 1.177524, 1.466404, 1.755898, 2.045997, 2.336693, 2.627977, 
    2.91984, 3.212274, 3.505269, 3.798816, 4.092907, 4.387532, 4.68268, 
    4.978343, 5.274512, 5.571175, 5.868323, 6.165946, 6.464034, 6.762576, 
    7.061561, 7.36098, 7.66082, 7.961073, 8.261726, 8.56277, 8.864192, 
    9.16598, 9.468125, 9.770616, 10.07344, 10.37658, 10.68004, 10.98379, 
    11.28783, 11.59214, 11.89671, 12.20154, 12.5066, 12.81189, 13.11739, 
    13.4231, 13.72899, 14.03506, 14.34129, 14.64768, 14.9542, 15.26085, 
    15.56762, 15.87448, 16.18144, 16.48846, 16.79556, 17.1027, 17.40988, 
    17.71708, 18.0243, 18.33151, 18.63871, 18.94589, 19.25302, 19.56011, 
    19.86712, 20.17406, 20.48092, 20.78766, 21.09429, 21.40079, 21.70716, 
    22.01337, 22.31941, 22.62527, 22.93094, 23.23641, 23.54167, 23.84669, 
    24.15148, 24.45602, 24.76029, 25.06428, 25.36798, 25.67139, 25.97449, 
    26.27726, 26.57969, 26.88178, 27.18351, 27.48487, 27.78586, 28.08645, 
    28.38664, 28.68641, 28.98576, 29.28468, 29.58315, 29.88116, 30.17871, 
    30.47578, 30.77237, 31.06846, 31.36404, 31.65911, 31.95365, 32.24765, 
    32.54111, 32.83402, 33.12637, 33.41814, 33.70933, 33.99993, 34.28994, 
    34.57933, 34.86811, 35.15628, 35.44381, 35.73069, 36.01694, 36.30253, 
    36.58746, 36.87172, 37.1553, 37.43821, 37.72042, 38.00193, 38.28274, 
    38.56285, 38.84223, 39.1209, 39.39884, 39.67604, 39.9525, 40.22823, 
    40.50319, 40.77741, 41.05086, 41.32355, 41.59546, 41.8666, 42.13697, 
    42.40654, 42.67533, 42.94333, 43.21053, 43.47692, 43.74252, 44.00731, 
    44.27128, 44.53444, 44.79678, 45.0583, 45.319, 45.57887, 45.83791, 
    46.09611, 46.35349, 46.61002, 46.86572, 47.12057, 47.37459, 47.62775, 
    47.88007, 48.13155, 48.38217, 48.63194, 48.88086, 49.12892, 49.37613, 
    49.62248, 49.86798, 50.11262, 50.3564, 50.59932, 50.84138, 51.08259, 
    51.32293, 51.56242, 51.80104, 52.03881, 52.27571, 52.51176, 52.74694, 
    52.98127, 53.21474, 53.44735, 53.6791, 53.91, 54.14004, 54.36923, 
    54.59756, 54.82504, 55.05167, 55.27744, 55.50237, 55.72645, 55.94968, 
    56.17207, 56.39361, 56.6143, 56.83416, 57.05318, 57.27136, 57.48871, 
    57.70522, 57.9209, 58.13575, 58.34977, 58.56297, 58.77534, 58.98689, 
    59.19762, 59.40753, 59.61662, 59.82491, 60.03238, 60.23904, 60.4449, 
    60.64996, 60.85422, 61.05767, 61.26033, 61.4622, 61.66328, 61.86357, 
    62.06308, 62.2618, 62.45974, 62.65691, 62.85331,
  -42.29303, -42.15498, -42.01643, -41.8774, -41.73788, -41.59785, -41.45733, 
    -41.31631, -41.17479, -41.03275, -40.89021, -40.74715, -40.60357, 
    -40.45948, -40.31487, -40.16972, -40.02405, -39.87785, -39.73112, 
    -39.58385, -39.43604, -39.28768, -39.13877, -38.98932, -38.83932, 
    -38.68876, -38.53764, -38.38596, -38.23371, -38.0809, -37.92751, 
    -37.77355, -37.61901, -37.46389, -37.30819, -37.1519, -36.99502, 
    -36.83754, -36.67947, -36.5208, -36.36152, -36.20164, -36.04115, 
    -35.88004, -35.71832, -35.55598, -35.39302, -35.22943, -35.06521, 
    -34.90035, -34.73487, -34.56874, -34.40197, -34.23455, -34.06649, 
    -33.89777, -33.72839, -33.55836, -33.38767, -33.2163, -33.04428, 
    -32.87157, -32.6982, -32.52414, -32.3494, -32.17398, -31.99786, 
    -31.82106, -31.64356, -31.46536, -31.28646, -31.10685, -30.92654, 
    -30.74551, -30.56377, -30.38131, -30.19813, -30.01423, -29.82959, 
    -29.64423, -29.45813, -29.2713, -29.08372, -28.8954, -28.70634, 
    -28.51652, -28.32595, -28.13463, -27.94254, -27.7497, -27.55609, 
    -27.36171, -27.16656, -26.97063, -26.77393, -26.57645, -26.37819, 
    -26.17913, -25.9793, -25.77867, -25.57724, -25.37502, -25.172, -24.96818, 
    -24.76356, -24.55812, -24.35188, -24.14482, -23.93695, -23.72826, 
    -23.51875, -23.30842, -23.09727, -22.88528, -22.67247, -22.45883, 
    -22.24435, -22.02904, -21.81289, -21.5959, -21.37807, -21.1594, 
    -20.93988, -20.71951, -20.49829, -20.27623, -20.05331, -19.82954, 
    -19.60491, -19.37943, -19.15309, -18.92589, -18.69783, -18.46891, 
    -18.23913, -18.00848, -17.77697, -17.54459, -17.31135, -17.07724, 
    -16.84227, -16.60642, -16.36971, -16.13213, -15.89368, -15.65437, 
    -15.41418, -15.17313, -14.9312, -14.68841, -14.44475, -14.20022, 
    -13.95483, -13.70856, -13.46144, -13.21344, -12.96459, -12.71486, 
    -12.46428, -12.21284, -11.96054, -11.70738, -11.45336, -11.19849, 
    -10.94277, -10.68619, -10.42877, -10.1705, -9.911386, -9.65143, 
    -9.390635, -9.129005, -8.866541, -8.603246, -8.339124, -8.074177, 
    -7.808409, -7.541824, -7.274425, -7.006216, -6.737201, -6.467384, 
    -6.196769, -5.92536, -5.653162, -5.38018, -5.106418, -4.831881, 
    -4.556574, -4.280502, -4.003672, -3.726087, -3.447754, -3.168678, 
    -2.888866, -2.608323, -2.327056, -2.045071, -1.762375, -1.478973, 
    -1.194874, -0.9100833, -0.6246088, -0.3384574, -0.05163664, 0.235846, 
    0.5239829, 0.8127661, 1.102188, 1.39224, 1.682914, 1.974202, 2.266095, 
    2.558584, 2.851661, 3.145317, 3.439543, 3.734329, 4.029665, 4.325544, 
    4.621954, 4.918887, 5.216331, 5.514279, 5.812718, 6.111639, 6.411032, 
    6.710885, 7.011189, 7.311933, 7.613105, 7.914695, 8.216692, 8.519084, 
    8.82186, 9.12501, 9.428521, 9.732382, 10.03658, 10.34111, 10.64595, 
    10.95109, 11.25652, 11.56223, 11.86821, 12.17444, 12.48092, 12.78762, 
    13.09454, 13.40166, 13.70898, 14.01648, 14.32414, 14.63195, 14.93991, 
    15.248, 15.5562, 15.8645, 16.17289, 16.48136, 16.7899, 17.09848, 17.4071, 
    17.71575, 18.02441, 18.33307, 18.64172, 18.95033, 19.25891, 19.56744, 
    19.87589, 20.18427, 20.49256, 20.80075, 21.10881, 21.41675, 21.72454, 
    22.03218, 22.33964, 22.64693, 22.95402, 23.26091, 23.56758, 23.87401, 
    24.18021, 24.48614, 24.79181, 25.0972, 25.40229, 25.70709, 26.01156, 
    26.31571, 26.61951, 26.92297, 27.22606, 27.52877, 27.83111, 28.13304, 
    28.43456, 28.73567, 29.03634, 29.33658, 29.63636, 29.93568, 30.23452, 
    30.53288, 30.83075, 31.12812, 31.42497, 31.72129, 32.01709, 32.31234, 
    32.60704, 32.90117, 33.19474, 33.48772, 33.78012, 34.07191, 34.36311, 
    34.65368, 34.94363, 35.23296, 35.52164, 35.80967, 36.09705, 36.38377, 
    36.66981, 36.95518, 37.23986, 37.52385, 37.80714, 38.08973, 38.3716, 
    38.65275, 38.93318, 39.21287, 39.49183, 39.77005, 40.04751, 40.32422, 
    40.60017, 40.87536, 41.14977, 41.42341, 41.69627, 41.96835, 42.23963, 
    42.51012, 42.77981, 43.04869, 43.31678, 43.58405, 43.8505, 44.11614, 
    44.38096, 44.64495, 44.90812, 45.17044, 45.43195, 45.69261, 45.95243, 
    46.21141, 46.46954, 46.72683, 46.98327, 47.23886, 47.4936, 47.74748, 
    48.0005, 48.25267, 48.50398, 48.75443, 49.00401, 49.25273, 49.50058, 
    49.74757, 49.9937, 50.23896, 50.48335, 50.72687, 50.96953, 51.21132, 
    51.45223, 51.69228, 51.93146, 52.16977, 52.40722, 52.64379, 52.87949, 
    53.11433, 53.3483, 53.58141, 53.81365, 54.04502, 54.27553, 54.50518, 
    54.73397, 54.96189, 55.18895, 55.41516, 55.6405, 55.86499, 56.08863, 
    56.31141, 56.53334, 56.75443, 56.97466, 57.19404, 57.41258, 57.63028, 
    57.84714, 58.06315, 58.27833, 58.49268, 58.70619, 58.91887, 59.13072, 
    59.34175, 59.55195, 59.76133, 59.96989, 60.17763, 60.38456, 60.59067, 
    60.79598, 61.00048, 61.20417, 61.40707, 61.60916, 61.81046, 62.01096, 
    62.21067, 62.4096, 62.60774, 62.8051, 63.00167,
  -42.44264, -42.3047, -42.16626, -42.02733, -41.88791, -41.74799, -41.60757, 
    -41.46664, -41.32521, -41.18328, -41.04083, -40.89786, -40.75438, 
    -40.61037, -40.46585, -40.32079, -40.17521, -40.02909, -39.88244, 
    -39.73524, -39.58751, -39.43923, -39.2904, -39.14102, -38.99109, 
    -38.84059, -38.68954, -38.53792, -38.38574, -38.23298, -38.07965, 
    -37.92575, -37.77126, -37.61619, -37.46053, -37.30429, -37.14745, 
    -36.99002, -36.83198, -36.67334, -36.5141, -36.35425, -36.19379, 
    -36.0327, -35.87101, -35.70868, -35.54573, -35.38216, -35.21795, 
    -35.0531, -34.88762, -34.72149, -34.55472, -34.3873, -34.21923, -34.0505, 
    -33.88111, -33.71106, -33.54034, -33.36895, -33.1969, -33.02416, 
    -32.85075, -32.67665, -32.50187, -32.3264, -32.15023, -31.97337, 
    -31.79581, -31.61755, -31.43858, -31.2589, -31.07851, -30.89741, 
    -30.71558, -30.53304, -30.34976, -30.16576, -29.98103, -29.79556, 
    -29.60935, -29.4224, -29.2347, -29.04626, -28.85706, -28.66711, -28.4764, 
    -28.28493, -28.09269, -27.89969, -27.70592, -27.51138, -27.31605, 
    -27.11995, -26.92307, -26.7254, -26.52694, -26.32769, -26.12765, 
    -25.9268, -25.72516, -25.52272, -25.31947, -25.11541, -24.91054, 
    -24.70486, -24.49836, -24.29104, -24.0829, -23.87394, -23.66415, 
    -23.45353, -23.24208, -23.0298, -22.81668, -22.60272, -22.38792, 
    -22.17228, -21.9558, -21.73846, -21.52028, -21.30125, -21.08136, 
    -20.86062, -20.63903, -20.41657, -20.19326, -19.96908, -19.74404, 
    -19.51814, -19.29137, -19.06373, -18.83523, -18.60586, -18.37561, 
    -18.1445, -17.91251, -17.67964, -17.44591, -17.21129, -16.97581, 
    -16.73944, -16.5022, -16.26408, -16.02508, -15.78521, -15.54446, 
    -15.30283, -15.06032, -14.81693, -14.57267, -14.32753, -14.08151, 
    -13.83462, -13.58685, -13.33821, -13.08869, -12.8383, -12.58704, 
    -12.33491, -12.08191, -11.82804, -11.5733, -11.31771, -11.06124, 
    -10.80392, -10.54574, -10.28671, -10.02681, -9.766071, -9.504479, 
    -9.242041, -8.978759, -8.714636, -8.449676, -8.183881, -7.917254, 
    -7.649801, -7.381524, -7.112426, -6.842512, -6.571785, -6.300251, 
    -6.027913, -5.754776, -5.480844, -5.206122, -4.930615, -4.654328, 
    -4.377267, -4.099436, -3.820841, -3.541488, -3.261383, -2.980531, 
    -2.698939, -2.416612, -2.133558, -1.849783, -1.565293, -1.280095, 
    -0.9941969, -0.7076052, -0.4203272, -0.1323706, 0.1562573, 0.4455485, 
    0.7354953, 1.02609, 1.317323, 1.609188, 1.901675, 2.194775, 2.488481, 
    2.782783, 3.077672, 3.373139, 3.669175, 3.96577, 4.262914, 4.560598, 
    4.858811, 5.157545, 5.456789, 5.756531, 6.056763, 6.357473, 6.658651, 
    6.960287, 7.262368, 7.564885, 7.867826, 8.17118, 8.474935, 8.77908, 
    9.083604, 9.388495, 9.693741, 9.999331, 10.30525, 10.61149, 10.91804, 
    11.22488, 11.53201, 11.8394, 12.14706, 12.45496, 12.76309, 13.07144, 
    13.38, 13.68875, 13.99769, 14.3068, 14.61606, 14.92546, 15.235, 15.54465, 
    15.85441, 16.16426, 16.47419, 16.78418, 17.09422, 17.4043, 17.71441, 
    18.02453, 18.33465, 18.64475, 18.95483, 19.26486, 19.57484, 19.88476, 
    20.19459, 20.50434, 20.81397, 21.12349, 21.43287, 21.74211, 22.05119, 
    22.3601, 22.66882, 22.97735, 23.28567, 23.59377, 23.90163, 24.20924, 
    24.51659, 24.82368, 25.13047, 25.43697, 25.74316, 26.04903, 26.35457, 
    26.65976, 26.96459, 27.26906, 27.57314, 27.87683, 28.18012, 28.483, 
    28.78544, 29.08746, 29.38902, 29.69012, 29.99076, 30.29092, 30.59058, 
    30.88974, 31.1884, 31.48653, 31.78413, 32.08118, 32.37769, 32.67364, 
    32.96901, 33.26381, 33.55802, 33.85163, 34.14463, 34.43702, 34.72879, 
    35.01992, 35.31041, 35.60026, 35.88944, 36.17797, 36.46582, 36.75299, 
    37.03947, 37.32526, 37.61034, 37.89472, 38.17838, 38.46132, 38.74353, 
    39.02501, 39.30574, 39.58573, 39.86496, 40.14344, 40.42115, 40.69809, 
    40.97425, 41.24963, 41.52423, 41.79803, 42.07104, 42.34326, 42.61466, 
    42.88526, 43.15505, 43.42402, 43.69216, 43.95948, 44.22598, 44.49164, 
    44.75647, 45.02046, 45.28361, 45.54591, 45.80737, 46.06798, 46.32774, 
    46.58664, 46.84468, 47.10187, 47.3582, 47.61366, 47.86826, 48.12199, 
    48.37485, 48.62684, 48.87796, 49.12822, 49.37759, 49.6261, 49.87373, 
    50.12048, 50.36636, 50.61137, 50.85549, 51.09874, 51.34111, 51.5826, 
    51.82321, 52.06295, 52.3018, 52.53978, 52.77689, 53.01311, 53.24846, 
    53.48294, 53.71654, 53.94926, 54.18111, 54.41209, 54.6422, 54.87143, 
    55.0998, 55.3273, 55.55393, 55.7797, 56.0046, 56.22864, 56.45182, 
    56.67414, 56.8956, 57.1162, 57.33595, 57.55485, 57.7729, 57.9901, 
    58.20645, 58.42196, 58.63662, 58.85045, 59.06343, 59.27559, 59.4869, 
    59.69739, 59.90705, 60.11588, 60.32389, 60.53108, 60.73745, 60.943, 
    61.14774, 61.35167, 61.55479, 61.75711, 61.95863, 62.15934, 62.35926, 
    62.55838, 62.75672, 62.95426, 63.15102,
  -42.5929, -42.45507, -42.31674, -42.17792, -42.0386, -41.89879, -41.75848, 
    -41.61765, -41.47633, -41.33449, -41.19213, -41.04927, -40.90588, 
    -40.76197, -40.61753, -40.47257, -40.32707, -40.18104, -40.03447, 
    -39.88736, -39.73971, -39.59151, -39.44275, -39.29345, -39.14359, 
    -38.99317, -38.84218, -38.69063, -38.53851, -38.38582, -38.23255, 
    -38.0787, -37.92427, -37.76926, -37.61365, -37.45745, -37.30066, 
    -37.14327, -36.98528, -36.82668, -36.66748, -36.50766, -36.34722, 
    -36.18617, -36.0245, -35.8622, -35.69927, -35.53571, -35.37151, 
    -35.20668, -35.0412, -34.87508, -34.70831, -34.54089, -34.37281, 
    -34.20407, -34.03467, -33.8646, -33.69387, -33.52246, -33.35038, 
    -33.17762, -33.00417, -32.83004, -32.65522, -32.4797, -32.30349, 
    -32.12658, -31.94896, -31.77064, -31.59161, -31.41187, -31.2314, 
    -31.05022, -30.86832, -30.68568, -30.50232, -30.31823, -30.13339, 
    -29.94782, -29.7615, -29.57444, -29.38663, -29.19806, -29.00874, 
    -28.81866, -28.62781, -28.4362, -28.24381, -28.05066, -27.85673, 
    -27.66202, -27.46653, -27.27026, -27.07319, -26.87534, -26.67669, 
    -26.47724, -26.27699, -26.07594, -25.87409, -25.67142, -25.46795, 
    -25.26366, -25.05855, -24.85262, -24.64587, -24.4383, -24.22989, 
    -24.02066, -23.81059, -23.59969, -23.38794, -23.17536, -22.96194, 
    -22.74766, -22.53255, -22.31658, -22.09976, -21.88208, -21.66355, 
    -21.44416, -21.22391, -21.0028, -20.78082, -20.55798, -20.33427, 
    -20.10969, -19.88424, -19.65792, -19.43073, -19.20265, -18.97371, 
    -18.74388, -18.51317, -18.28159, -18.04912, -17.81577, -17.58154, 
    -17.34642, -17.11042, -16.87354, -16.63577, -16.39711, -16.15756, 
    -15.91713, -15.67581, -15.43361, -15.19051, -14.94653, -14.70167, 
    -14.45591, -14.20927, -13.96175, -13.71334, -13.46404, -13.21387, 
    -12.9628, -12.71086, -12.45804, -12.20434, -11.94976, -11.69431, 
    -11.43798, -11.18078, -10.9227, -10.66376, -10.40396, -10.14328, 
    -9.88175, -9.619356, -9.356107, -9.092003, -8.827048, -8.561246, 
    -8.294599, -8.02711, -7.758783, -7.489622, -7.219631, -6.948812, 
    -6.677172, -6.404713, -6.13144, -5.857357, -5.582469, -5.306781, 
    -5.030298, -4.753025, -4.474967, -4.196129, -3.916517, -3.636137, 
    -3.354995, -3.073095, -2.790446, -2.507052, -2.22292, -1.938058, 
    -1.652471, -1.366166, -1.079152, -0.7914338, -0.50302, -0.2139181, 
    0.07586446, 0.3663198, 0.65744, 0.9492169, 1.241642, 1.534707, 1.828404, 
    2.122724, 2.417657, 2.713195, 3.009328, 3.306048, 3.603345, 3.901209, 
    4.199631, 4.4986, 4.798108, 5.098143, 5.398695, 5.699754, 6.001309, 
    6.30335, 6.605866, 6.908845, 7.212278, 7.516153, 7.820458, 8.125183, 
    8.430315, 8.735843, 9.041756, 9.348041, 9.654686, 9.96168, 10.26901, 
    10.57667, 10.88463, 11.1929, 11.50145, 11.81028, 12.11937, 12.42871, 
    12.73829, 13.04809, 13.3581, 13.66831, 13.9787, 14.28927, 14.59999, 
    14.91086, 15.22186, 15.53298, 15.84421, 16.15553, 16.46693, 16.77839, 
    17.08991, 17.40147, 17.71305, 18.02464, 18.33624, 18.64782, 18.95937, 
    19.27088, 19.58233, 19.89372, 20.20503, 20.51624, 20.82734, 21.13832, 
    21.44917, 21.75987, 22.07041, 22.38077, 22.69095, 23.00093, 23.3107, 
    23.62024, 23.92954, 24.23859, 24.54737, 24.85588, 25.1641, 25.47202, 
    25.77962, 26.0869, 26.39384, 26.70043, 27.00666, 27.31251, 27.61798, 
    27.92305, 28.22771, 28.53194, 28.83575, 29.13911, 29.44202, 29.74446, 
    30.04642, 30.3479, 30.64888, 30.94935, 31.2493, 31.54873, 31.84761, 
    32.14595, 32.44372, 32.74092, 33.03756, 33.3336, 33.62904, 33.92387, 
    34.21809, 34.51169, 34.80466, 35.09698, 35.38865, 35.67967, 35.97002, 
    36.25969, 36.54869, 36.83699, 37.1246, 37.4115, 37.69769, 37.98317, 
    38.26791, 38.55193, 38.83521, 39.11774, 39.39952, 39.68054, 39.9608, 
    40.24029, 40.519, 40.79694, 41.07409, 41.35044, 41.62601, 41.90076, 
    42.17472, 42.44786, 42.7202, 42.99171, 43.26239, 43.53225, 43.80128, 
    44.06948, 44.33683, 44.60335, 44.86901, 45.13383, 45.3978, 45.66092, 
    45.92318, 46.18457, 46.44511, 46.70478, 46.96358, 47.22152, 47.47858, 
    47.73477, 47.99009, 48.24453, 48.49809, 48.75077, 49.00258, 49.2535, 
    49.50354, 49.75269, 50.00096, 50.24835, 50.49485, 50.74046, 50.98519, 
    51.22903, 51.47198, 51.71404, 51.95522, 52.19551, 52.43492, 52.67344, 
    52.91107, 53.14781, 53.38367, 53.61865, 53.85274, 54.08595, 54.31828, 
    54.54972, 54.78029, 55.00998, 55.23879, 55.46672, 55.69378, 55.91996, 
    56.14528, 56.36972, 56.59329, 56.81599, 57.03783, 57.25881, 57.47892, 
    57.69818, 57.91657, 58.13411, 58.3508, 58.56663, 58.78162, 58.99575, 
    59.20905, 59.42149, 59.6331, 59.84388, 60.05381, 60.26291, 60.47119, 
    60.67863, 60.88525, 61.09105, 61.29603, 61.50019, 61.70354, 61.90607, 
    62.1078, 62.30872, 62.50884, 62.70816, 62.90669, 63.10442, 63.30136,
  -42.74382, -42.6061, -42.46788, -42.32917, -42.18997, -42.05027, -41.91006, 
    -41.76934, -41.62812, -41.48638, -41.34413, -41.20136, -41.05807, 
    -40.91426, -40.76992, -40.62505, -40.47964, -40.3337, -40.18722, 
    -40.0402, -39.89263, -39.74451, -39.59584, -39.44661, -39.29683, 
    -39.14648, -38.99557, -38.84409, -38.69204, -38.53941, -38.38621, 
    -38.23242, -38.07805, -37.92309, -37.76754, -37.6114, -37.45466, 
    -37.29731, -37.13937, -36.98081, -36.82165, -36.66187, -36.50146, 
    -36.34045, -36.1788, -36.01653, -35.85362, -35.69009, -35.52591, 
    -35.36109, -35.19563, -35.02951, -34.86275, -34.69532, -34.52724, 
    -34.35851, -34.1891, -34.01902, -33.84827, -33.67685, -33.50474, 
    -33.33195, -33.15848, -32.98431, -32.80946, -32.6339, -32.45765, 
    -32.28069, -32.10302, -31.92464, -31.74555, -31.56574, -31.38521, 
    -31.20396, -31.02198, -30.83926, -30.65582, -30.47163, -30.2867, 
    -30.10103, -29.91461, -29.72744, -29.53951, -29.35083, -29.16138, 
    -28.97117, -28.78019, -28.58844, -28.39591, -28.20261, -28.00853, 
    -27.81366, -27.618, -27.42156, -27.22432, -27.02628, -26.82744, -26.6278, 
    -26.42736, -26.2261, -26.02403, -25.82115, -25.61745, -25.41293, 
    -25.20759, -25.00142, -24.79442, -24.58659, -24.37792, -24.16842, 
    -23.95807, -23.74689, -23.53485, -23.32198, -23.10825, -22.89367, 
    -22.67823, -22.46194, -22.24478, -22.02677, -21.80789, -21.58815, 
    -21.36753, -21.14605, -20.9237, -20.70047, -20.47637, -20.25139, 
    -20.02553, -19.79879, -19.57117, -19.34266, -19.11327, -18.88299, 
    -18.65183, -18.41977, -18.18683, -17.953, -17.71827, -17.48265, 
    -17.24614, -17.00873, -16.77043, -16.53123, -16.29114, -16.05015, 
    -15.80826, -15.56548, -15.3218, -15.07723, -14.83176, -14.58539, 
    -14.33813, -14.08997, -13.84091, -13.59097, -13.34013, -13.08839, 
    -12.83577, -12.58225, -12.32785, -12.07256, -11.81638, -11.55932, 
    -11.30138, -11.04255, -10.78285, -10.52226, -10.26081, -9.998481, 
    -9.735283, -9.471218, -9.206288, -8.940497, -8.673849, -8.406344, 
    -8.137988, -7.868784, -7.598735, -7.327845, -7.056117, -6.783557, 
    -6.510168, -6.235953, -5.960919, -5.68507, -5.40841, -5.130944, 
    -4.852678, -4.573617, -4.293765, -4.013129, -3.731714, -3.449527, 
    -3.166572, -2.882858, -2.598388, -2.313171, -2.027213, -1.740521, 
    -1.453101, -1.164961, -0.8761073, -0.5865486, -0.2962919, -0.005344956, 
    0.2862843, 0.5785879, 0.8715576, 1.165185, 1.459462, 1.754379, 2.049927, 
    2.346099, 2.642884, 2.940274, 3.238258, 3.536828, 3.835974, 4.135685, 
    4.435953, 4.736765, 5.038114, 5.339987, 5.642375, 5.945267, 6.248652, 
    6.552518, 6.856856, 7.161654, 7.4669, 7.772584, 8.078692, 8.385216, 
    8.692141, 8.999456, 9.30715, 9.61521, 9.923623, 10.23238, 10.54146, 
    10.85087, 11.16057, 11.47057, 11.78084, 12.09139, 12.40218, 12.71322, 
    13.02448, 13.33596, 13.64764, 13.95951, 14.27155, 14.58375, 14.8961, 
    15.20858, 15.52119, 15.8339, 16.14671, 16.45959, 16.77255, 17.08556, 
    17.3986, 17.71168, 18.02476, 18.33785, 18.65092, 18.96396, 19.27696, 
    19.5899, 19.90278, 20.21557, 20.52827, 20.84086, 21.15332, 21.46565, 
    21.77782, 22.08984, 22.40168, 22.71332, 23.02477, 23.336, 23.647, 
    23.95775, 24.26825, 24.57849, 24.88844, 25.1981, 25.50745, 25.81648, 
    26.12519, 26.43354, 26.74155, 27.04918, 27.35644, 27.6633, 27.96976, 
    28.2758, 28.58141, 28.88659, 29.19131, 29.49558, 29.79937, 30.10268, 
    30.40549, 30.7078, 31.00959, 31.31085, 31.61158, 31.91176, 32.21138, 
    32.51044, 32.80892, 33.10681, 33.4041, 33.70079, 33.99686, 34.29232, 
    34.58713, 34.88131, 35.17483, 35.46769, 35.75989, 36.05141, 36.34225, 
    36.6324, 36.92184, 37.21059, 37.49862, 37.78592, 38.07249, 38.35834, 
    38.64344, 38.92779, 39.21138, 39.49422, 39.77628, 40.05757, 40.33809, 
    40.61781, 40.89675, 41.17489, 41.45223, 41.72876, 42.00448, 42.27938, 
    42.55347, 42.82673, 43.09916, 43.37075, 43.64151, 43.91142, 44.1805, 
    44.44872, 44.71608, 44.9826, 45.24825, 45.51305, 45.77697, 46.04004, 
    46.30222, 46.56354, 46.82399, 47.08355, 47.34224, 47.60004, 47.85696, 
    48.113, 48.36815, 48.62241, 48.87579, 49.12827, 49.37986, 49.63056, 
    49.88037, 50.12928, 50.3773, 50.62442, 50.87064, 51.11597, 51.36041, 
    51.60395, 51.84658, 52.08833, 52.32917, 52.56913, 52.80818, 53.04634, 
    53.28361, 53.51998, 53.75546, 53.99004, 54.22374, 54.45654, 54.68845, 
    54.91948, 55.14961, 55.37886, 55.60723, 55.83471, 56.06131, 56.28703, 
    56.51188, 56.73584, 56.95893, 57.18114, 57.40249, 57.62296, 57.84257, 
    58.06131, 58.27919, 58.49621, 58.71236, 58.92767, 59.14211, 59.35571, 
    59.56845, 59.78035, 59.9914, 60.20161, 60.41098, 60.61952, 60.82722, 
    61.03409, 61.24013, 61.44534, 61.64973, 61.8533, 62.05605, 62.25799, 
    62.45912, 62.65944, 62.85895, 63.05766, 63.25557, 63.45269,
  -42.8954, -42.75779, -42.61969, -42.4811, -42.34201, -42.20242, -42.06232, 
    -41.92171, -41.7806, -41.63897, -41.49682, -41.35416, -41.21097, 
    -41.06726, -40.92302, -40.77824, -40.63293, -40.48708, -40.34069, 
    -40.19376, -40.04628, -39.89825, -39.74966, -39.60052, -39.45081, 
    -39.30054, -39.14971, -38.9983, -38.84632, -38.69377, -38.54063, 
    -38.38691, -38.2326, -38.07771, -37.92221, -37.76613, -37.60944, 
    -37.45215, -37.29425, -37.13574, -36.97662, -36.81688, -36.65652, 
    -36.49554, -36.33393, -36.17168, -36.00881, -35.84529, -35.68114, 
    -35.51633, -35.35089, -35.18479, -35.01803, -34.85062, -34.68254, 
    -34.5138, -34.34439, -34.1743, -34.00354, -33.8321, -33.65998, -33.48717, 
    -33.31367, -33.13948, -32.96459, -32.789, -32.61271, -32.4357, -32.25799, 
    -32.07956, -31.90041, -31.72054, -31.53995, -31.35863, -31.17657, 
    -30.99378, -30.81025, -30.62598, -30.44096, -30.2552, -30.06867, 
    -29.8814, -29.69336, -29.50456, -29.315, -29.12466, -28.93355, -28.74167, 
    -28.549, -28.35555, -28.16132, -27.96629, -27.77048, -27.57386, 
    -27.37645, -27.17823, -26.97921, -26.77938, -26.57874, -26.37728, 
    -26.17501, -25.97191, -25.76799, -25.56324, -25.35767, -25.15126, 
    -24.94401, -24.73593, -24.527, -24.31723, -24.10661, -23.89515, 
    -23.68283, -23.46966, -23.25563, -23.04074, -22.82499, -22.60837, 
    -22.39089, -22.17253, -21.95331, -21.73322, -21.51224, -21.29039, 
    -21.06766, -20.84405, -20.61956, -20.39417, -20.16791, -19.94075, 
    -19.7127, -19.48376, -19.25393, -19.02321, -18.79158, -18.55906, 
    -18.32564, -18.09132, -17.8561, -17.61998, -17.38296, -17.14503, 
    -16.9062, -16.66646, -16.42582, -16.18427, -15.94182, -15.69846, 
    -15.4542, -15.20903, -14.96295, -14.71597, -14.46808, -14.21929, 
    -13.96959, -13.71899, -13.46748, -13.21508, -12.96177, -12.70756, 
    -12.45245, -12.19645, -11.93954, -11.68175, -11.42306, -11.16348, 
    -10.903, -10.64165, -10.3794, -10.11628, -9.852271, -9.587388, -9.32163, 
    -9.054998, -8.787498, -8.519134, -8.249906, -7.979819, -7.708876, 
    -7.437082, -7.16444, -6.890954, -6.61663, -6.341469, -6.065478, 
    -5.788661, -5.511022, -5.232567, -4.953301, -4.673229, -4.392357, 
    -4.11069, -3.828233, -3.544993, -3.260976, -2.976188, -2.690635, 
    -2.404325, -2.117262, -1.829456, -1.540911, -1.251637, -0.961639, 
    -0.6709259, -0.3795049, -0.08738377, 0.2054294, 0.4989265, 0.7930992, 
    1.087939, 1.383438, 1.679586, 1.976375, 2.273797, 2.57184, 2.870497, 
    3.169758, 3.469613, 3.770052, 4.071065, 4.372643, 4.674774, 4.977448, 
    5.280656, 5.584386, 5.888628, 6.193369, 6.498601, 6.80431, 7.110487, 
    7.417119, 7.724194, 8.031702, 8.33963, 8.647966, 8.956699, 9.265816, 
    9.575304, 9.885153, 10.19535, 10.50588, 10.81673, 11.12789, 11.43935, 
    11.75109, 12.0631, 12.37536, 12.68788, 13.00062, 13.31358, 13.62674, 
    13.9401, 14.25363, 14.56733, 14.88117, 15.19515, 15.50926, 15.82347, 
    16.13778, 16.45218, 16.76664, 17.08115, 17.39571, 17.71029, 18.02488, 
    18.33948, 18.65405, 18.9686, 19.28311, 19.59756, 19.91194, 20.22623, 
    20.54043, 20.85452, 21.16848, 21.48231, 21.79598, 22.10948, 22.42281, 
    22.73594, 23.04887, 23.36157, 23.67405, 23.98627, 24.29824, 24.60994, 
    24.92135, 25.23246, 25.54326, 25.85374, 26.16388, 26.47367, 26.78311, 
    27.09216, 27.40083, 27.70911, 28.01697, 28.32441, 28.63141, 28.93797, 
    29.24408, 29.54971, 29.85487, 30.15953, 30.46369, 30.76734, 31.07047, 
    31.37305, 31.6751, 31.97659, 32.27751, 32.57786, 32.87762, 33.17678, 
    33.47535, 33.77329, 34.07061, 34.3673, 34.66335, 34.95874, 35.25348, 
    35.54755, 35.84093, 36.13364, 36.42565, 36.71696, 37.00756, 37.29744, 
    37.5866, 37.87503, 38.16272, 38.44967, 38.73586, 39.02129, 39.30595, 
    39.58985, 39.87297, 40.1553, 40.43684, 40.71759, 40.99753, 41.27667, 
    41.55499, 41.8325, 42.10919, 42.38505, 42.66008, 42.93427, 43.20762, 
    43.48013, 43.75179, 44.0226, 44.29255, 44.56164, 44.82987, 45.09723, 
    45.36373, 45.62934, 45.89409, 46.15796, 46.42094, 46.68305, 46.94427, 
    47.2046, 47.46404, 47.72259, 47.98024, 48.237, 48.49287, 48.74783, 
    49.0019, 49.25507, 49.50733, 49.75869, 50.00915, 50.25871, 50.50735, 
    50.7551, 51.00194, 51.24787, 51.4929, 51.73702, 51.98023, 52.22254, 
    52.46395, 52.70444, 52.94404, 53.18272, 53.42051, 53.65739, 53.89337, 
    54.12845, 54.36263, 54.5959, 54.82828, 55.05976, 55.29035, 55.52004, 
    55.74884, 55.97674, 56.20376, 56.42989, 56.65512, 56.87948, 57.10295, 
    57.32554, 57.54726, 57.76809, 57.98805, 58.20713, 58.42535, 58.64269, 
    58.85917, 59.07479, 59.28954, 59.50343, 59.71647, 59.92865, 60.13999, 
    60.35047, 60.5601, 60.7689, 60.97685, 61.18396, 61.39024, 61.59569, 
    61.8003, 62.00409, 62.20706, 62.40921, 62.61053, 62.81105, 63.01075, 
    63.20964, 63.40773, 63.60502,
  -43.04763, -42.91015, -42.77217, -42.63369, -42.49472, -42.35524, 
    -42.21526, -42.07477, -41.93377, -41.79224, -41.65021, -41.50765, 
    -41.36457, -41.22096, -41.07682, -40.93214, -40.78693, -40.64119, 
    -40.49489, -40.34805, -40.20066, -40.05272, -39.90422, -39.75516, 
    -39.60554, -39.45536, -39.3046, -39.15327, -39.00137, -38.84889, 
    -38.69582, -38.54218, -38.38794, -38.2331, -38.07767, -37.92165, 
    -37.76502, -37.60778, -37.44994, -37.29148, -37.1324, -36.97271, 
    -36.81239, -36.65145, -36.48987, -36.32767, -36.16482, -36.00134, 
    -35.8372, -35.67243, -35.507, -35.34091, -35.17417, -35.00677, -34.8387, 
    -34.66996, -34.50055, -34.33046, -34.1597, -33.98825, -33.81611, 
    -33.64328, -33.46976, -33.29555, -33.12063, -32.94501, -32.76868, 
    -32.59163, -32.41388, -32.2354, -32.0562, -31.87628, -31.69562, 
    -31.51423, -31.33211, -31.14925, -30.96564, -30.78129, -30.59618, 
    -30.41032, -30.22371, -30.03633, -29.84818, -29.65928, -29.46959, 
    -29.27914, -29.0879, -28.89589, -28.70308, -28.50949, -28.31511, 
    -28.11993, -27.92396, -27.72718, -27.5296, -27.33121, -27.13201, 
    -26.93199, -26.73115, -26.5295, -26.32702, -26.12371, -25.91957, 
    -25.7146, -25.50879, -25.30215, -25.09466, -24.88632, -24.67714, 
    -24.46711, -24.25622, -24.04448, -23.83188, -23.61841, -23.40409, 
    -23.18889, -22.97283, -22.75589, -22.53808, -22.31939, -22.09982, 
    -21.87938, -21.65805, -21.43583, -21.21273, -20.98873, -20.76385, 
    -20.53807, -20.3114, -20.08382, -19.85535, -19.62598, -19.39571, 
    -19.16454, -18.93246, -18.69947, -18.46557, -18.23077, -17.99506, 
    -17.75843, -17.5209, -17.28245, -17.04309, -16.80281, -16.56162, 
    -16.31952, -16.0765, -15.83257, -15.58772, -15.34195, -15.09527, 
    -14.84767, -14.59916, -14.34973, -14.09938, -13.84813, -13.59596, 
    -13.34287, -13.08888, -12.83397, -12.57816, -12.32144, -12.06381, 
    -11.80527, -11.54583, -11.28549, -11.02425, -10.76212, -10.49908, 
    -10.23516, -9.970338, -9.704632, -9.43804, -9.170565, -8.90221, 
    -8.632979, -8.362875, -8.091901, -7.820061, -7.547358, -7.273796, 
    -6.99938, -6.724113, -6.448, -6.171046, -5.893255, -5.614632, -5.335182, 
    -5.054909, -4.77382, -4.49192, -4.209214, -3.925708, -3.641408, 
    -3.356321, -3.070451, -2.783807, -2.496394, -2.208219, -1.91929, 
    -1.629612, -1.339194, -1.048042, -0.7561651, -0.4635701, -0.170265, 
    0.1237421, 0.4184429, 0.7138292, 1.009892, 1.306624, 1.604014, 1.902055, 
    2.200737, 2.500051, 2.799987, 3.100536, 3.401688, 3.703432, 4.00576, 
    4.30866, 4.612122, 4.916136, 5.220691, 5.525776, 5.831381, 6.137493, 
    6.444103, 6.751198, 7.058767, 7.366798, 7.67528, 7.984201, 8.293549, 
    8.603312, 8.913476, 9.224031, 9.534964, 9.846262, 10.15791, 10.4699, 
    10.78222, 11.09485, 11.40778, 11.721, 12.03449, 12.34825, 12.66225, 
    12.97649, 13.29095, 13.60562, 13.92048, 14.23551, 14.55072, 14.86608, 
    15.18158, 15.4972, 15.81293, 16.12877, 16.44468, 16.76066, 17.0767, 
    17.39278, 17.70888, 18.025, 18.34112, 18.65722, 18.9733, 19.28933, 
    19.6053, 19.9212, 20.23702, 20.55273, 20.86834, 21.18381, 21.49915, 
    21.81433, 22.12934, 22.44417, 22.75881, 23.07323, 23.38743, 23.7014, 
    24.01511, 24.32856, 24.64174, 24.95462, 25.26721, 25.57947, 25.89141, 
    26.203, 26.51425, 26.82512, 27.13561, 27.44571, 27.75541, 28.06469, 
    28.37355, 28.68196, 28.98992, 29.29741, 29.60443, 29.91096, 30.217, 
    30.52252, 30.82752, 31.13199, 31.43592, 31.73929, 32.0421, 32.34434, 
    32.64599, 32.94704, 33.2475, 33.54734, 33.84655, 34.14513, 34.44307, 
    34.74036, 35.03698, 35.33294, 35.62822, 35.92281, 36.21671, 36.5099, 
    36.80238, 37.09415, 37.38518, 37.67548, 37.96504, 38.25385, 38.54191, 
    38.8292, 39.11572, 39.40147, 39.68643, 39.97061, 40.25399, 40.53656, 
    40.81834, 41.0993, 41.37944, 41.65876, 41.93725, 42.21491, 42.49173, 
    42.76771, 43.04284, 43.31713, 43.59055, 43.86312, 44.13482, 44.40566, 
    44.67562, 44.94472, 45.21293, 45.48027, 45.74672, 46.01229, 46.27696, 
    46.54075, 46.80364, 47.06564, 47.32674, 47.58693, 47.84623, 48.10462, 
    48.36211, 48.61869, 48.87436, 49.12912, 49.38297, 49.63591, 49.88793, 
    50.13905, 50.38924, 50.63853, 50.88689, 51.13435, 51.38089, 51.62651, 
    51.87121, 52.11501, 52.35788, 52.59984, 52.84088, 53.08101, 53.32023, 
    53.55853, 53.79593, 54.0324, 54.26797, 54.50263, 54.73638, 54.96923, 
    55.20116, 55.4322, 55.66233, 55.89156, 56.11988, 56.34731, 56.57384, 
    56.79948, 57.02422, 57.24808, 57.47104, 57.69312, 57.91431, 58.13462, 
    58.35404, 58.57259, 58.79026, 59.00706, 59.22299, 59.43805, 59.65224, 
    59.86557, 60.07803, 60.28964, 60.50039, 60.71029, 60.91933, 61.12754, 
    61.33489, 61.5414, 61.74708, 61.95192, 62.15593, 62.3591, 62.56145, 
    62.76298, 62.96368, 63.16357, 63.36264, 63.56091, 63.75836,
  -43.20053, -43.06318, -42.92532, -42.78696, -42.64811, -42.50875, 
    -42.36889, -42.22851, -42.08762, -41.94622, -41.80429, -41.66185, 
    -41.51888, -41.37537, -41.23134, -41.08677, -40.94166, -40.79601, 
    -40.64982, -40.50307, -40.35578, -40.20793, -40.05952, -39.91056, 
    -39.76102, -39.61093, -39.46025, -39.30901, -39.15718, -39.00478, 
    -38.85179, -38.69822, -38.54405, -38.38929, -38.23392, -38.07796, 
    -37.92139, -37.76422, -37.60643, -37.44802, -37.289, -37.12936, 
    -36.96909, -36.80819, -36.64665, -36.48448, -36.32167, -36.15822, 
    -35.99412, -35.82937, -35.66396, -35.4979, -35.33117, -35.16378, 
    -34.99573, -34.827, -34.65759, -34.4875, -34.31673, -34.14528, -33.97313, 
    -33.8003, -33.62676, -33.45252, -33.27758, -33.10193, -32.92556, 
    -32.74849, -32.57069, -32.39217, -32.21292, -32.03295, -31.85224, 
    -31.67079, -31.4886, -31.30567, -31.12199, -30.93755, -30.75237, 
    -30.56642, -30.37971, -30.19223, -30.00399, -29.81497, -29.62518, 
    -29.43461, -29.24325, -29.05111, -28.85817, -28.66444, -28.46992, 
    -28.27459, -28.07846, -27.88152, -27.68377, -27.48521, -27.28583, 
    -27.08563, -26.88461, -26.68276, -26.48007, -26.27656, -26.07221, 
    -25.86702, -25.66098, -25.4541, -25.24637, -25.03779, -24.82836, 
    -24.61806, -24.40691, -24.19489, -23.98201, -23.76826, -23.55363, 
    -23.33813, -23.12176, -22.90451, -22.68637, -22.46735, -22.24744, 
    -22.02665, -21.80496, -21.58238, -21.35891, -21.13453, -20.90926, 
    -20.68308, -20.456, -20.22802, -19.99913, -19.76933, -19.53862, 
    -19.30699, -19.07446, -18.841, -18.60663, -18.37135, -18.13514, 
    -17.89802, -17.65997, -17.42101, -17.18111, -16.9403, -16.69856, 
    -16.4559, -16.21232, -15.9678, -15.72237, -15.476, -15.22871, -14.9805, 
    -14.73136, -14.4813, -14.23031, -13.97839, -13.72556, -13.4718, 
    -13.21711, -12.96151, -12.70499, -12.44755, -12.18919, -11.92991, 
    -11.66972, -11.40862, -11.14661, -10.88369, -10.61986, -10.35513, 
    -10.0895, -9.822964, -9.555535, -9.287212, -9.017999, -8.747898, 
    -8.476912, -8.205047, -7.932303, -7.658686, -7.3842, -7.108848, 
    -6.832634, -6.555563, -6.27764, -5.998868, -5.719254, -5.438802, 
    -5.157516, -4.875403, -4.592468, -4.308716, -4.024153, -3.738786, 
    -3.45262, -3.165662, -2.877917, -2.589394, -2.300098, -2.010036, 
    -1.719216, -1.427645, -1.135331, -0.8422799, -0.5485011, -0.254002, 
    0.04120917, 0.3371241, 0.6337345, 0.9310315, 1.229007, 1.52765, 1.826954, 
    2.126909, 2.427504, 2.728731, 3.030581, 3.333041, 3.636104, 3.939758, 
    4.243994, 4.5488, 4.854167, 5.160082, 5.466536, 5.773517, 6.081014, 
    6.389015, 6.697509, 7.006485, 7.31593, 7.625834, 7.936182, 8.246964, 
    8.558167, 8.86978, 9.181788, 9.49418, 9.806943, 10.12006, 10.43353, 
    10.74733, 11.06144, 11.37587, 11.69058, 12.00558, 12.32083, 12.63635, 
    12.9521, 13.26807, 13.58425, 13.90063, 14.2172, 14.53393, 14.85082, 
    15.16785, 15.48501, 15.80228, 16.11964, 16.4371, 16.75462, 17.0722, 
    17.38982, 17.70746, 18.02512, 18.34278, 18.66043, 18.97804, 19.29561, 
    19.61312, 19.93056, 20.24792, 20.56517, 20.88231, 21.19932, 21.51618, 
    21.83289, 22.14942, 22.46577, 22.78193, 23.09787, 23.41358, 23.72905, 
    24.04427, 24.35922, 24.67389, 24.98826, 25.30233, 25.61608, 25.92949, 
    26.24256, 26.55526, 26.86759, 27.17954, 27.49109, 27.80223, 28.11294, 
    28.42322, 28.73305, 29.04242, 29.35132, 29.65974, 29.96766, 30.27508, 
    30.58198, 30.88835, 31.19417, 31.49945, 31.80417, 32.10831, 32.41188, 
    32.71484, 33.01721, 33.31896, 33.62009, 33.92058, 34.22043, 34.51963, 
    34.81817, 35.11604, 35.41323, 35.70973, 36.00554, 36.30064, 36.59502, 
    36.88868, 37.18162, 37.47382, 37.76527, 38.05597, 38.34591, 38.63509, 
    38.92348, 39.21111, 39.49794, 39.78398, 40.06922, 40.35365, 40.63728, 
    40.92008, 41.20206, 41.48322, 41.76354, 42.04302, 42.32166, 42.59945, 
    42.87638, 43.15246, 43.42768, 43.70203, 43.97551, 44.24811, 44.51984, 
    44.79068, 45.06064, 45.32972, 45.5979, 45.86518, 46.13158, 46.39706, 
    46.66166, 46.92534, 47.18811, 47.44999, 47.71094, 47.97099, 48.23011, 
    48.48833, 48.74562, 49.002, 49.25746, 49.512, 49.76561, 50.0183, 
    50.27007, 50.52091, 50.77083, 51.01982, 51.26789, 51.51503, 51.76125, 
    52.00654, 52.25091, 52.49435, 52.73687, 52.97845, 53.21912, 53.45887, 
    53.69769, 53.93559, 54.17257, 54.40863, 54.64377, 54.87799, 55.1113, 
    55.34369, 55.57517, 55.80574, 56.0354, 56.26414, 56.49199, 56.71892, 
    56.94495, 57.17008, 57.39431, 57.61765, 57.84009, 58.06163, 58.28229, 
    58.50206, 58.72094, 58.93893, 59.15604, 59.37228, 59.58764, 59.80213, 
    60.01574, 60.22849, 60.44037, 60.65139, 60.86154, 61.07084, 61.27929, 
    61.48688, 61.69363, 61.89953, 62.10459, 62.30881, 62.51219, 62.71474, 
    62.91646, 63.11736, 63.31742, 63.51667, 63.71511, 63.91273,
  -43.3541, -43.21687, -43.07914, -42.94091, -42.80219, -42.66295, -42.52321, 
    -42.38295, -42.24218, -42.10089, -41.95908, -41.81675, -41.67389, 
    -41.5305, -41.38658, -41.24212, -41.09711, -40.95157, -40.80548, 
    -40.65884, -40.51164, -40.36389, -40.21558, -40.0667, -39.91727, 
    -39.76725, -39.61667, -39.46551, -39.31377, -39.16145, -39.00854, 
    -38.85504, -38.70095, -38.54626, -38.39097, -38.23507, -38.07857, 
    -37.92146, -37.76373, -37.60538, -37.44642, -37.28683, -37.12661, 
    -36.96575, -36.80426, -36.64214, -36.47937, -36.31595, -36.15188, 
    -35.98716, -35.82178, -35.65575, -35.48904, -35.32167, -35.15363, 
    -34.98491, -34.81551, -34.64543, -34.47467, -34.30321, -34.13106, 
    -33.95821, -33.78466, -33.61041, -33.43544, -33.25977, -33.08338, 
    -32.90627, -32.72844, -32.54988, -32.37059, -32.19056, -32.0098, 
    -31.82829, -31.64605, -31.46305, -31.2793, -31.09479, -30.90952, 
    -30.72349, -30.5367, -30.34913, -30.16079, -29.97166, -29.78176, 
    -29.59108, -29.3996, -29.20733, -29.01427, -28.82041, -28.62574, 
    -28.43027, -28.23399, -28.0369, -27.83899, -27.64025, -27.4407, 
    -27.24032, -27.03911, -26.83707, -26.63419, -26.43047, -26.22591, 
    -26.0205, -25.81424, -25.60713, -25.39916, -25.19034, -24.98065, 
    -24.7701, -24.55868, -24.3464, -24.13323, -23.9192, -23.70428, -23.48848, 
    -23.2718, -23.05423, -22.83577, -22.61642, -22.39618, -22.17504, -21.953, 
    -21.73005, -21.50621, -21.28146, -21.0558, -20.82923, -20.60174, 
    -20.37335, -20.14404, -19.91381, -19.68266, -19.45059, -19.2176, 
    -18.98368, -18.74884, -18.51307, -18.27637, -18.03875, -17.80019, 
    -17.56071, -17.32029, -17.07894, -16.83665, -16.59343, -16.34928, 
    -16.10419, -15.85817, -15.61121, -15.36331, -15.11448, -14.86471, 
    -14.61401, -14.36237, -14.1098, -13.8563, -13.60186, -13.34649, 
    -13.09018, -12.83295, -12.57479, -12.3157, -12.05568, -11.79474, 
    -11.53287, -11.27008, -11.00638, -10.74175, -10.47621, -10.20976, 
    -9.9424, -9.674129, -9.404955, -9.134879, -8.863903, -8.592032, -8.31927, 
    -8.045619, -7.771083, -7.495666, -7.219373, -6.942206, -6.664172, 
    -6.385273, -6.105515, -5.824904, -5.543443, -5.261137, -4.977993, 
    -4.694016, -4.409211, -4.123584, -3.837141, -3.549889, -3.261833, 
    -2.972981, -2.683338, -2.392912, -2.10171, -1.809738, -1.517005, 
    -1.223518, -0.929284, -0.6343115, -0.3386083, -0.04218278, 0.2549568, 
    0.5528019, 0.8513438, 1.150573, 1.450482, 1.75106, 2.052299, 2.354188, 
    2.656718, 2.959879, 3.263662, 3.568055, 3.873049, 4.178633, 4.484796, 
    4.791528, 5.098817, 5.406653, 5.715024, 6.02392, 6.333327, 6.643235, 
    6.953632, 7.264506, 7.575845, 7.887636, 8.199868, 8.512527, 8.825602, 
    9.139079, 9.452946, 9.767189, 10.0818, 10.39675, 10.71205, 11.02767, 
    11.3436, 11.65982, 11.97633, 12.29311, 12.61015, 12.92743, 13.24493, 
    13.56265, 13.88057, 14.19868, 14.51696, 14.83539, 15.15397, 15.47268, 
    15.7915, 16.11042, 16.42943, 16.74851, 17.06764, 17.38682, 17.70603, 
    18.02525, 18.34447, 18.66367, 18.98284, 19.30197, 19.62104, 19.94003, 
    20.25894, 20.57775, 20.89643, 21.21499, 21.5334, 21.85165, 22.16973, 
    22.48762, 22.80531, 23.12278, 23.44002, 23.75701, 24.07375, 24.39022, 
    24.7064, 25.02228, 25.33785, 25.65309, 25.96799, 26.28254, 26.59673, 
    26.91053, 27.22395, 27.53696, 27.84955, 28.16171, 28.47343, 28.7847, 
    29.0955, 29.40582, 29.71565, 30.02498, 30.33379, 30.64208, 30.94983, 
    31.25703, 31.56367, 31.86975, 32.17524, 32.48014, 32.78443, 33.08812, 
    33.39118, 33.69361, 33.9954, 34.29653, 34.597, 34.8968, 35.19593, 
    35.49436, 35.79209, 36.08912, 36.38543, 36.68102, 36.97588, 37.26999, 
    37.56336, 37.85597, 38.14782, 38.4389, 38.72921, 39.01873, 39.30745, 
    39.59538, 39.88251, 40.16882, 40.45432, 40.73899, 41.02284, 41.30585, 
    41.58802, 41.86935, 42.14983, 42.42945, 42.70821, 42.98611, 43.26313, 
    43.53929, 43.81457, 44.08897, 44.36248, 44.6351, 44.90683, 45.17766, 
    45.44759, 45.71663, 45.98475, 46.25197, 46.51828, 46.78367, 47.04815, 
    47.31171, 47.57436, 47.83607, 48.09687, 48.35674, 48.61568, 48.8737, 
    49.13079, 49.38694, 49.64217, 49.89646, 50.14981, 50.40224, 50.65373, 
    50.90428, 51.1539, 51.40258, 51.65033, 51.89714, 52.14302, 52.38796, 
    52.63197, 52.87504, 53.11718, 53.35838, 53.59865, 53.83799, 54.0764, 
    54.31388, 54.55043, 54.78605, 55.02074, 55.25451, 55.48736, 55.71928, 
    55.95029, 56.18037, 56.40954, 56.63779, 56.86513, 57.09155, 57.31707, 
    57.54168, 57.76538, 57.98818, 58.21008, 58.43108, 58.65118, 58.87039, 
    59.08871, 59.30613, 59.52268, 59.73833, 59.95311, 60.16701, 60.38004, 
    60.59219, 60.80347, 61.01388, 61.22343, 61.43212, 61.63995, 61.84692, 
    62.05305, 62.25832, 62.46275, 62.66634, 62.86908, 63.071, 63.27207, 
    63.47232, 63.67175, 63.87035, 64.06813,
  -43.50834, -43.37124, -43.23365, -43.09555, -42.95695, -42.81784, 
    -42.67822, -42.53809, -42.39744, -42.25627, -42.11458, -41.97237, 
    -41.82962, -41.68635, -41.54254, -41.39819, -41.2533, -41.10786, 
    -40.96188, -40.81534, -40.66825, -40.5206, -40.37239, -40.22361, 
    -40.07426, -39.92435, -39.77386, -39.62279, -39.47113, -39.3189, 
    -39.16607, -39.01265, -38.85864, -38.70403, -38.54881, -38.39299, 
    -38.23656, -38.07951, -37.92185, -37.76357, -37.60466, -37.44513, 
    -37.28496, -37.12416, -36.96272, -36.80064, -36.63791, -36.47454, 
    -36.3105, -36.14582, -35.98048, -35.81446, -35.64779, -35.48044, 
    -35.31242, -35.14371, -34.97433, -34.80426, -34.6335, -34.46204, 
    -34.28989, -34.11704, -33.94348, -33.76921, -33.59423, -33.41854, 
    -33.24213, -33.06499, -32.88713, -32.70853, -32.5292, -32.34913, 
    -32.16832, -31.98676, -31.80446, -31.6214, -31.43758, -31.253, -31.06766, 
    -30.88155, -30.69467, -30.50701, -30.31858, -30.12936, -29.93935, 
    -29.74856, -29.55697, -29.36458, -29.17139, -28.9774, -28.7826, 
    -28.58698, -28.39056, -28.19331, -27.99524, -27.79635, -27.59662, 
    -27.39607, -27.19467, -26.99244, -26.78937, -26.58545, -26.38068, 
    -26.17505, -25.96858, -25.76124, -25.55304, -25.34398, -25.13404, 
    -24.92324, -24.71156, -24.499, -24.28557, -24.07125, -23.85604, 
    -23.63994, -23.42296, -23.20508, -22.9863, -22.76662, -22.54604, 
    -22.32455, -22.10216, -21.87886, -21.65465, -21.42952, -21.20348, 
    -20.97651, -20.74863, -20.51982, -20.29009, -20.05944, -19.82785, 
    -19.59534, -19.36189, -19.12751, -18.8922, -18.65595, -18.41877, 
    -18.18064, -17.94158, -17.70157, -17.46062, -17.21873, -16.9759, 
    -16.73213, -16.4874, -16.24174, -15.99513, -15.74757, -15.49907, 
    -15.24962, -14.99922, -14.74788, -14.4956, -14.24237, -13.98819, 
    -13.73307, -13.47701, -13.22001, -12.96206, -12.70318, -12.44335, 
    -12.18259, -11.92089, -11.65826, -11.39469, -11.1302, -10.86477, 
    -10.59842, -10.33115, -10.06295, -9.79384, -9.523809, -9.252866, 
    -8.981011, -8.708251, -8.434587, -8.160024, -7.884563, -7.608211, 
    -7.33097, -7.052846, -6.773841, -6.493962, -6.213212, -5.931596, 
    -5.64912, -5.365788, -5.081606, -4.796579, -4.510714, -4.224015, 
    -3.936489, -3.648142, -3.358981, -3.069012, -2.778241, -2.486677, 
    -2.194325, -1.901193, -1.607288, -1.312618, -1.017192, -0.7210153, 
    -0.4240979, -0.1264475, 0.1719273, 0.4710179, 0.7708156, 1.071311, 
    1.372496, 1.67436, 1.976894, 2.280089, 2.583934, 2.88842, 3.193537, 
    3.499273, 3.805619, 4.112565, 4.420098, 4.728209, 5.036886, 5.346118, 
    5.655894, 5.966202, 6.27703, 6.588366, 6.900199, 7.212516, 7.525305, 
    7.838554, 8.15225, 8.466381, 8.780933, 9.095895, 9.411252, 9.726993, 
    10.0431, 10.35957, 10.67638, 10.99351, 11.31097, 11.62872, 11.94676, 
    12.26508, 12.58366, 12.90248, 13.22153, 13.54081, 13.86028, 14.17995, 
    14.49979, 14.81979, 15.13993, 15.46021, 15.7806, 16.10109, 16.42167, 
    16.74233, 17.06304, 17.38379, 17.70458, 18.02537, 18.34617, 18.66695, 
    18.9877, 19.3084, 19.62904, 19.94961, 20.27009, 20.59047, 20.91072, 
    21.23084, 21.55082, 21.87063, 22.19027, 22.50971, 22.82895, 23.14797, 
    23.46675, 23.78529, 24.10356, 24.42156, 24.73927, 25.05667, 25.37376, 
    25.69052, 26.00693, 26.32298, 26.63866, 26.95395, 27.26885, 27.58334, 
    27.8974, 28.21103, 28.5242, 28.83692, 29.14916, 29.46091, 29.77217, 
    30.08292, 30.39314, 30.70283, 31.01198, 31.32057, 31.62859, 31.93603, 
    32.24288, 32.54913, 32.85477, 33.15979, 33.46417, 33.76791, 34.07101, 
    34.37344, 34.67519, 34.97627, 35.27665, 35.57634, 35.87532, 36.17358, 
    36.47112, 36.76791, 37.06397, 37.35928, 37.65383, 37.94761, 38.24062, 
    38.53285, 38.82429, 39.11493, 39.40477, 39.69381, 39.98203, 40.26942, 
    40.55599, 40.84172, 41.12661, 41.41066, 41.69386, 41.9762, 42.25768, 
    42.53829, 42.81804, 43.0969, 43.37489, 43.65199, 43.9282, 44.20351, 
    44.47794, 44.75146, 45.02407, 45.29578, 45.56659, 45.83647, 46.10544, 
    46.37349, 46.64062, 46.90682, 47.1721, 47.43645, 47.69986, 47.96235, 
    48.2239, 48.48451, 48.74419, 49.00293, 49.26072, 49.51758, 49.77349, 
    50.02846, 50.28249, 50.53557, 50.7877, 51.03889, 51.28914, 51.53844, 
    51.78679, 52.0342, 52.28066, 52.52618, 52.77075, 53.01438, 53.25706, 
    53.4988, 53.7396, 53.97945, 54.21837, 54.45635, 54.69339, 54.92949, 
    55.16465, 55.39888, 55.63218, 55.86455, 56.09599, 56.3265, 56.55608, 
    56.78474, 57.01247, 57.23929, 57.46519, 57.69017, 57.91425, 58.1374, 
    58.35965, 58.58099, 58.80143, 59.02097, 59.2396, 59.45734, 59.67419, 
    59.89014, 60.10521, 60.31939, 60.53268, 60.7451, 60.95664, 61.16731, 
    61.37711, 61.58603, 61.79409, 62.0013, 62.20764, 62.41312, 62.61776, 
    62.82155, 63.02449, 63.22659, 63.42785, 63.62827, 63.82786, 64.02663, 
    64.22456,
  -43.66326, -43.52629, -43.38883, -43.25087, -43.1124, -42.97342, -42.83393, 
    -42.69392, -42.5534, -42.41236, -42.27079, -42.1287, -41.98608, 
    -41.84292, -41.69922, -41.55499, -41.41021, -41.26489, -41.11901, 
    -40.97258, -40.8256, -40.67805, -40.52995, -40.38128, -40.23203, 
    -40.08221, -39.93182, -39.78084, -39.62928, -39.47713, -39.32439, 
    -39.17106, -39.01713, -38.8626, -38.70746, -38.55171, -38.39536, 
    -38.23838, -38.08079, -37.92257, -37.76373, -37.60426, -37.44415, 
    -37.28341, -37.12202, -36.95999, -36.79731, -36.63398, -36.46999, 
    -36.30535, -36.14004, -35.97406, -35.80741, -35.64009, -35.47209, 
    -35.30341, -35.13404, -34.96398, -34.79323, -34.62178, -34.44963, 
    -34.27678, -34.10322, -33.92895, -33.75396, -33.57825, -33.40181, 
    -33.22466, -33.04676, -32.86813, -32.68877, -32.50866, -32.3278, 
    -32.1462, -31.96384, -31.78073, -31.59685, -31.4122, -31.22679, 
    -31.04061, -30.85365, -30.6659, -30.47738, -30.28806, -30.09796, 
    -29.90705, -29.71535, -29.52285, -29.32954, -29.13542, -28.94049, 
    -28.74474, -28.54817, -28.35077, -28.15255, -27.9535, -27.7536, 
    -27.55288, -27.35131, -27.14889, -26.94562, -26.74151, -26.53653, 
    -26.3307, -26.12401, -25.91644, -25.70802, -25.49871, -25.28854, 
    -25.07748, -24.86555, -24.65272, -24.43901, -24.22441, -24.00892, 
    -23.79253, -23.57524, -23.35705, -23.13796, -22.91795, -22.69704, 
    -22.47521, -22.25247, -22.02881, -21.80424, -21.57873, -21.35231, 
    -21.12496, -20.89667, -20.66746, -20.43731, -20.20623, -19.97421, 
    -19.74125, -19.50736, -19.27252, -19.03673, -18.8, -18.56233, -18.32371, 
    -18.08413, -17.84361, -17.60213, -17.35971, -17.11633, -16.872, 
    -16.62671, -16.38046, -16.13327, -15.88511, -15.636, -15.38593, 
    -15.13491, -14.88293, -14.63, -14.37611, -14.12126, -13.86546, -13.60871, 
    -13.351, -13.09234, -12.83273, -12.57217, -12.31066, -12.0482, -11.7848, 
    -11.52046, -11.25517, -10.98894, -10.72178, -10.45368, -10.18464, 
    -9.914681, -9.64379, -9.371975, -9.099238, -8.825583, -8.551013, 
    -8.275532, -7.999143, -7.721849, -7.443657, -7.164568, -6.884588, 
    -6.603722, -6.321973, -6.039347, -5.755848, -5.471483, -5.186256, 
    -4.900173, -4.613239, -4.325461, -4.036844, -3.747395, -3.45712, 
    -3.166026, -2.874119, -2.581407, -2.287896, -1.993594, -1.698508, 
    -1.402647, -1.106017, -0.8086268, -0.5104848, -0.2115991, 0.0880217, 
    0.3883688, 0.6894334, 0.9912064, 1.293679, 1.59684, 1.900682, 2.205195, 
    2.510368, 2.816191, 3.122654, 3.429747, 3.737458, 4.045779, 4.354696, 
    4.664199, 4.974278, 5.28492, 5.596114, 5.907849, 6.220111, 6.532891, 
    6.846174, 7.15995, 7.474205, 7.788927, 8.104103, 8.419721, 8.735767, 
    9.052229, 9.369093, 9.686345, 10.00397, 10.32196, 10.6403, 10.95897, 
    11.27797, 11.59727, 11.91686, 12.23673, 12.55687, 12.87725, 13.19787, 
    13.51871, 13.83976, 14.161, 14.48242, 14.804, 15.12573, 15.44759, 
    15.76957, 16.09166, 16.41383, 16.73608, 17.05838, 17.38073, 17.70311, 
    18.0255, 18.34789, 18.67026, 18.99261, 19.3149, 19.63714, 19.9593, 
    20.28136, 20.60333, 20.92517, 21.24688, 21.56843, 21.88982, 22.21103, 
    22.53205, 22.85286, 23.17344, 23.49379, 23.81388, 24.13371, 24.45326, 
    24.77251, 25.09146, 25.41008, 25.72836, 26.0463, 26.36386, 26.68106, 
    26.99786, 27.31425, 27.63023, 27.94578, 28.26089, 28.57554, 28.88972, 
    29.20341, 29.51662, 29.82932, 30.1415, 30.45315, 30.76426, 31.07481, 
    31.3848, 31.69421, 32.00303, 32.31126, 32.61887, 32.92587, 33.23223, 
    33.53795, 33.84302, 34.14743, 34.45116, 34.75422, 35.05658, 35.35824, 
    35.65919, 35.95942, 36.25893, 36.5577, 36.85572, 37.15299, 37.4495, 
    37.74524, 38.0402, 38.33438, 38.62776, 38.92035, 39.21213, 39.50309, 
    39.79324, 40.08255, 40.37104, 40.65868, 40.94548, 41.23143, 41.51652, 
    41.80075, 42.08411, 42.3666, 42.64821, 42.92894, 43.20877, 43.48772, 
    43.76577, 44.04292, 44.31917, 44.59451, 44.86893, 45.14244, 45.41503, 
    45.6867, 45.95745, 46.22726, 46.49615, 46.7641, 47.03112, 47.2972, 
    47.56233, 47.82653, 48.08978, 48.35209, 48.61345, 48.87386, 49.13332, 
    49.39183, 49.64938, 49.90599, 50.16164, 50.41633, 50.67007, 50.92286, 
    51.17468, 51.42556, 51.67547, 51.92443, 52.17243, 52.41948, 52.66557, 
    52.91071, 53.15489, 53.39812, 53.6404, 53.88172, 54.12209, 54.36152, 
    54.59999, 54.83751, 55.07409, 55.30973, 55.54442, 55.77817, 56.01098, 
    56.24285, 56.47378, 56.70378, 56.93285, 57.16098, 57.38819, 57.61447, 
    57.83982, 58.06425, 58.28777, 58.51036, 58.73204, 58.95282, 59.17268, 
    59.39163, 59.60968, 59.82682, 60.04307, 60.25842, 60.47288, 60.68645, 
    60.89913, 61.11093, 61.32184, 61.53188, 61.74104, 61.94934, 62.15676, 
    62.36332, 62.56901, 62.77385, 62.97783, 63.18097, 63.38325, 63.58468, 
    63.78528, 63.98504, 64.18396, 64.38205,
  -43.81886, -43.68203, -43.5447, -43.40687, -43.26854, -43.12969, -42.99033, 
    -42.85046, -42.71007, -42.56915, -42.42772, -42.28575, -42.14325, 
    -42.00021, -41.85664, -41.71252, -41.56786, -41.42266, -41.2769, 
    -41.13058, -40.98371, -40.83627, -40.68827, -40.5397, -40.39056, 
    -40.24084, -40.09055, -39.93967, -39.78821, -39.63615, -39.48351, 
    -39.33027, -39.17642, -39.02197, -38.86692, -38.71125, -38.55497, 
    -38.39808, -38.24055, -38.08241, -37.92363, -37.76423, -37.60418, 
    -37.4435, -37.28217, -37.12019, -36.95757, -36.79428, -36.63034, 
    -36.46574, -36.30047, -36.13453, -35.96792, -35.80063, -35.63266, 
    -35.464, -35.29465, -35.12461, -34.95388, -34.78244, -34.6103, -34.43745, 
    -34.26389, -34.08961, -33.91462, -33.7389, -33.56245, -33.38527, 
    -33.20735, -33.0287, -32.8493, -32.66916, -32.48827, -32.30661, 
    -32.12421, -31.94104, -31.7571, -31.5724, -31.38692, -31.20066, 
    -31.01362, -30.8258, -30.63719, -30.44778, -30.25758, -30.06658, 
    -29.87477, -29.68216, -29.48873, -29.29449, -29.09943, -28.90355, 
    -28.70684, -28.5093, -28.31092, -28.11171, -27.91166, -27.71076, 
    -27.50902, -27.30642, -27.10297, -26.89865, -26.69348, -26.48744, 
    -26.28053, -26.07275, -25.8641, -25.65456, -25.44415, -25.23284, 
    -25.02065, -24.80757, -24.59359, -24.37872, -24.16294, -23.94626, 
    -23.72867, -23.51017, -23.29076, -23.07044, -22.84919, -22.62703, 
    -22.40394, -22.17993, -21.95499, -21.72911, -21.50231, -21.27457, 
    -21.04589, -20.81627, -20.58571, -20.3542, -20.12175, -19.88835, -19.654, 
    -19.4187, -19.18245, -18.94524, -18.70708, -18.46796, -18.22788, 
    -17.98684, -17.74484, -17.50187, -17.25795, -17.01306, -16.7672, 
    -16.52038, -16.2726, -16.02384, -15.77413, -15.52344, -15.27179, 
    -15.01917, -14.76558, -14.51103, -14.25552, -13.99903, -13.74158, 
    -13.48317, -13.2238, -12.96346, -12.70216, -12.4399, -12.17669, 
    -11.91251, -11.64738, -11.3813, -11.11427, -10.84629, -10.57736, 
    -10.30748, -10.03667, -9.764915, -9.492224, -9.218599, -8.944045, 
    -8.668565, -8.39216, -8.114838, -7.836598, -7.557447, -7.27739, 
    -6.996428, -6.714568, -6.431815, -6.148172, -5.863645, -5.578239, 
    -5.29196, -5.004813, -4.716804, -4.427938, -4.138223, -3.847663, 
    -3.556266, -3.264038, -2.970986, -2.677117, -2.382438, -2.086957, 
    -1.790681, -1.493617, -1.195775, -0.8971605, -0.5977834, -0.2976518, 
    0.003225795, 0.3048405, 0.6071833, 0.9102451, 1.214016, 1.518488, 
    1.82365, 2.129492, 2.436005, 2.743178, 3.051001, 3.359463, 3.668554, 
    3.978262, 4.288577, 4.599487, 4.910981, 5.223047, 5.535674, 5.84885, 
    6.162562, 6.476799, 6.791549, 7.106798, 7.422534, 7.738745, 8.055417, 
    8.372538, 8.690094, 9.008072, 9.326458, 9.64524, 9.964403, 10.28393, 
    10.60382, 10.92404, 11.24459, 11.56546, 11.88662, 12.20806, 12.52977, 
    12.85174, 13.17394, 13.49637, 13.81901, 14.14184, 14.46486, 14.78804, 
    15.11137, 15.43484, 15.75842, 16.08212, 16.4059, 16.72975, 17.05367, 
    17.37763, 17.70162, 18.02563, 18.34963, 18.67362, 18.99757, 19.32148, 
    19.64532, 19.96909, 20.29277, 20.61634, 20.93978, 21.26309, 21.58625, 
    21.90924, 22.23204, 22.55465, 22.87704, 23.19921, 23.52114, 23.84281, 
    24.1642, 24.48532, 24.80613, 25.12663, 25.4468, 25.76663, 26.08611, 
    26.40521, 26.72393, 27.04226, 27.36017, 27.67765, 27.99471, 28.31131, 
    28.62744, 28.9431, 29.25827, 29.57294, 29.8871, 30.20073, 30.51381, 
    30.82635, 31.13833, 31.44973, 31.76055, 32.07077, 32.38038, 32.68937, 
    32.99773, 33.30545, 33.61253, 33.91893, 34.22467, 34.52972, 34.83408, 
    35.13774, 35.44069, 35.74292, 36.04442, 36.34518, 36.64519, 36.94445, 
    37.24294, 37.54066, 37.8376, 38.13375, 38.4291, 38.72366, 39.0174, 
    39.31032, 39.60242, 39.89368, 40.18411, 40.47369, 40.76242, 41.05029, 
    41.3373, 41.62344, 41.90871, 42.1931, 42.4766, 42.75921, 43.04093, 
    43.32175, 43.60167, 43.88067, 44.15877, 44.43594, 44.7122, 44.98754, 
    45.26194, 45.53542, 45.80796, 46.07957, 46.35023, 46.61996, 46.88874, 
    47.15657, 47.42345, 47.68938, 47.95436, 48.21839, 48.48145, 48.74356, 
    49.0047, 49.26489, 49.52411, 49.78237, 50.03967, 50.296, 50.55136, 
    50.80576, 51.05919, 51.31166, 51.56316, 51.81369, 52.06326, 52.31186, 
    52.55949, 52.80616, 53.05186, 53.2966, 53.54037, 53.78318, 54.02503, 
    54.26592, 54.50585, 54.74482, 54.98283, 55.21989, 55.45599, 55.69114, 
    55.92533, 56.15858, 56.39088, 56.62224, 56.85265, 57.08212, 57.31065, 
    57.53825, 57.7649, 57.99063, 58.21542, 58.43929, 58.66223, 58.88425, 
    59.10535, 59.32553, 59.5448, 59.76315, 59.98059, 60.19713, 60.41277, 
    60.6275, 60.84134, 61.05428, 61.26633, 61.47749, 61.68777, 61.89716, 
    62.10568, 62.31332, 62.52009, 62.72599, 62.93103, 63.13521, 63.33852, 
    63.54099, 63.7426, 63.94336, 64.14328, 64.34236, 64.5406,
  -43.97513, -43.83844, -43.70126, -43.56357, -43.42537, -43.28667, 
    -43.14745, -43.00771, -42.86745, -42.72667, -42.58536, -42.44352, 
    -42.30115, -42.15824, -42.01479, -41.8708, -41.72626, -41.58117, 
    -41.43553, -41.28933, -41.14257, -40.99525, -40.84736, -40.6989, 
    -40.54987, -40.40026, -40.25007, -40.09929, -39.94793, -39.79597, 
    -39.64342, -39.49027, -39.33652, -39.18216, -39.02719, -38.87161, 
    -38.71541, -38.55859, -38.40115, -38.24308, -38.08438, -37.92504, 
    -37.76506, -37.60445, -37.44318, -37.28126, -37.11869, -36.95546, 
    -36.79158, -36.62702, -36.4618, -36.2959, -36.12932, -35.96207, 
    -35.79413, -35.6255, -35.45618, -35.28616, -35.11544, -34.94402, 
    -34.77189, -34.59905, -34.4255, -34.25122, -34.07622, -33.90049, 
    -33.72403, -33.54684, -33.3689, -33.19023, -33.01081, -32.83063, 
    -32.6497, -32.46801, -32.28556, -32.10234, -31.91836, -31.73359, 
    -31.54805, -31.36173, -31.17462, -30.98672, -30.79803, -30.60853, 
    -30.41824, -30.22714, -30.03523, -29.84251, -29.64897, -29.45461, 
    -29.25943, -29.06342, -28.86657, -28.66889, -28.47037, -28.27101, 
    -28.07079, -27.86973, -27.66782, -27.46504, -27.26141, -27.0569, 
    -26.85154, -26.64529, -26.43818, -26.23018, -26.0213, -25.81153, 
    -25.60088, -25.38934, -25.17689, -24.96355, -24.74931, -24.53416, 
    -24.3181, -24.10113, -23.88325, -23.66445, -23.44473, -23.22408, 
    -23.00251, -22.78001, -22.55658, -22.33221, -22.10691, -21.88067, 
    -21.65349, -21.42536, -21.19629, -20.96626, -20.73529, -20.50336, 
    -20.27048, -20.03664, -19.80184, -19.56609, -19.32936, -19.09168, 
    -18.85303, -18.61341, -18.37283, -18.13127, -17.88874, -17.64524, 
    -17.40077, -17.15532, -16.9089, -16.66151, -16.41313, -16.16378, 
    -15.91346, -15.66215, -15.40987, -15.15661, -14.90238, -14.64716, 
    -14.39097, -14.1338, -13.87566, -13.61654, -13.35645, -13.09538, 
    -12.83335, -12.57034, -12.30636, -12.04141, -11.77549, -11.50862, 
    -11.24077, -10.97197, -10.70221, -10.43149, -10.15982, -9.887197, 
    -9.613626, -9.339111, -9.063654, -8.787257, -8.509926, -8.231664, 
    -7.952473, -7.672359, -7.391326, -7.109377, -6.826518, -6.542753, 
    -6.258087, -5.972525, -5.686072, -5.398734, -5.110515, -4.821423, 
    -4.531462, -4.24064, -3.948961, -3.656434, -3.363064, -3.068858, 
    -2.773823, -2.477968, -2.181298, -1.883821, -1.585546, -1.28648, 
    -0.9866313, -0.6860086, -0.3846203, -0.0824749, 0.2204185, 0.524051, 
    0.8284132, 1.133496, 1.439289, 1.745783, 2.052968, 2.360833, 2.669369, 
    2.978565, 3.288409, 3.598892, 3.910002, 4.221728, 4.534059, 4.846983, 
    5.160488, 5.474563, 5.789195, 6.104372, 6.420082, 6.736312, 7.05305, 
    7.370283, 7.687998, 8.006183, 8.324821, 8.643904, 8.963415, 9.283341, 
    9.603669, 9.924384, 10.24547, 10.56692, 10.88872, 11.21084, 11.53328, 
    11.85603, 12.17906, 12.50237, 12.82593, 13.14973, 13.47377, 13.79802, 
    14.12247, 14.4471, 14.77189, 15.09685, 15.42193, 15.74715, 16.07246, 
    16.39787, 16.72336, 17.04891, 17.3745, 17.70012, 18.02575, 18.35139, 
    18.67701, 19.00259, 19.32813, 19.65361, 19.979, 20.3043, 20.6295, 
    20.95457, 21.27949, 21.60427, 21.92887, 22.25329, 22.5775, 22.9015, 
    23.22527, 23.54879, 23.87206, 24.19504, 24.51774, 24.84013, 25.16221, 
    25.48395, 25.80534, 26.12637, 26.44703, 26.76729, 27.08715, 27.4066, 
    27.72561, 28.04418, 28.36229, 28.67993, 28.99709, 29.31374, 29.62989, 
    29.94552, 30.26061, 30.57516, 30.88914, 31.20255, 31.51539, 31.82762, 
    32.13925, 32.45026, 32.76065, 33.07039, 33.37948, 33.68791, 33.99567, 
    34.30275, 34.60913, 34.91481, 35.21978, 35.52403, 35.82755, 36.13032, 
    36.43235, 36.73361, 37.03411, 37.33384, 37.63278, 37.93093, 38.22828, 
    38.52482, 38.82055, 39.11545, 39.40953, 39.70276, 39.99516, 40.2867, 
    40.57738, 40.86721, 41.15617, 41.44424, 41.73144, 42.01775, 42.30318, 
    42.5877, 42.87132, 43.15404, 43.43584, 43.71673, 43.9967, 44.27574, 
    44.55386, 44.83104, 45.10729, 45.3826, 45.65696, 45.93039, 46.20286, 
    46.47438, 46.74495, 47.01455, 47.28321, 47.5509, 47.81762, 48.08338, 
    48.34818, 48.612, 48.87486, 49.13675, 49.39766, 49.6576, 49.91656, 
    50.17455, 50.43156, 50.6876, 50.94266, 51.19674, 51.44984, 51.70197, 
    51.95312, 52.20329, 52.45249, 52.70071, 52.94795, 53.19421, 53.43951, 
    53.68383, 53.92717, 54.16954, 54.41095, 54.65138, 54.89084, 55.12934, 
    55.36687, 55.60344, 55.83905, 56.0737, 56.30738, 56.54011, 56.77189, 
    57.00271, 57.23258, 57.46151, 57.68948, 57.91652, 58.14261, 58.36777, 
    58.59198, 58.81527, 59.03762, 59.25904, 59.47954, 59.69912, 59.91777, 
    60.13551, 60.35234, 60.56825, 60.78326, 60.99736, 61.21056, 61.42286, 
    61.63426, 61.84478, 62.0544, 62.26314, 62.471, 62.67797, 62.88408, 
    63.08931, 63.29367, 63.49717, 63.69981, 63.90159, 64.10252, 64.3026, 
    64.50183, 64.70022,
  -44.13209, -43.99555, -43.85851, -43.72097, -43.58291, -43.44434, 
    -43.30526, -43.16566, -43.02554, -42.8849, -42.74372, -42.60202, 
    -42.45978, -42.317, -42.17368, -42.02982, -41.8854, -41.74044, -41.59492, 
    -41.44884, -41.3022, -41.15499, -41.00723, -40.85888, -40.70996, 
    -40.56046, -40.41037, -40.2597, -40.10844, -39.95658, -39.80413, 
    -39.65108, -39.49743, -39.34316, -39.18828, -39.03279, -38.87668, 
    -38.71994, -38.56258, -38.40459, -38.24597, -38.0867, -37.9268, 
    -37.76625, -37.60505, -37.4432, -37.28069, -37.11752, -36.95368, 
    -36.78918, -36.624, -36.45815, -36.29162, -36.1244, -35.9565, -35.78791, 
    -35.61862, -35.44863, -35.27793, -35.10653, -34.93442, -34.76159, 
    -34.58804, -34.41377, -34.23877, -34.06304, -33.88658, -33.70937, 
    -33.53143, -33.35273, -33.17329, -32.99309, -32.81213, -32.6304, 
    -32.44791, -32.26465, -32.08062, -31.8958, -31.7102, -31.52381, 
    -31.33664, -31.14866, -30.95989, -30.77032, -30.57994, -30.38875, 
    -30.19674, -30.00392, -29.81027, -29.6158, -29.42049, -29.22435, 
    -29.02738, -28.82956, -28.6309, -28.43139, -28.23102, -28.0298, 
    -27.82771, -27.62477, -27.42095, -27.21626, -27.0107, -26.80426, 
    -26.59694, -26.38873, -26.17963, -25.96964, -25.75875, -25.54697, 
    -25.33428, -25.12068, -24.90617, -24.69076, -24.47442, -24.25717, 
    -24.03899, -23.81989, -23.59986, -23.3789, -23.157, -22.93417, -22.7104, 
    -22.48568, -22.26002, -22.03341, -21.80586, -21.57734, -21.34788, 
    -21.11745, -20.88607, -20.65372, -20.42041, -20.18614, -19.95089, 
    -19.71468, -19.47749, -19.23933, -19.00019, -18.76008, -18.51899, 
    -18.27692, -18.03387, -17.78983, -17.54482, -17.29881, -17.05182, 
    -16.80385, -16.55489, -16.30494, -16.05401, -15.80209, -15.54917, 
    -15.29527, -15.04039, -14.78451, -14.52765, -14.26979, -14.01095, 
    -13.75113, -13.49032, -13.22852, -12.96574, -12.70198, -12.43723, 
    -12.17151, -11.9048, -11.63712, -11.36847, -11.09884, -10.82825, 
    -10.55668, -10.28415, -10.01066, -9.736201, -9.46079, -9.184424, 
    -8.907108, -8.628844, -8.349638, -8.06949, -7.788408, -7.506393, 
    -7.223452, -6.939588, -6.654805, -6.369109, -6.082505, -5.794998, 
    -5.506593, -5.217296, -4.927113, -4.63605, -4.344112, -4.051307, 
    -3.757641, -3.46312, -3.167751, -2.871542, -2.574499, -2.276631, 
    -1.977944, -1.678447, -1.378148, -1.077055, -0.7751755, -0.4725195, 
    -0.1690952, 0.1350883, 0.440022, 0.7456964, 1.052102, 1.359229, 1.667067, 
    1.975607, 2.284838, 2.59475, 2.905332, 3.216572, 3.528461, 3.840987, 
    4.154139, 4.467904, 4.782272, 5.09723, 5.412767, 5.72887, 6.045527, 
    6.362726, 6.680453, 6.998696, 7.317442, 7.636677, 7.956389, 8.276565, 
    8.597189, 8.91825, 9.239733, 9.561623, 9.883907, 10.20657, 10.5296, 
    10.85298, 11.1767, 11.50074, 11.82509, 12.14973, 12.47464, 12.79982, 
    13.12525, 13.45091, 13.77678, 14.10286, 14.42913, 14.75556, 15.08215, 
    15.40888, 15.73574, 16.0627, 16.38976, 16.71689, 17.04409, 17.37133, 
    17.6986, 18.02589, 18.35317, 18.68044, 19.00768, 19.33486, 19.66198, 
    19.98903, 20.31598, 20.64281, 20.96952, 21.29609, 21.6225, 21.94873, 
    22.27478, 22.60062, 22.92624, 23.25163, 23.57677, 23.90165, 24.22624, 
    24.55054, 24.87453, 25.19819, 25.52152, 25.84449, 26.1671, 26.48932, 
    26.81115, 27.13256, 27.45356, 27.77411, 28.09422, 28.41385, 28.73301, 
    29.05168, 29.36984, 29.68748, 30.0046, 30.32117, 30.63718, 30.95263, 
    31.26749, 31.58177, 31.89544, 32.20849, 32.52092, 32.8327, 33.14384, 
    33.45432, 33.76412, 34.07325, 34.38168, 34.6894, 34.99641, 35.3027, 
    35.60826, 35.91308, 36.21714, 36.52045, 36.82298, 37.12474, 37.4257, 
    37.72588, 38.02525, 38.3238, 38.62154, 38.91845, 39.21453, 39.50977, 
    39.80415, 40.09768, 40.39035, 40.68215, 40.97307, 41.26312, 41.55227, 
    41.84054, 42.1279, 42.41436, 42.69991, 42.98455, 43.26827, 43.55106, 
    43.83293, 44.11387, 44.39387, 44.67292, 44.95104, 45.2282, 45.50442, 
    45.77968, 46.05398, 46.32732, 46.5997, 46.87111, 47.14156, 47.41103, 
    47.67953, 47.94706, 48.2136, 48.47918, 48.74376, 49.00737, 49.27, 
    49.53164, 49.79229, 50.05196, 50.31065, 50.56834, 50.82505, 51.08077, 
    51.3355, 51.58924, 51.842, 52.09377, 52.34455, 52.59434, 52.84314, 
    53.09096, 53.33779, 53.58364, 53.8285, 54.07238, 54.31528, 54.55719, 
    54.79813, 55.03809, 55.27707, 55.51508, 55.75211, 55.98817, 56.22326, 
    56.45739, 56.69054, 56.92274, 57.15397, 57.38424, 57.61356, 57.84192, 
    58.06932, 58.29578, 58.52129, 58.74586, 58.96948, 59.19217, 59.41391, 
    59.63472, 59.85461, 60.07356, 60.2916, 60.5087, 60.72489, 60.94017, 
    61.15453, 61.36798, 61.58053, 61.79217, 62.00292, 62.21277, 62.42173, 
    62.6298, 62.83698, 63.04328, 63.2487, 63.45325, 63.65693, 63.85974, 
    64.06168, 64.26277, 64.46301, 64.66238, 64.86091,
  -44.28974, -44.15335, -44.01646, -43.87906, -43.74115, -43.60273, 
    -43.46379, -43.32434, -43.18436, -43.04385, -42.90281, -42.76125, 
    -42.61914, -42.4765, -42.33331, -42.18958, -42.04529, -41.90046, 
    -41.75506, -41.60911, -41.46259, -41.31551, -41.16786, -41.01963, 
    -40.87082, -40.72144, -40.57146, -40.4209, -40.26975, -40.118, -39.96566, 
    -39.81271, -39.65915, -39.50498, -39.3502, -39.1948, -39.03878, 
    -38.88214, -38.72486, -38.56695, -38.40841, -38.24923, -38.0894, 
    -37.92892, -37.76779, -37.60601, -37.44356, -37.28045, -37.11668, 
    -36.95223, -36.78711, -36.62131, -36.45483, -36.28765, -36.11979, 
    -35.95123, -35.78198, -35.61202, -35.44135, -35.26998, -35.09789, 
    -34.92507, -34.75154, -34.57728, -34.40229, -34.22656, -34.05009, 
    -33.87288, -33.69493, -33.51622, -33.33675, -33.15653, -32.97555, 
    -32.79379, -32.61127, -32.42797, -32.24389, -32.05902, -31.87337, 
    -31.68693, -31.49969, -31.31165, -31.1228, -30.93315, -30.74269, 
    -30.55141, -30.35931, -30.16638, -29.97263, -29.77805, -29.58263, 
    -29.38637, -29.18927, -28.99132, -28.79252, -28.59286, -28.39235, 
    -28.19097, -27.98872, -27.7856, -27.58162, -27.37675, -27.171, -26.96436, 
    -26.75684, -26.54842, -26.3391, -26.12889, -25.91777, -25.70575, 
    -25.49282, -25.27897, -25.0642, -24.84852, -24.63191, -24.41437, 
    -24.19591, -23.97651, -23.75617, -23.5349, -23.31268, -23.08952, 
    -22.86541, -22.64035, -22.41433, -22.18736, -21.95943, -21.73054, 
    -21.50068, -21.26986, -21.03807, -20.8053, -20.57157, -20.33685, 
    -20.10116, -19.86449, -19.62684, -19.38821, -19.14859, -18.90798, 
    -18.66639, -18.4238, -18.18023, -17.93566, -17.69009, -17.44354, 
    -17.19598, -16.94743, -16.69789, -16.44734, -16.1958, -15.94326, 
    -15.68971, -15.43517, -15.17963, -14.92309, -14.66555, -14.40701, 
    -14.14748, -13.88694, -13.62541, -13.36288, -13.09936, -12.83484, 
    -12.56933, -12.30282, -12.03533, -11.76685, -11.49738, -11.22692, 
    -10.95549, -10.68307, -10.40968, -10.13531, -9.859964, -9.583652, 
    -9.306375, -9.028133, -8.748933, -8.468777, -8.187668, -7.905611, 
    -7.62261, -7.338669, -7.053793, -6.767987, -6.481255, -6.193602, 
    -5.905033, -5.615555, -5.325172, -5.033891, -4.741717, -4.448657, 
    -4.154716, -3.859902, -3.564221, -3.267681, -2.970288, -2.672049, 
    -2.372972, -2.073066, -1.772337, -1.470794, -1.168445, -0.8652994, 
    -0.5613647, -0.2566502, 0.04883488, 0.3550814, 0.6620799, 0.9698206, 
    1.278294, 1.587489, 1.897397, 2.208007, 2.519307, 2.831289, 3.143939, 
    3.457248, 3.771204, 4.085795, 4.40101, 4.716836, 5.033263, 5.350277, 
    5.667867, 5.98602, 6.304722, 6.623961, 6.943725, 7.264, 7.584772, 
    7.906029, 8.227757, 8.54994, 8.872567, 9.195623, 9.519094, 9.842965, 
    10.16722, 10.49185, 10.81684, 11.14217, 11.46782, 11.79379, 12.12005, 
    12.4466, 12.77341, 13.10048, 13.42778, 13.7553, 14.08303, 14.41095, 
    14.73904, 15.06729, 15.39568, 15.72419, 16.05282, 16.38154, 16.71035, 
    17.03921, 17.36812, 17.69706, 18.02602, 18.35497, 18.68391, 19.01282, 
    19.34167, 19.67046, 19.99917, 20.32778, 20.65628, 20.98465, 21.31287, 
    21.64094, 21.96882, 22.29652, 22.62401, 22.95127, 23.2783, 23.60507, 
    23.93158, 24.2578, 24.58371, 24.90932, 25.23459, 25.55952, 25.88409, 
    26.20829, 26.5321, 26.85551, 27.1785, 27.50105, 27.82317, 28.14482, 
    28.466, 28.7867, 29.10689, 29.42657, 29.74573, 30.06434, 30.38241, 
    30.69991, 31.01683, 31.33316, 31.64889, 31.96401, 32.2785, 32.59235, 
    32.90556, 33.21811, 33.52998, 33.84117, 34.15167, 34.46147, 34.77055, 
    35.07891, 35.38653, 35.69341, 35.99954, 36.3049, 36.60949, 36.9133, 
    37.21632, 37.51855, 37.81996, 38.12056, 38.42034, 38.71928, 39.01739, 
    39.31464, 39.61105, 39.90659, 40.20127, 40.49507, 40.78799, 41.08002, 
    41.37117, 41.66141, 41.95074, 42.23917, 42.52667, 42.81326, 43.09892, 
    43.38365, 43.66744, 43.95029, 44.2322, 44.51316, 44.79316, 45.07221, 
    45.3503, 45.62743, 45.90358, 46.17877, 46.45299, 46.72623, 46.99849, 
    47.26977, 47.54007, 47.80938, 48.07771, 48.34505, 48.61139, 48.87675, 
    49.14111, 49.40448, 49.66685, 49.92822, 50.1886, 50.44798, 50.70636, 
    50.96374, 51.22012, 51.4755, 51.72989, 51.98327, 52.23565, 52.48704, 
    52.73743, 52.98682, 53.23521, 53.4826, 53.729, 53.97441, 54.21882, 
    54.46224, 54.70467, 54.94611, 55.18656, 55.42602, 55.6645, 55.902, 
    56.13851, 56.37405, 56.6086, 56.84219, 57.0748, 57.30643, 57.53711, 
    57.76681, 57.99555, 58.22333, 58.45015, 58.67601, 58.90092, 59.12489, 
    59.3479, 59.56997, 59.79109, 60.01128, 60.23053, 60.44884, 60.66624, 
    60.8827, 61.09824, 61.31285, 61.52656, 61.73935, 61.95123, 62.1622, 
    62.37227, 62.58145, 62.78972, 62.9971, 63.2036, 63.40921, 63.61394, 
    63.81779, 64.02077, 64.22288, 64.42412, 64.6245, 64.82402, 65.02269,
  -44.44808, -44.31184, -44.1751, -44.03786, -43.9001, -43.76183, -43.62304, 
    -43.48373, -43.34389, -43.20353, -43.06263, -42.92121, -42.77924, 
    -42.63673, -42.49369, -42.35009, -42.20594, -42.06123, -41.91597, 
    -41.77015, -41.62376, -41.4768, -41.32927, -41.18116, -41.03248, 
    -40.88321, -40.73335, -40.58291, -40.43187, -40.28023, -40.12799, 
    -39.97515, -39.82169, -39.66763, -39.51295, -39.35765, -39.20172, 
    -39.04517, -38.88799, -38.73016, -38.5717, -38.41261, -38.25286, 
    -38.09246, -37.9314, -37.76969, -37.60732, -37.44427, -37.28056, 
    -37.11618, -36.95111, -36.78537, -36.61894, -36.45182, -36.284, 
    -36.11549, -35.94627, -35.77634, -35.60571, -35.43436, -35.26229, 
    -35.08951, -34.91599, -34.74174, -34.56676, -34.39104, -34.21458, 
    -34.03737, -33.85941, -33.68069, -33.50122, -33.32098, -33.13997, 
    -32.95819, -32.77563, -32.5923, -32.40818, -32.22327, -32.03757, 
    -31.85107, -31.66377, -31.47567, -31.28676, -31.09703, -30.90649, 
    -30.71513, -30.52294, -30.32992, -30.13607, -29.94138, -29.74586, 
    -29.54948, -29.35225, -29.15418, -28.95524, -28.75545, -28.55478, 
    -28.35325, -28.15085, -27.94757, -27.74341, -27.53836, -27.33242, 
    -27.1256, -26.91788, -26.70925, -26.49973, -26.2893, -26.07795, -25.8657, 
    -25.65252, -25.43843, -25.22341, -25.00746, -24.79058, -24.57277, 
    -24.35402, -24.13432, -23.91368, -23.6921, -23.46956, -23.24608, 
    -23.02163, -22.79623, -22.56986, -22.34253, -22.11423, -21.88495, 
    -21.65471, -21.42349, -21.19129, -20.95811, -20.72395, -20.48881, 
    -20.25267, -20.01555, -19.77744, -19.53833, -19.29823, -19.05713, 
    -18.81503, -18.57193, -18.32783, -18.08273, -17.83662, -17.58951, 
    -17.34139, -17.09227, -16.84213, -16.59099, -16.33884, -16.08568, 
    -15.83151, -15.57632, -15.32013, -15.06293, -14.80471, -14.54548, 
    -14.28525, -14.024, -13.76175, -13.49849, -13.23422, -12.96894, 
    -12.70266, -12.43537, -12.16709, -11.8978, -11.62751, -11.35623, 
    -11.08395, -10.81068, -10.53642, -10.26117, -9.984932, -9.707716, 
    -9.429522, -9.150352, -8.870209, -8.589098, -8.307022, -8.023985, 
    -7.739992, -7.455046, -7.169153, -6.882316, -6.594541, -6.305832, 
    -6.016196, -5.725636, -5.43416, -5.141773, -4.848481, -4.554289, 
    -4.259205, -3.963235, -3.666386, -3.368665, -3.070078, -2.770634, 
    -2.47034, -2.169203, -1.867232, -1.564435, -1.26082, -0.956396, 
    -0.6511714, -0.3451555, -0.03835716, 0.2692141, 0.5775487, 0.886637, 
    1.196469, 1.507034, 1.818323, 2.130324, 2.443027, 2.756422, 3.070496, 
    3.385239, 3.700638, 4.016684, 4.333363, 4.650663, 4.968573, 5.28708, 
    5.606172, 5.925835, 6.246058, 6.566825, 6.888126, 7.209947, 7.532272, 
    7.855091, 8.178387, 8.502148, 8.826359, 9.151006, 9.476074, 9.80155, 
    10.12742, 10.45366, 10.78027, 11.10723, 11.43452, 11.76212, 12.09003, 
    12.41823, 12.7467, 13.07542, 13.40438, 13.73357, 14.06297, 14.39255, 
    14.72232, 15.05225, 15.38232, 15.71252, 16.04283, 16.37324, 16.70372, 
    17.03428, 17.36488, 17.69551, 18.02615, 18.3568, 18.68742, 19.01801, 
    19.34856, 19.67904, 20.00943, 20.33972, 20.6699, 20.99995, 21.32985, 
    21.65959, 21.98915, 22.31852, 22.64767, 22.97659, 23.30528, 23.63371, 
    23.96185, 24.28972, 24.61728, 24.94451, 25.27142, 25.59797, 25.92415, 
    26.24996, 26.57537, 26.90038, 27.22496, 27.5491, 27.87278, 28.19601, 
    28.51875, 28.84099, 29.16273, 29.48395, 29.80463, 30.12477, 30.44434, 
    30.76334, 31.08175, 31.39957, 31.71677, 32.03335, 32.3493, 32.66459, 
    32.97923, 33.2932, 33.60648, 33.91908, 34.23096, 34.54214, 34.85259, 
    35.1623, 35.47128, 35.77949, 36.08694, 36.39362, 36.6995, 37.0046, 
    37.3089, 37.61239, 37.91505, 38.21689, 38.5179, 38.81806, 39.11737, 
    39.41582, 39.7134, 40.01011, 40.30594, 40.60088, 40.89494, 41.18808, 
    41.48033, 41.77166, 42.06207, 42.35156, 42.64013, 42.92775, 43.21444, 
    43.50018, 43.78498, 44.06882, 44.3517, 44.63363, 44.91459, 45.19458, 
    45.47359, 45.75163, 46.02869, 46.30477, 46.57986, 46.85397, 47.12708, 
    47.3992, 47.67033, 47.94046, 48.20959, 48.47772, 48.74485, 49.01097, 
    49.27608, 49.5402, 49.8033, 50.0654, 50.32648, 50.58656, 50.84562, 
    51.10368, 51.36072, 51.61676, 51.87178, 52.12579, 52.37879, 52.63079, 
    52.88177, 53.13174, 53.38071, 53.62867, 53.87562, 54.12157, 54.36651, 
    54.61045, 54.85339, 55.09533, 55.33627, 55.57622, 55.81517, 56.05312, 
    56.29009, 56.52607, 56.76106, 56.99506, 57.22809, 57.46013, 57.6912, 
    57.92129, 58.1504, 58.37855, 58.60573, 58.83194, 59.0572, 59.28149, 
    59.50483, 59.72721, 59.94865, 60.16914, 60.38868, 60.60728, 60.82495, 
    61.04168, 61.25748, 61.47235, 61.68631, 61.89933, 62.11145, 62.32264, 
    62.53293, 62.74231, 62.95079, 63.15837, 63.36506, 63.57085, 63.77576, 
    63.97978, 64.18292, 64.38519, 64.58659, 64.78711, 64.98677, 65.18557,
  -44.60711, -44.47104, -44.33445, -44.19736, -44.05975, -43.92163, -43.783, 
    -43.64384, -43.50415, -43.36393, -43.22319, -43.08191, -42.94008, 
    -42.79772, -42.65481, -42.51135, -42.36734, -42.22277, -42.07764, 
    -41.93195, -41.78569, -41.63887, -41.49147, -41.34348, -41.19492, 
    -41.04578, -40.89604, -40.74572, -40.59479, -40.44327, -40.29114, 
    -40.13841, -39.98507, -39.83111, -39.67653, -39.52133, -39.36551, 
    -39.20905, -39.05196, -38.89423, -38.73586, -38.57685, -38.41719, 
    -38.25687, -38.09589, -37.93426, -37.77196, -37.60899, -37.44535, 
    -37.28103, -37.11603, -36.95034, -36.78397, -36.6169, -36.44913, 
    -36.28067, -36.11149, -35.94161, -35.77102, -35.5997, -35.42766, 
    -35.2549, -35.08141, -34.90718, -34.73222, -34.55651, -34.38005, 
    -34.20285, -34.02488, -33.84616, -33.66668, -33.48643, -33.3054, 
    -33.1236, -32.94102, -32.75765, -32.5735, -32.38855, -32.20281, 
    -32.01626, -31.82891, -31.64075, -31.45177, -31.26198, -31.07136, 
    -30.87992, -30.68765, -30.49454, -30.3006, -30.10581, -29.91017, 
    -29.71369, -29.51634, -29.31814, -29.11908, -28.91915, -28.71834, 
    -28.51666, -28.3141, -28.11066, -27.90633, -27.70111, -27.495, -27.28799, 
    -27.08007, -26.87125, -26.66152, -26.45087, -26.2393, -26.02682, 
    -25.81341, -25.59907, -25.3838, -25.16759, -24.95045, -24.73236, 
    -24.51332, -24.29334, -24.0724, -23.85051, -23.62766, -23.40385, 
    -23.17907, -22.95333, -22.72661, -22.49892, -22.27025, -22.0406, 
    -21.80997, -21.57836, -21.34576, -21.11217, -20.87759, -20.64201, 
    -20.40543, -20.16786, -19.92928, -19.6897, -19.44912, -19.20753, 
    -18.96493, -18.72132, -18.4767, -18.23107, -17.98442, -17.73675, 
    -17.48807, -17.23837, -16.98765, -16.73591, -16.48315, -16.22937, 
    -15.97457, -15.71874, -15.46189, -15.20403, -14.94513, -14.68522, 
    -14.42428, -14.16233, -13.89935, -13.63535, -13.37033, -13.1043, 
    -12.83724, -12.56918, -12.30009, -12.03, -11.75889, -11.48677, -11.21365, 
    -10.93952, -10.66438, -10.38825, -10.11112, -9.832998, -9.553883, 
    -9.273778, -8.992689, -8.710618, -8.42757, -8.143548, -7.858557, -7.5726, 
    -7.285683, -6.997809, -6.708985, -6.419214, -6.128502, -5.836855, 
    -5.544278, -5.250777, -4.956358, -4.661027, -4.364791, -4.067657, 
    -3.76963, -3.470718, -3.170929, -2.87027, -2.568748, -2.266371, 
    -1.963148, -1.659086, -1.354195, -1.048481, -0.7419558, -0.4346267, 
    -0.1265034, 0.1824045, 0.4920876, 0.8025358, 1.113739, 1.425687, 1.73837, 
    2.051776, 2.365896, 2.680717, 2.996229, 3.312419, 3.629278, 3.946792, 
    4.26495, 4.58374, 4.903148, 5.223164, 5.543773, 5.864963, 6.186721, 
    6.509035, 6.831889, 7.155271, 7.479167, 7.803564, 8.128447, 8.453801, 
    8.779613, 9.105869, 9.432553, 9.759651, 10.08715, 10.41503, 10.74328, 
    11.07188, 11.40082, 11.73009, 12.05966, 12.38953, 12.71966, 13.05007, 
    13.38071, 13.71158, 14.04266, 14.37395, 14.70541, 15.03703, 15.3688, 
    15.7007, 16.03271, 16.36483, 16.69702, 17.02928, 17.36159, 17.69393, 
    18.02629, 18.35864, 18.69098, 19.02328, 19.35553, 19.68771, 20.01981, 
    20.35181, 20.68369, 21.01544, 21.34704, 21.67847, 22.00972, 22.34077, 
    22.67161, 23.00222, 23.33257, 23.66267, 23.99249, 24.32202, 24.65123, 
    24.98012, 25.30867, 25.63686, 25.96468, 26.29212, 26.61915, 26.94577, 
    27.27195, 27.59769, 27.92298, 28.24778, 28.5721, 28.89592, 29.21922, 
    29.54199, 29.86421, 30.18588, 30.50698, 30.8275, 31.14742, 31.46673, 
    31.78542, 32.10348, 32.42089, 32.73764, 33.05373, 33.36913, 33.68384, 
    33.99785, 34.31114, 34.62371, 34.93554, 35.24662, 35.55695, 35.86651, 
    36.1753, 36.4833, 36.7905, 37.09689, 37.40248, 37.70724, 38.01117, 
    38.31426, 38.6165, 38.91788, 39.21841, 39.51806, 39.81683, 40.11472, 
    40.41171, 40.70781, 41.00299, 41.29726, 41.59062, 41.88305, 42.17455, 
    42.46511, 42.75473, 43.04341, 43.33113, 43.6179, 43.9037, 44.18854, 
    44.47241, 44.7553, 45.03722, 45.31815, 45.5981, 45.87706, 46.15503, 
    46.432, 46.70797, 46.98295, 47.25692, 47.52988, 47.80184, 48.07279, 
    48.34272, 48.61165, 48.87955, 49.14645, 49.41232, 49.67718, 49.94102, 
    50.20383, 50.46563, 50.7264, 50.98615, 51.24488, 51.50259, 51.75928, 
    52.01494, 52.26958, 52.5232, 52.7758, 53.02738, 53.27794, 53.52747, 
    53.776, 54.0235, 54.26999, 54.51546, 54.75993, 55.00337, 55.24582, 
    55.48724, 55.72767, 55.96709, 56.20551, 56.44292, 56.67934, 56.91476, 
    57.14919, 57.38262, 57.61507, 57.84652, 58.077, 58.30649, 58.535, 
    58.76254, 58.9891, 59.21469, 59.43932, 59.66298, 59.88567, 60.10741, 
    60.3282, 60.54803, 60.76692, 60.98486, 61.20185, 61.41791, 61.63304, 
    61.84723, 62.06049, 62.27283, 62.48425, 62.69475, 62.90434, 63.11302, 
    63.32079, 63.52766, 63.73364, 63.93872, 64.14291, 64.34621, 64.54862, 
    64.75016, 64.95083, 65.15063, 65.34955,
  -44.76685, -44.63093, -44.4945, -44.35757, -44.22012, -44.08216, -43.94368, 
    -43.80467, -43.66514, -43.52508, -43.38448, -43.24335, -43.10167, 
    -42.95945, -42.81669, -42.67337, -42.5295, -42.38508, -42.24009, 
    -42.09454, -41.94841, -41.80172, -41.65445, -41.5066, -41.35817, 
    -41.20914, -41.05954, -40.90933, -40.75853, -40.60712, -40.45512, 
    -40.3025, -40.14927, -39.99542, -39.84095, -39.68586, -39.53014, 
    -39.37378, -39.21679, -39.05916, -38.90089, -38.74197, -38.58239, 
    -38.42216, -38.26127, -38.09972, -37.9375, -37.7746, -37.61104, 
    -37.44679, -37.28185, -37.11623, -36.94992, -36.78291, -36.6152, 
    -36.44678, -36.27766, -36.10782, -35.93727, -35.76599, -35.59399, 
    -35.42126, -35.2478, -35.07359, -34.89865, -34.72295, -34.54651, 
    -34.36931, -34.19136, -34.01264, -33.83315, -33.65289, -33.47185, 
    -33.29004, -33.10743, -32.92404, -32.73986, -32.55487, -32.36909, 
    -32.1825, -31.9951, -31.80689, -31.61785, -31.428, -31.23731, -31.0458, 
    -30.85344, -30.66025, -30.46622, -30.27133, -30.07559, -29.879, 
    -29.68154, -29.48322, -29.28403, -29.08397, -28.88303, -28.68121, 
    -28.4785, -28.2749, -28.07041, -27.86502, -27.65873, -27.45154, 
    -27.24343, -27.03441, -26.82448, -26.61362, -26.40184, -26.18913, 
    -25.97548, -25.7609, -25.54539, -25.32892, -25.11152, -24.89316, 
    -24.67384, -24.45357, -24.23234, -24.01015, -23.78698, -23.56285, 
    -23.33775, -23.11166, -22.8846, -22.65655, -22.42752, -22.1975, 
    -21.96649, -21.73449, -21.50148, -21.26748, -21.03248, -20.79647, 
    -20.55946, -20.32143, -20.0824, -19.84235, -19.60129, -19.35921, 
    -19.11611, -18.87199, -18.62685, -18.38068, -18.13349, -17.88527, 
    -17.63603, -17.38575, -17.13445, -16.88211, -16.62874, -16.37434, 
    -16.11891, -15.86244, -15.60494, -15.34641, -15.08684, -14.82624, 
    -14.5646, -14.30193, -14.03823, -13.77349, -13.50773, -13.24093, 
    -12.9731, -12.70425, -12.43437, -12.16346, -11.89153, -11.61857, 
    -11.3446, -11.06961, -10.7936, -10.51658, -10.23855, -9.959517, 
    -9.679476, -9.398433, -9.116391, -8.833357, -8.549331, -8.264318, 
    -7.978323, -7.69135, -7.403402, -7.114486, -6.824605, -6.533765, 
    -6.241971, -5.949229, -5.655543, -5.36092, -5.065367, -4.768888, 
    -4.471492, -4.173184, -3.873971, -3.57386, -3.272859, -2.970974, 
    -2.668215, -2.364588, -2.060102, -1.754765, -1.448585, -1.141572, 
    -0.8337337, -0.52508, -0.2156199, 0.09463693, 0.4056807, 0.7175016, 
    1.030089, 1.343433, 1.657523, 1.972348, 2.287898, 2.60416, 2.921123, 
    3.238777, 3.557109, 3.876107, 4.195758, 4.516052, 4.836975, 5.158514, 
    5.480658, 5.803391, 6.126702, 6.450576, 6.775001, 7.099962, 7.425446, 
    7.751438, 8.077925, 8.404891, 8.732323, 9.060205, 9.388523, 9.717261, 
    10.04641, 10.37594, 10.70585, 11.03612, 11.36673, 11.69768, 12.02893, 
    12.36048, 12.69231, 13.02441, 13.35675, 13.68933, 14.02212, 14.35511, 
    14.68829, 15.02163, 15.35512, 15.68874, 16.02248, 16.35632, 16.69024, 
    17.02423, 17.35827, 17.69234, 18.02642, 18.36051, 18.69457, 19.0286, 
    19.36258, 19.69649, 20.03032, 20.36404, 20.69764, 21.03111, 21.36443, 
    21.69757, 22.03053, 22.36329, 22.69583, 23.02814, 23.3602, 23.69198, 
    24.02349, 24.35469, 24.68559, 25.01615, 25.34636, 25.67621, 26.00569, 
    26.33477, 26.66344, 26.99169, 27.3195, 27.64686, 27.97375, 28.30016, 
    28.62607, 28.95148, 29.27635, 29.60069, 29.92448, 30.2477, 30.57034, 
    30.89239, 31.21383, 31.53465, 31.85485, 32.1744, 32.49329, 32.81152, 
    33.12906, 33.44592, 33.76207, 34.0775, 34.39221, 34.70618, 35.01941, 
    35.33187, 35.64357, 35.95449, 36.26463, 36.57396, 36.88248, 37.19019, 
    37.49707, 37.80312, 38.10832, 38.41267, 38.71616, 39.01879, 39.32053, 
    39.62139, 39.92136, 40.22043, 40.5186, 40.81585, 41.11218, 41.40759, 
    41.70206, 41.9956, 42.28819, 42.57983, 42.87052, 43.16025, 43.44902, 
    43.73681, 44.02363, 44.30947, 44.59433, 44.87819, 45.16107, 45.44296, 
    45.72384, 46.00372, 46.2826, 46.56047, 46.83733, 47.11318, 47.38801, 
    47.66182, 47.93461, 48.20638, 48.47712, 48.74685, 49.01554, 49.2832, 
    49.54984, 49.81544, 50.08001, 50.34355, 50.60606, 50.86753, 51.12797, 
    51.38737, 51.64574, 51.90308, 52.15939, 52.41465, 52.66889, 52.9221, 
    53.17427, 53.42541, 53.67553, 53.92461, 54.17266, 54.41969, 54.6657, 
    54.91068, 55.15463, 55.39757, 55.63949, 55.88039, 56.12028, 56.35915, 
    56.59702, 56.83387, 57.06972, 57.30457, 57.53841, 57.77125, 58.0031, 
    58.23396, 58.46382, 58.69269, 58.92058, 59.14749, 59.37342, 59.59837, 
    59.82235, 60.04536, 60.2674, 60.48848, 60.7086, 60.92776, 61.14597, 
    61.36323, 61.57954, 61.79491, 62.00934, 62.22284, 62.4354, 62.64703, 
    62.85775, 63.06754, 63.27641, 63.48437, 63.69143, 63.89757, 64.10282, 
    64.30717, 64.51063, 64.7132, 64.91487, 65.11568, 65.3156, 65.51466,
  -44.92728, -44.79153, -44.65527, -44.5185, -44.38121, -44.24341, -44.10509, 
    -43.96624, -43.82686, -43.68695, -43.54651, -43.40553, -43.26401, 
    -43.12194, -42.97933, -42.83616, -42.69244, -42.54815, -42.40331, 
    -42.25789, -42.11191, -41.96535, -41.81822, -41.67051, -41.52221, 
    -41.37332, -41.22383, -41.07376, -40.92308, -40.7718, -40.61992, 
    -40.46742, -40.3143, -40.16057, -40.00621, -39.85123, -39.69562, 
    -39.53937, -39.38249, -39.22496, -39.06678, -38.90796, -38.74848, 
    -38.58834, -38.42754, -38.26608, -38.10394, -37.94112, -37.77763, 
    -37.61346, -37.4486, -37.28305, -37.1168, -36.94985, -36.7822, -36.61384, 
    -36.44477, -36.27499, -36.10448, -35.93325, -35.76128, -35.58859, 
    -35.41516, -35.24098, -35.06606, -34.89039, -34.71397, -34.53679, 
    -34.35884, -34.18012, -34.00064, -33.82037, -33.63933, -33.4575, 
    -33.27488, -33.09147, -32.90726, -32.72225, -32.53643, -32.3498, 
    -32.16236, -31.9741, -31.78501, -31.59509, -31.40434, -31.21276, 
    -31.02033, -30.82706, -30.63294, -30.43796, -30.24213, -30.04543, 
    -29.84787, -29.64943, -29.45012, -29.24994, -29.04886, -28.8469, 
    -28.64405, -28.4403, -28.23565, -28.0301, -27.82364, -27.61626, 
    -27.40797, -27.19876, -26.98862, -26.77756, -26.56556, -26.35263, 
    -26.13876, -25.92395, -25.70818, -25.49147, -25.2738, -25.05518, 
    -24.83559, -24.61503, -24.39351, -24.17102, -23.94755, -23.7231, 
    -23.49767, -23.27125, -23.04384, -22.81544, -22.58605, -22.35566, 
    -22.12427, -21.89188, -21.65848, -21.42407, -21.18865, -20.95221, 
    -20.71476, -20.47629, -20.2368, -19.99629, -19.75475, -19.51218, 
    -19.26858, -19.02395, -18.77829, -18.5316, -18.28386, -18.0351, 
    -17.78529, -17.53444, -17.28255, -17.02962, -16.77564, -16.52062, 
    -16.26456, -16.00745, -15.74929, -15.49009, -15.22985, -14.96855, 
    -14.70622, -14.44283, -14.1784, -13.91293, -13.64641, -13.37885, 
    -13.11025, -12.84061, -12.56992, -12.2982, -12.02544, -11.75165, 
    -11.47683, -11.20097, -10.92409, -10.64618, -10.36724, -10.08729, 
    -9.806318, -9.524332, -9.241335, -8.95733, -8.672321, -8.386312, 
    -8.099308, -7.811312, -7.522329, -7.232363, -6.941419, -6.649503, 
    -6.35662, -6.062775, -5.767973, -5.472221, -5.175525, -4.877891, 
    -4.579325, -4.279835, -3.979426, -3.678107, -3.375884, -3.072765, 
    -2.768758, -2.463871, -2.158111, -1.851488, -1.544009, -1.235684, 
    -0.9265221, -0.6165318, -0.3057229, 0.005895053, 0.3183122, 0.6315184, 
    0.9455033, 1.260257, 1.575767, 1.892025, 2.209018, 2.526735, 2.845165, 
    3.164296, 3.484116, 3.804613, 4.125774, 4.447588, 4.770041, 5.093121, 
    5.416813, 5.741107, 6.065986, 6.391439, 6.717451, 7.044009, 7.371098, 
    7.698703, 8.026812, 8.355408, 8.684476, 9.014004, 9.343974, 9.674372, 
    10.00518, 10.33639, 10.66798, 10.99993, 11.33224, 11.66488, 11.99783, 
    12.33109, 12.66464, 12.99845, 13.33251, 13.66682, 14.00134, 14.33606, 
    14.67097, 15.00605, 15.34128, 15.67664, 16.01213, 16.34771, 16.68338, 
    17.01912, 17.35491, 17.69073, 18.02656, 18.3624, 18.69821, 19.03399, 
    19.36972, 19.70538, 20.04095, 20.37641, 20.71176, 21.04697, 21.38202, 
    21.7169, 22.05159, 22.38608, 22.72034, 23.05437, 23.38814, 23.72164, 
    24.05485, 24.38776, 24.72035, 25.0526, 25.3845, 25.71603, 26.04717, 
    26.37792, 26.70825, 27.03815, 27.36761, 27.6966, 28.02512, 28.35315, 
    28.68068, 29.00768, 29.33415, 29.66008, 29.98544, 30.31023, 30.63443, 
    30.95803, 31.28101, 31.60336, 31.92507, 32.24613, 32.56652, 32.88623, 
    33.20525, 33.52357, 33.84118, 34.15805, 34.47419, 34.78958, 35.10421, 
    35.41808, 35.73116, 36.04345, 36.35494, 36.66562, 36.97548, 37.28451, 
    37.5927, 37.90005, 38.20654, 38.51216, 38.81691, 39.12077, 39.42375, 
    39.72583, 40.02701, 40.32727, 40.62661, 40.92503, 41.22252, 41.51907, 
    41.81467, 42.10932, 42.40302, 42.69574, 42.98751, 43.2783, 43.56811, 
    43.85693, 44.14478, 44.43162, 44.71747, 45.00232, 45.28617, 45.569, 
    45.85083, 46.13164, 46.41143, 46.69021, 46.96796, 47.24467, 47.52037, 
    47.79503, 48.06866, 48.34126, 48.61281, 48.88333, 49.15281, 49.42125, 
    49.68864, 49.95499, 50.2203, 50.48457, 50.74778, 51.00996, 51.27108, 
    51.53116, 51.7902, 52.04819, 52.30513, 52.56103, 52.81588, 53.06969, 
    53.32246, 53.57419, 53.82487, 54.07452, 54.32312, 54.57069, 54.81722, 
    55.06272, 55.30719, 55.55062, 55.79302, 56.0344, 56.27475, 56.51408, 
    56.75239, 56.98968, 57.22596, 57.46122, 57.69547, 57.92871, 58.16094, 
    58.39217, 58.62241, 58.85164, 59.07988, 59.30713, 59.53339, 59.75867, 
    59.98296, 60.20628, 60.42862, 60.64999, 60.87039, 61.08982, 61.3083, 
    61.52581, 61.74238, 61.95799, 62.17265, 62.38638, 62.59916, 62.81101, 
    63.02192, 63.23191, 63.44098, 63.64912, 63.85635, 64.06267, 64.26808, 
    64.47259, 64.67619, 64.87891, 65.08073, 65.28166, 65.48171, 65.68088,
  -45.08842, -44.95283, -44.81674, -44.68014, -44.54302, -44.40538, 
    -44.26722, -44.12854, -43.98932, -43.84957, -43.70929, -43.56847, 
    -43.4271, -43.28519, -43.14272, -42.99971, -42.85614, -42.712, -42.5673, 
    -42.42204, -42.2762, -42.12978, -41.98279, -41.83521, -41.68705, 
    -41.5383, -41.38895, -41.23901, -41.08846, -40.93731, -40.78555, 
    -40.63317, -40.48018, -40.32657, -40.17233, -40.01746, -39.86197, 
    -39.70583, -39.54905, -39.39163, -39.23356, -39.07483, -38.91545, 
    -38.75541, -38.59471, -38.43333, -38.27128, -38.10855, -37.94514, 
    -37.78105, -37.61627, -37.45079, -37.28461, -37.11773, -36.95015, 
    -36.78185, -36.61284, -36.44311, -36.27265, -36.10147, -35.92955, 
    -35.7569, -35.5835, -35.40936, -35.23447, -35.05883, -34.88243, 
    -34.70526, -34.52733, -34.34863, -34.16915, -33.98888, -33.80784, 
    -33.626, -33.44337, -33.25995, -33.07572, -32.89069, -32.70484, 
    -32.51817, -32.33069, -32.14238, -31.95325, -31.76328, -31.57247, 
    -31.38082, -31.18832, -30.99498, -30.80077, -30.60571, -30.40979, 
    -30.21299, -30.01532, -29.81678, -29.61736, -29.41704, -29.21584, 
    -29.01375, -28.81075, -28.60686, -28.40206, -28.19634, -27.98971, 
    -27.78217, -27.5737, -27.3643, -27.15397, -26.9427, -26.7305, -26.51735, 
    -26.30325, -26.08821, -25.8722, -25.65524, -25.43732, -25.21843, 
    -24.99857, -24.77774, -24.55593, -24.33314, -24.10936, -23.8846, 
    -23.65885, -23.4321, -23.20435, -22.97561, -22.74586, -22.5151, 
    -22.28333, -22.05055, -21.81676, -21.58194, -21.34611, -21.10925, 
    -20.87136, -20.63245, -20.3925, -20.15152, -19.90951, -19.66645, 
    -19.42236, -19.17723, -18.93105, -18.68382, -18.43555, -18.18623, 
    -17.93586, -17.68444, -17.43196, -17.17844, -16.92385, -16.66822, 
    -16.41152, -16.15377, -15.89496, -15.63509, -15.37417, -15.11219, 
    -14.84915, -14.58505, -14.31989, -14.05368, -13.78641, -13.51808, 
    -13.2487, -12.97827, -12.70678, -12.43425, -12.16066, -11.88603, 
    -11.61035, -11.33362, -11.05586, -10.77705, -10.49721, -10.21634, 
    -9.93443, -9.651496, -9.367537, -9.082558, -8.796561, -8.509551, 
    -8.221531, -7.932506, -7.642481, -7.351459, -7.059446, -6.766447, 
    -6.472467, -6.177512, -5.881587, -5.584698, -5.286851, -4.988052, 
    -4.688309, -4.387627, -4.086014, -3.783477, -3.480023, -3.175659, 
    -2.870394, -2.564236, -2.257192, -1.949272, -1.640483, -1.330836, 
    -1.020338, -0.7089992, -0.3968292, -0.08383764, 0.2299655, 0.5445699, 
    0.8599654, 1.176141, 1.493087, 1.81079, 2.129241, 2.448428, 2.768339, 
    3.088962, 3.410286, 3.732297, 4.054984, 4.378333, 4.702332, 5.026968, 
    5.352227, 5.678096, 6.004562, 6.331611, 6.659227, 6.987399, 7.316111, 
    7.645348, 7.975095, 8.305339, 8.636065, 8.967255, 9.298897, 9.630973, 
    9.963469, 10.29637, 10.62966, 10.96332, 11.29733, 11.63169, 11.96637, 
    12.30135, 12.63663, 12.97218, 13.30798, 13.64403, 13.9803, 14.31677, 
    14.65344, 14.99028, 15.32727, 15.6644, 16.00165, 16.339, 16.67644, 
    17.01395, 17.3515, 17.68909, 18.0267, 18.36431, 18.70189, 19.03945, 
    19.37694, 19.71437, 20.05171, 20.38894, 20.72605, 21.06302, 21.39983, 
    21.73646, 22.07291, 22.40914, 22.74515, 23.08092, 23.41643, 23.75166, 
    24.0866, 24.42122, 24.75553, 25.08949, 25.42309, 25.75632, 26.08915, 
    26.42159, 26.75359, 27.08517, 27.41628, 27.74693, 28.0771, 28.40677, 
    28.73592, 29.06455, 29.39263, 29.72016, 30.04712, 30.37349, 30.69926, 
    31.02443, 31.34896, 31.67286, 31.99611, 32.31868, 32.64059, 32.9618, 
    33.28231, 33.60211, 33.92118, 34.23951, 34.5571, 34.87392, 35.18998, 
    35.50525, 35.81973, 36.1334, 36.44626, 36.7583, 37.06951, 37.37988, 
    37.68938, 37.99804, 38.30582, 38.61272, 38.91874, 39.22387, 39.52808, 
    39.83139, 40.13379, 40.43525, 40.73579, 41.03538, 41.33403, 41.63173, 
    41.92846, 42.22423, 42.51904, 42.81286, 43.10571, 43.39756, 43.68842, 
    43.97829, 44.26716, 44.55502, 44.84187, 45.1277, 45.41252, 45.69632, 
    45.97909, 46.26083, 46.54155, 46.82122, 47.09986, 47.37746, 47.65402, 
    47.92954, 48.20401, 48.47743, 48.7498, 49.02112, 49.29139, 49.5606, 
    49.82876, 50.09586, 50.3619, 50.6269, 50.89083, 51.1537, 51.41552, 
    51.67627, 51.93597, 52.19461, 52.4522, 52.70872, 52.9642, 53.21861, 
    53.47197, 53.72428, 53.97554, 54.22574, 54.4749, 54.723, 54.97006, 
    55.21607, 55.46104, 55.70497, 55.94786, 56.18971, 56.43053, 56.67031, 
    56.90906, 57.14679, 57.38348, 57.61916, 57.85381, 58.08744, 58.32006, 
    58.55167, 58.78226, 59.01186, 59.24044, 59.46803, 59.69462, 59.92022, 
    60.14482, 60.36845, 60.59108, 60.81274, 61.03341, 61.25312, 61.47186, 
    61.68963, 61.90644, 62.12229, 62.33718, 62.55113, 62.76413, 62.97618, 
    63.1873, 63.39748, 63.60674, 63.81506, 64.02246, 64.22894, 64.43452, 
    64.63918, 64.84293, 65.04578, 65.24773, 65.44879, 65.64896, 65.84824,
  -45.25026, -45.11485, -44.97893, -44.8425, -44.70555, -44.56808, -44.43009, 
    -44.29157, -44.15252, -44.01294, -43.87281, -43.73215, -43.59095, 
    -43.44919, -43.30689, -43.16403, -43.02061, -42.87663, -42.73208, 
    -42.58696, -42.44127, -42.29501, -42.14816, -42.00072, -41.8527, 
    -41.70409, -41.55488, -41.40508, -41.25466, -41.10365, -40.95201, 
    -40.79977, -40.6469, -40.49341, -40.3393, -40.18455, -40.02917, 
    -39.87315, -39.71649, -39.55918, -39.40121, -39.2426, -39.08332, 
    -38.92338, -38.76277, -38.60149, -38.43954, -38.2769, -38.11358, 
    -37.94957, -37.78487, -37.61947, -37.45337, -37.28656, -37.11905, 
    -36.95082, -36.78187, -36.6122, -36.4418, -36.27067, -36.0988, -35.92619, 
    -35.75284, -35.57874, -35.40389, -35.22828, -35.0519, -34.87476, 
    -34.69685, -34.51816, -34.33869, -34.15844, -33.97739, -33.79556, 
    -33.61292, -33.42949, -33.24524, -33.06018, -32.87431, -32.68762, 
    -32.50011, -32.31176, -32.12258, -31.93256, -31.7417, -31.54999, 
    -31.35743, -31.16401, -30.96973, -30.77459, -30.57858, -30.38169, 
    -30.18392, -29.98528, -29.78574, -29.58531, -29.38399, -29.18176, 
    -28.97863, -28.7746, -28.56964, -28.36378, -28.15699, -27.94927, 
    -27.74062, -27.53104, -27.32052, -27.10906, -26.89665, -26.68329, 
    -26.46897, -26.2537, -26.03746, -25.82026, -25.60208, -25.38293, 
    -25.16281, -24.9417, -24.7196, -24.49652, -24.27244, -24.04737, -23.8213, 
    -23.59422, -23.36614, -23.13705, -22.90695, -22.67583, -22.44369, 
    -22.21052, -21.97634, -21.74112, -21.50487, -21.26759, -21.02927, 
    -20.78992, -20.54952, -20.30808, -20.06559, -19.82205, -19.57746, 
    -19.33182, -19.08513, -18.83738, -18.58857, -18.3387, -18.08777, 
    -17.83577, -17.58272, -17.32859, -17.0734, -16.81715, -16.55982, 
    -16.30143, -16.04196, -15.78143, -15.51983, -15.25715, -14.99341, 
    -14.7286, -14.46271, -14.19576, -13.92773, -13.65864, -13.38848, 
    -13.11726, -12.84496, -12.57161, -12.29719, -12.02171, -11.74517, 
    -11.46758, -11.18893, -10.90923, -10.62847, -10.34667, -10.06383, 
    -9.779943, -9.495018, -9.209059, -8.922069, -8.634051, -8.345011, 
    -8.054951, -7.763877, -7.471793, -7.178704, -6.884615, -6.589532, 
    -6.293459, -5.996402, -5.698368, -5.399363, -5.099391, -4.798461, 
    -4.49658, -4.193753, -3.889988, -3.585293, -3.279675, -2.973142, 
    -2.665703, -2.357364, -2.048136, -1.738026, -1.427044, -1.115198, 
    -0.8024991, -0.4889557, -0.174578, 0.1406239, 0.4566398, 0.7734591, 
    1.091071, 1.409465, 1.728629, 2.048553, 2.369224, 2.69063, 3.012761, 
    3.335603, 3.659144, 3.983372, 4.308273, 4.633834, 4.960043, 5.286886, 
    5.614348, 5.942417, 6.271079, 6.600318, 6.930121, 7.260473, 7.59136, 
    7.922766, 8.254676, 8.587076, 8.91995, 9.253282, 9.587055, 9.921256, 
    10.25587, 10.59087, 10.92626, 11.26201, 11.5981, 11.93452, 12.27125, 
    12.60828, 12.94559, 13.28316, 13.62097, 13.95901, 14.29726, 14.6357, 
    14.97431, 15.31309, 15.652, 15.99104, 16.33018, 16.66941, 17.00871, 
    17.34806, 17.68744, 18.02684, 18.36624, 18.70562, 19.04497, 19.38425, 
    19.72347, 20.0626, 20.40162, 20.74051, 21.07926, 21.41785, 21.75626, 
    22.09448, 22.43248, 22.77026, 23.10779, 23.44505, 23.78203, 24.11872, 
    24.45509, 24.79113, 25.12682, 25.46214, 25.79709, 26.13164, 26.46577, 
    26.79948, 27.13274, 27.46554, 27.79786, 28.12969, 28.46102, 28.79182, 
    29.12209, 29.4518, 29.78095, 30.10952, 30.43749, 30.76486, 31.0916, 
    31.41771, 31.74317, 32.06796, 32.39208, 32.71551, 33.03824, 33.36026, 
    33.68155, 34.00211, 34.32191, 34.64095, 34.95922, 35.27671, 35.5934, 
    35.90929, 36.22436, 36.53861, 36.85202, 37.16459, 37.47629, 37.78714, 
    38.09711, 38.4062, 38.71439, 39.02169, 39.32808, 39.63355, 39.9381, 
    40.24172, 40.5444, 40.84613, 41.1469, 41.44672, 41.74558, 42.04346, 
    42.34036, 42.63628, 42.9312, 43.22513, 43.51806, 43.80999, 44.1009, 
    44.3908, 44.67968, 44.96753, 45.25436, 45.54016, 45.82492, 46.10864, 
    46.39132, 46.67295, 46.95354, 47.23308, 47.51156, 47.78899, 48.06536, 
    48.34067, 48.61492, 48.88811, 49.16023, 49.43129, 49.70128, 49.9702, 
    50.23806, 50.50484, 50.77056, 51.0352, 51.29877, 51.56128, 51.82272, 
    52.08308, 52.34237, 52.6006, 52.85775, 53.11384, 53.36886, 53.62281, 
    53.87571, 54.12753, 54.37829, 54.62799, 54.87664, 55.12422, 55.37075, 
    55.61622, 55.86065, 56.10402, 56.34634, 56.58762, 56.82785, 57.06704, 
    57.30519, 57.54231, 57.7784, 58.01345, 58.24747, 58.48048, 58.71245, 
    58.94341, 59.17336, 59.40229, 59.63021, 59.85713, 60.08304, 60.30796, 
    60.53188, 60.7548, 60.97674, 61.19769, 61.41766, 61.63666, 61.85468, 
    62.07173, 62.28782, 62.50294, 62.7171, 62.93031, 63.14257, 63.35388, 
    63.56425, 63.77369, 63.98219, 64.18976, 64.3964, 64.60213, 64.80693, 
    65.01083, 65.21381, 65.41589, 65.61707, 65.81736, 66.01675,
  -45.41282, -45.27758, -45.14184, -45.00558, -44.86881, -44.73151, 
    -44.59369, -44.45534, -44.31646, -44.17704, -44.03709, -43.8966, 
    -43.75555, -43.61396, -43.47182, -43.32912, -43.18586, -43.04203, 
    -42.89764, -42.75268, -42.60714, -42.46103, -42.31433, -42.16705, 
    -42.01917, -41.8707, -41.72164, -41.57197, -41.4217, -41.27082, 
    -41.11932, -40.96721, -40.81447, -40.66111, -40.50713, -40.3525, 
    -40.19725, -40.04135, -39.8848, -39.72761, -39.56976, -39.41125, 
    -39.25208, -39.09225, -38.93175, -38.77057, -38.60871, -38.44617, 
    -38.28294, -38.11902, -37.95441, -37.78909, -37.62307, -37.45634, 
    -37.2889, -37.12075, -36.95187, -36.78226, -36.61192, -36.44085, 
    -36.26904, -36.09648, -35.92318, -35.74912, -35.57431, -35.39873, 
    -35.22239, -35.04528, -34.86739, -34.68872, -34.50927, -34.32903, 
    -34.14799, -33.96616, -33.78353, -33.60009, -33.41583, -33.23076, 
    -33.04487, -32.85816, -32.67061, -32.48223, -32.29301, -32.10295, 
    -31.91204, -31.72028, -31.52765, -31.33417, -31.13982, -30.9446, 
    -30.74851, -30.55153, -30.35368, -30.15493, -29.95529, -29.75475, 
    -29.5533, -29.35096, -29.1477, -28.94352, -28.73843, -28.53241, 
    -28.32546, -28.11758, -27.90876, -27.699, -27.48829, -27.27664, 
    -27.06403, -26.85046, -26.63593, -26.42043, -26.20396, -25.98652, 
    -25.7681, -25.54869, -25.3283, -25.10693, -24.88455, -24.66118, 
    -24.43681, -24.21143, -23.98504, -23.75764, -23.52923, -23.2998, 
    -23.06934, -22.83786, -22.60535, -22.37181, -22.13723, -21.90161, 
    -21.66496, -21.42726, -21.18851, -20.94871, -20.70786, -20.46596, 
    -20.223, -19.97898, -19.7339, -19.48776, -19.24055, -18.99228, -18.74293, 
    -18.49251, -18.24102, -17.98846, -17.73482, -17.4801, -17.2243, 
    -16.96743, -16.70947, -16.45044, -16.19032, -15.92912, -15.66684, 
    -15.40347, -15.13902, -14.87349, -14.60688, -14.33918, -14.07041, 
    -13.80054, -13.5296, -13.25758, -12.98449, -12.71031, -12.43506, 
    -12.15873, -11.88133, -11.60286, -11.32332, -11.04272, -10.76105, 
    -10.47832, -10.19453, -9.90969, -9.623796, -9.336851, -9.048862, 
    -8.759832, -8.469766, -8.178665, -7.886537, -7.593384, -7.299213, 
    -7.004027, -6.707833, -6.410635, -6.11244, -5.813252, -5.51308, 
    -5.211927, -4.909802, -4.606711, -4.302662, -3.99766, -3.691714, 
    -3.384832, -3.07702, -2.768289, -2.458645, -2.148097, -1.836654, 
    -1.524326, -1.211121, -0.8970492, -0.5821201, -0.2663435, 0.05027031, 
    0.3677109, 0.6859676, 1.00503, 1.324886, 1.645525, 1.966935, 2.289105, 
    2.612023, 2.935676, 3.260053, 3.58514, 3.910924, 4.237393, 4.564534, 
    4.892332, 5.220775, 5.549848, 5.879538, 6.20983, 6.540709, 6.872162, 
    7.204174, 7.536728, 7.869812, 8.203407, 8.537501, 8.872076, 9.207118, 
    9.542609, 9.878535, 10.21488, 10.55162, 10.88875, 11.22625, 11.5641, 
    11.90228, 12.24079, 12.57959, 12.91867, 13.25803, 13.59762, 13.93746, 
    14.2775, 14.61774, 14.95816, 15.29874, 15.63946, 15.9803, 16.32125, 
    16.6623, 17.00341, 17.34457, 17.68577, 18.02699, 18.3682, 18.7094, 
    19.05055, 19.39165, 19.73268, 20.07362, 20.41445, 20.75515, 21.0957, 
    21.43609, 21.7763, 22.11631, 22.45611, 22.79567, 23.13498, 23.47402, 
    23.81278, 24.15123, 24.48936, 24.82716, 25.1646, 25.50167, 25.83835, 
    26.17463, 26.51049, 26.84591, 27.18088, 27.51538, 27.8494, 28.18291, 
    28.51591, 28.84838, 29.18031, 29.51167, 29.84246, 30.17265, 30.50225, 
    30.83122, 31.15956, 31.48726, 31.81429, 32.14066, 32.46633, 32.79131, 
    33.11557, 33.43911, 33.76191, 34.08396, 34.40525, 34.72576, 35.04549, 
    35.36443, 35.68256, 35.99987, 36.31635, 36.63199, 36.94679, 37.26072, 
    37.57379, 37.88598, 38.19728, 38.50769, 38.81718, 39.12577, 39.43344, 
    39.74017, 40.04597, 40.35082, 40.65472, 40.95766, 41.25963, 41.56063, 
    41.86065, 42.15968, 42.45771, 42.75475, 43.05079, 43.34581, 43.63982, 
    43.93282, 44.22478, 44.51572, 44.80562, 45.09449, 45.38231, 45.66909, 
    45.95482, 46.23949, 46.52311, 46.80568, 47.08718, 47.36761, 47.64698, 
    47.92528, 48.20251, 48.47867, 48.75375, 49.02776, 49.30069, 49.57254, 
    49.8433, 50.11299, 50.3816, 50.64912, 50.91557, 51.18093, 51.44521, 
    51.7084, 51.97051, 52.23154, 52.49149, 52.75035, 53.00813, 53.26484, 
    53.52046, 53.77501, 54.02848, 54.28087, 54.5322, 54.78244, 55.03162, 
    55.27973, 55.52677, 55.77274, 56.01765, 56.26151, 56.5043, 56.74603, 
    56.98671, 57.22635, 57.46492, 57.70246, 57.93895, 58.1744, 58.40882, 
    58.6422, 58.87454, 59.10586, 59.33615, 59.56543, 59.79368, 60.02092, 
    60.24715, 60.47237, 60.69658, 60.91979, 61.14201, 61.36323, 61.58347, 
    61.80272, 62.02098, 62.23827, 62.45458, 62.66993, 62.8843, 63.09772, 
    63.31018, 63.52169, 63.73224, 63.94185, 64.15052, 64.35825, 64.56506, 
    64.77093, 64.97588, 65.17991, 65.38303, 65.58523, 65.78653, 65.98692, 
    66.18642,
  -45.57609, -45.44104, -45.30547, -45.1694, -45.0328, -44.89568, -44.75803, 
    -44.61986, -44.48115, -44.34191, -44.20213, -44.0618, -43.92093, 
    -43.7795, -43.63752, -43.49499, -43.35189, -43.20823, -43.064, -42.9192, 
    -42.77382, -42.62786, -42.48131, -42.33418, -42.18646, -42.03814, 
    -41.88922, -41.7397, -41.58957, -41.43883, -41.28747, -41.1355, -40.9829, 
    -40.82967, -40.67582, -40.52133, -40.3662, -40.21042, -40.054, -39.89693, 
    -39.7392, -39.58081, -39.42175, -39.26203, -39.10163, -38.94056, 
    -38.7788, -38.61636, -38.45324, -38.28941, -38.12489, -37.95966, 
    -37.79373, -37.62708, -37.45972, -37.29164, -37.12284, -36.9533, 
    -36.78303, -36.61202, -36.44027, -36.26777, -36.09452, -35.92051, 
    -35.74574, -35.57021, -35.39391, -35.21683, -35.03897, -34.86033, 
    -34.6809, -34.50068, -34.31966, -34.13783, -33.9552, -33.77176, -33.5875, 
    -33.40242, -33.21652, -33.02979, -32.84222, -32.65381, -32.46455, 
    -32.27446, -32.0835, -31.89169, -31.69901, -31.50547, -31.31106, 
    -31.11577, -30.91959, -30.72254, -30.52459, -30.32575, -30.12601, 
    -29.92536, -29.7238, -29.52134, -29.31795, -29.11364, -28.90841, 
    -28.70224, -28.49514, -28.2871, -28.07812, -27.86818, -27.6573, 
    -27.44545, -27.23265, -27.01888, -26.80413, -26.58842, -26.37172, 
    -26.15405, -25.93538, -25.71573, -25.49508, -25.27343, -25.05078, 
    -24.82713, -24.60246, -24.37678, -24.15008, -23.92237, -23.69362, 
    -23.46385, -23.23305, -23.00121, -22.76833, -22.53441, -22.29945, 
    -22.06344, -21.82638, -21.58826, -21.34908, -21.10885, -20.86756, 
    -20.6252, -20.38177, -20.13727, -19.8917, -19.64506, -19.39733, 
    -19.14853, -18.89865, -18.64769, -18.39564, -18.14251, -17.88828, 
    -17.63297, -17.37657, -17.11908, -16.8605, -16.60082, -16.34005, 
    -16.07818, -15.81522, -15.55116, -15.28601, -15.01976, -14.75242, 
    -14.48398, -14.21444, -13.94381, -13.67209, -13.39927, -13.12536, 
    -12.85036, -12.57428, -12.2971, -12.01884, -11.73949, -11.45906, 
    -11.17755, -10.89496, -10.6113, -10.32656, -10.04076, -9.753889, 
    -9.465956, -9.176964, -8.886915, -8.595817, -8.30367, -8.01048, 
    -7.716253, -7.420992, -7.124702, -6.82739, -6.529059, -6.229717, 
    -5.929369, -5.628021, -5.325679, -5.02235, -4.718041, -4.412759, 
    -4.106511, -3.799304, -3.491147, -3.182047, -2.872013, -2.561052, 
    -2.249174, -1.936387, -1.622701, -1.308125, -0.9926676, -0.6763399, 
    -0.3591516, -0.04111278, 0.2777659, 0.5974737, 0.9179996, 1.239333, 
    1.561461, 1.884373, 2.208057, 2.532501, 2.857693, 3.183619, 3.510268, 
    3.837626, 4.165679, 4.494416, 4.823821, 5.153882, 5.484583, 5.815911, 
    6.147851, 6.48039, 6.813511, 7.1472, 7.481441, 7.816221, 8.151522, 
    8.487329, 8.823626, 9.160397, 9.497625, 9.835296, 10.17339, 10.5119, 
    10.85079, 11.19006, 11.52969, 11.86966, 12.20995, 12.55055, 12.89143, 
    13.23259, 13.574, 13.91564, 14.2575, 14.59956, 14.9418, 15.28421, 
    15.62676, 15.96943, 16.31222, 16.65509, 16.99804, 17.34104, 17.68408, 
    18.02713, 18.37018, 18.71322, 19.05621, 19.39915, 19.74201, 20.08478, 
    20.42744, 20.76997, 21.11234, 21.45456, 21.79659, 22.13842, 22.48003, 
    22.8214, 23.16251, 23.50335, 23.8439, 24.18414, 24.52406, 24.86363, 
    25.20284, 25.54168, 25.88012, 26.21815, 26.55575, 26.89291, 27.2296, 
    27.56582, 27.90155, 28.23677, 28.57147, 28.90562, 29.23922, 29.57225, 
    29.9047, 30.23654, 30.56777, 30.89837, 31.22833, 31.55763, 31.88626, 
    32.2142, 32.54145, 32.86798, 33.19379, 33.51887, 33.84319, 34.16676, 
    34.48955, 34.81155, 35.13276, 35.45315, 35.77273, 36.09148, 36.40938, 
    36.72644, 37.04263, 37.35794, 37.67238, 37.98592, 38.29857, 38.6103, 
    38.92112, 39.231, 39.53996, 39.84796, 40.15502, 40.46111, 40.76624, 
    41.0704, 41.37357, 41.67575, 41.97694, 42.27713, 42.57632, 42.87449, 
    43.17164, 43.46777, 43.76286, 44.05693, 44.34995, 44.64193, 44.93287, 
    45.22275, 45.51157, 45.79934, 46.08604, 46.37168, 46.65624, 46.93974, 
    47.22215, 47.50349, 47.78375, 48.06293, 48.34101, 48.61802, 48.89394, 
    49.16877, 49.4425, 49.71515, 49.98669, 50.25715, 50.52651, 50.79478, 
    51.06195, 51.32803, 51.593, 51.85689, 52.11967, 52.38137, 52.64197, 
    52.90147, 53.15989, 53.4172, 53.67343, 53.92857, 54.18262, 54.43558, 
    54.68746, 54.93825, 55.18796, 55.43659, 55.68414, 55.93062, 56.17602, 
    56.42035, 56.6636, 56.9058, 57.14692, 57.38699, 57.626, 57.86395, 
    58.10084, 58.33669, 58.57148, 58.80524, 59.03795, 59.26963, 59.50026, 
    59.72987, 59.95845, 60.18601, 60.41255, 60.63807, 60.86257, 61.08607, 
    61.30856, 61.53005, 61.75054, 61.97004, 62.18855, 62.40607, 62.6226, 
    62.83817, 63.05275, 63.26637, 63.47903, 63.69072, 63.90145, 64.11124, 
    64.32008, 64.52796, 64.73492, 64.94093, 65.14602, 65.35018, 65.55342, 
    65.75574, 65.95716, 66.15766, 66.35726,
  -45.74008, -45.60521, -45.46983, -45.33393, -45.19752, -45.06058, 
    -44.92311, -44.78512, -44.64659, -44.50753, -44.36792, -44.22776, 
    -44.08707, -43.94581, -43.80401, -43.66164, -43.51871, -43.37522, 
    -43.23115, -43.08651, -42.94129, -42.79549, -42.64911, -42.50213, 
    -42.35456, -42.2064, -42.05763, -41.90826, -41.75828, -41.60769, 
    -41.45647, -41.30464, -41.15219, -40.9991, -40.84538, -40.69102, 
    -40.53603, -40.38038, -40.22409, -40.06714, -39.90953, -39.75126, 
    -39.59233, -39.43272, -39.27244, -39.11148, -38.94983, -38.78749, 
    -38.62447, -38.46074, -38.29632, -38.13119, -37.96535, -37.79879, 
    -37.63151, -37.46351, -37.29478, -37.12532, -36.95513, -36.78419, 
    -36.6125, -36.44007, -36.26687, -36.09292, -35.91821, -35.74272, 
    -35.56646, -35.38942, -35.21159, -35.03299, -34.85358, -34.67338, 
    -34.49238, -34.31057, -34.12795, -33.94452, -33.76026, -33.57518, 
    -33.38926, -33.20252, -33.01493, -32.8265, -32.63722, -32.44709, 
    -32.25609, -32.06424, -31.87151, -31.67792, -31.48344, -31.28809, 
    -31.09184, -30.89471, -30.69668, -30.49775, -30.29791, -30.09716, 
    -29.8955, -29.69291, -29.48941, -29.28498, -29.07961, -28.8733, 
    -28.66605, -28.45786, -28.24871, -28.03861, -27.82755, -27.61552, 
    -27.40252, -27.18855, -26.9736, -26.75768, -26.54076, -26.32285, 
    -26.10395, -25.88405, -25.66315, -25.44124, -25.21832, -24.99438, 
    -24.76942, -24.54345, -24.31644, -24.08841, -23.85934, -23.62923, 
    -23.39808, -23.16589, -22.93265, -22.69836, -22.46301, -22.22661, 
    -21.98915, -21.75062, -21.51102, -21.27035, -21.02861, -20.7858, 
    -20.5419, -20.29693, -20.05087, -19.80372, -19.55549, -19.30617, 
    -19.05576, -18.80425, -18.55164, -18.29794, -18.04314, -17.78723, 
    -17.53023, -17.27212, -17.01291, -16.75259, -16.49116, -16.22863, 
    -15.96499, -15.70024, -15.43438, -15.16741, -14.89934, -14.63016, 
    -14.35986, -14.08846, -13.81596, -13.54234, -13.26762, -12.9918, 
    -12.71487, -12.43684, -12.15771, -11.87748, -11.59616, -11.31374, 
    -11.03023, -10.74563, -10.45994, -10.17317, -9.88532, -9.596392, 
    -9.306391, -9.01532, -8.723182, -8.429983, -8.135727, -7.840418, 
    -7.544061, -7.246661, -6.948223, -6.648753, -6.348256, -6.046739, 
    -5.744207, -5.440667, -5.136126, -4.830589, -4.524065, -4.216561, 
    -3.908084, -3.598642, -3.288242, -2.976894, -2.664606, -2.351386, 
    -2.037243, -1.722187, -1.406227, -1.089373, -0.7716336, -0.4530204, 
    -0.1335433, 0.1867871, 0.5079599, 0.829964, 1.152788, 1.47642, 1.800849, 
    2.126063, 2.452049, 2.778795, 3.106287, 3.434514, 3.763462, 4.093117, 
    4.423466, 4.754496, 5.086191, 5.418538, 5.751523, 6.08513, 6.419345, 
    6.754154, 7.08954, 7.425487, 7.761981, 8.099007, 8.436546, 8.774586, 
    9.113107, 9.452093, 9.791529, 10.1314, 10.47168, 10.81236, 11.15343, 
    11.49485, 11.83663, 12.17873, 12.52115, 12.86385, 13.20683, 13.55008, 
    13.89355, 14.23725, 14.58116, 14.92525, 15.2695, 15.6139, 15.95843, 
    16.30307, 16.6478, 16.99261, 17.33747, 17.68237, 18.02728, 18.37219, 
    18.71708, 19.06194, 19.40673, 19.75145, 20.09608, 20.44059, 20.78497, 
    21.1292, 21.47326, 21.81713, 22.16079, 22.50424, 22.84744, 23.19038, 
    23.53304, 23.8754, 24.21746, 24.55918, 24.90055, 25.24155, 25.58217, 
    25.92239, 26.26219, 26.60156, 26.94047, 27.27892, 27.61688, 27.95434, 
    28.29128, 28.62769, 28.96355, 29.29885, 29.63356, 29.96768, 30.30119, 
    30.63408, 30.96632, 31.29791, 31.62884, 31.95908, 32.28862, 32.61745, 
    32.94556, 33.27294, 33.59957, 33.92543, 34.25052, 34.57483, 34.89833, 
    35.22103, 35.5429, 35.86394, 36.18414, 36.50348, 36.82195, 37.13955, 
    37.45626, 37.77208, 38.087, 38.40099, 38.71407, 39.02621, 39.33741, 
    39.64766, 39.95694, 40.26527, 40.57262, 40.87899, 41.18436, 41.48875, 
    41.79213, 42.0945, 42.39586, 42.69619, 42.9955, 43.29377, 43.59101, 
    43.8872, 44.18234, 44.47643, 44.76946, 45.06143, 45.35234, 45.64217, 
    45.93092, 46.21861, 46.5052, 46.79072, 47.07515, 47.35848, 47.64073, 
    47.92188, 48.20193, 48.48089, 48.75875, 49.0355, 49.31115, 49.5857, 
    49.85913, 50.13147, 50.40269, 50.67281, 50.94182, 51.20972, 51.47651, 
    51.74219, 52.00677, 52.27023, 52.53259, 52.79384, 53.05398, 53.31302, 
    53.57096, 53.82779, 54.08352, 54.33814, 54.59167, 54.8441, 55.09544, 
    55.34568, 55.59483, 55.84289, 56.08986, 56.33575, 56.58055, 56.82428, 
    57.06692, 57.30849, 57.54899, 57.78842, 58.02678, 58.26408, 58.50031, 
    58.73549, 58.96962, 59.20269, 59.43472, 59.6657, 59.89564, 60.12455, 
    60.35242, 60.57926, 60.80508, 61.02987, 61.25365, 61.47641, 61.69816, 
    61.9189, 62.13864, 62.35739, 62.57514, 62.7919, 63.00767, 63.22246, 
    63.43628, 63.64912, 63.861, 64.07191, 64.28186, 64.49085, 64.6989, 
    64.906, 65.11215, 65.31738, 65.52166, 65.72502, 65.92746, 66.12897, 
    66.32958, 66.52927,
  -45.90479, -45.77011, -45.63492, -45.49921, -45.36298, -45.22623, 
    -45.08895, -44.95113, -44.81279, -44.6739, -44.53447, -44.3945, 
    -44.25398, -44.1129, -43.97127, -43.82907, -43.68632, -43.543, -43.3991, 
    -43.25463, -43.10957, -42.96394, -42.81772, -42.67091, -42.52349, 
    -42.37549, -42.22688, -42.07766, -41.92784, -41.77739, -41.62633, 
    -41.47465, -41.32234, -41.1694, -41.01582, -40.8616, -40.70674, 
    -40.55123, -40.39507, -40.23825, -40.08077, -39.92263, -39.76382, 
    -39.60433, -39.44417, -39.28332, -39.12179, -38.95956, -38.79665, 
    -38.63303, -38.4687, -38.30367, -38.13793, -37.97147, -37.80428, 
    -37.63637, -37.46772, -37.29834, -37.12822, -36.95736, -36.78574, 
    -36.61337, -36.44025, -36.26635, -36.09169, -35.91626, -35.74005, 
    -35.56305, -35.38527, -35.2067, -35.02733, -34.84716, -34.66618, 
    -34.48439, -34.30179, -34.11836, -33.93411, -33.74903, -33.56312, 
    -33.37636, -33.18876, -33.00031, -32.81101, -32.62085, -32.42982, 
    -32.23793, -32.04516, -31.85152, -31.65699, -31.46157, -31.26526, 
    -31.06806, -30.86995, -30.67093, -30.471, -30.27016, -30.0684, -29.86571, 
    -29.66208, -29.45753, -29.25203, -29.04559, -28.8382, -28.62985, 
    -28.42055, -28.21029, -27.99905, -27.78684, -27.57366, -27.3595, 
    -27.14435, -26.92821, -26.71108, -26.49295, -26.27381, -26.05367, 
    -25.83252, -25.61035, -25.38716, -25.16295, -24.93771, -24.71144, 
    -24.48413, -24.25578, -24.02639, -23.79596, -23.56447, -23.33193, 
    -23.09833, -22.86367, -22.62794, -22.39115, -22.15328, -21.91434, 
    -21.67432, -21.43323, -21.19104, -20.94778, -20.70342, -20.45797, 
    -20.21143, -19.96378, -19.71504, -19.4652, -19.21425, -18.9622, 
    -18.70904, -18.45477, -18.19939, -17.9429, -17.68529, -17.42657, 
    -17.16672, -16.90576, -16.64368, -16.38049, -16.11617, -15.85072, 
    -15.58416, -15.31647, -15.04767, -14.77774, -14.50669, -14.23452, 
    -13.96122, -13.68681, -13.41127, -13.13462, -12.85685, -12.57797, 
    -12.29797, -12.01686, -11.73463, -11.4513, -11.16687, -10.88132, 
    -10.59468, -10.30694, -10.01811, -9.72818, -9.437164, -9.145064, 
    -8.851884, -8.557627, -8.262297, -7.9659, -7.66844, -7.369922, -7.070352, 
    -6.769734, -6.468076, -6.165381, -5.861658, -5.556911, -5.251147, 
    -4.944375, -4.6366, -4.327829, -4.018072, -3.707334, -3.395625, 
    -3.082953, -2.769325, -2.454752, -2.139242, -1.822804, -1.505448, 
    -1.187183, -0.8680198, -0.5479685, -0.2270396, 0.09475634, 0.4174082, 
    0.7409047, 1.065235, 1.390386, 1.716347, 2.043105, 2.370649, 2.698964, 
    3.02804, 3.357861, 3.688416, 4.01969, 4.351669, 4.68434, 5.017688, 
    5.3517, 5.686359, 6.021652, 6.357563, 6.694077, 7.031179, 7.368853, 
    7.707082, 8.045852, 8.385145, 8.724945, 9.065237, 9.406002, 9.747225, 
    10.08889, 10.43097, 10.77346, 11.11634, 11.45959, 11.80319, 12.14713, 
    12.49138, 12.83593, 13.18076, 13.52586, 13.87119, 14.21676, 14.56252, 
    14.90848, 15.25461, 15.60088, 15.94729, 16.29381, 16.64042, 16.98711, 
    17.33385, 17.68063, 18.02743, 18.37422, 18.721, 19.06774, 19.41441, 
    19.76101, 20.10752, 20.4539, 20.80016, 21.14626, 21.49218, 21.83792, 
    22.18345, 22.52875, 22.8738, 23.21859, 23.5631, 23.9073, 24.25118, 
    24.59473, 24.93792, 25.28074, 25.62317, 25.96519, 26.30678, 26.64793, 
    26.98862, 27.32884, 27.66856, 28.00777, 28.34646, 28.6846, 29.02218, 
    29.35919, 29.69561, 30.03143, 30.36662, 30.70118, 31.03509, 31.36833, 
    31.70089, 32.03276, 32.36392, 32.69436, 33.02406, 33.35302, 33.68121, 
    34.00864, 34.33527, 34.6611, 34.98612, 35.31032, 35.63369, 35.9562, 
    36.27786, 36.59866, 36.91856, 37.23759, 37.55571, 37.87292, 38.18921, 
    38.50457, 38.819, 39.13248, 39.445, 39.75655, 40.06713, 40.37674, 
    40.68535, 40.99297, 41.29958, 41.60518, 41.90977, 42.21333, 42.51586, 
    42.81736, 43.11781, 43.41721, 43.71556, 44.01286, 44.30909, 44.60424, 
    44.89833, 45.19134, 45.48327, 45.77411, 46.06387, 46.35253, 46.6401, 
    46.92657, 47.21193, 47.4962, 47.77935, 48.0614, 48.34233, 48.62216, 
    48.90087, 49.17846, 49.45493, 49.73029, 50.00453, 50.27764, 50.54964, 
    50.82051, 51.09026, 51.35889, 51.6264, 51.89279, 52.15805, 52.42219, 
    52.68521, 52.94712, 53.2079, 53.46757, 53.72611, 53.98355, 54.23986, 
    54.49507, 54.74916, 55.00215, 55.25402, 55.5048, 55.75446, 56.00303, 
    56.2505, 56.49687, 56.74215, 56.98633, 57.22943, 57.47144, 57.71236, 
    57.95221, 58.19098, 58.42868, 58.6653, 58.90086, 59.13535, 59.36878, 
    59.60116, 59.83248, 60.06275, 60.29197, 60.52015, 60.7473, 60.9734, 
    61.19848, 61.42253, 61.64556, 61.86757, 62.08856, 62.30854, 62.52752, 
    62.74549, 62.96247, 63.17845, 63.39344, 63.60745, 63.82048, 64.03253, 
    64.24361, 64.45372, 64.66287, 64.87106, 65.07831, 65.2846, 65.48994, 
    65.69435, 65.89783, 66.10037, 66.30199, 66.50269, 66.70248,
  -46.07022, -45.93574, -45.80074, -45.66522, -45.52918, -45.39262, 
    -45.25553, -45.1179, -44.97974, -44.84104, -44.7018, -44.562, -44.42167, 
    -44.28077, -44.13932, -43.9973, -43.85472, -43.71157, -43.56785, 
    -43.42355, -43.27867, -43.13321, -42.98715, -42.8405, -42.69326, 
    -42.54542, -42.39697, -42.24791, -42.09824, -41.94796, -41.79705, 
    -41.64552, -41.49336, -41.34056, -41.18713, -41.03306, -40.87834, 
    -40.72297, -40.56695, -40.41027, -40.25292, -40.09491, -39.93623, 
    -39.77687, -39.61683, -39.4561, -39.29469, -39.13258, -38.96978, 
    -38.80627, -38.64205, -38.47713, -38.31148, -38.14512, -37.97803, 
    -37.81021, -37.64165, -37.47236, -37.30233, -37.13154, -36.96, -36.7877, 
    -36.61465, -36.44082, -36.26622, -36.09084, -35.91469, -35.73774, 
    -35.56001, -35.38148, -35.20215, -35.02201, -34.84106, -34.6593, 
    -34.47672, -34.29331, -34.10907, -33.924, -33.73809, -33.55133, 
    -33.36372, -33.17526, -32.98594, -32.79576, -32.60471, -32.41278, 
    -32.21997, -32.02628, -31.83171, -31.63623, -31.43987, -31.24259, 
    -31.04441, -30.84532, -30.64531, -30.44437, -30.24251, -30.03971, 
    -29.83598, -29.63131, -29.42569, -29.21912, -29.01159, -28.8031, 
    -28.59365, -28.38322, -28.17182, -27.95944, -27.74608, -27.53173, 
    -27.31638, -27.10004, -26.8827, -26.66434, -26.44498, -26.2246, -26.0032, 
    -25.78078, -25.55733, -25.33285, -25.10733, -24.88077, -24.65316, 
    -24.42451, -24.1948, -23.96404, -23.73221, -23.49932, -23.26537, 
    -23.03034, -22.79424, -22.55706, -22.3188, -22.07945, -21.83902, 
    -21.59749, -21.35487, -21.11115, -20.86633, -20.62041, -20.37339, 
    -20.12525, -19.87601, -19.62564, -19.37417, -19.12158, -18.86786, 
    -18.61303, -18.35707, -18.09999, -17.84177, -17.58243, -17.32197, 
    -17.06037, -16.79763, -16.53377, -16.26877, -16.00263, -15.73537, 
    -15.46696, -15.19742, -14.92675, -14.65494, -14.38199, -14.10791, 
    -13.83269, -13.55634, -13.27886, -13.00025, -12.72051, -12.43964, 
    -12.15764, -11.87451, -11.59027, -11.3049, -11.01841, -10.73081, 
    -10.4421, -10.15227, -9.861341, -9.569306, -9.276172, -8.981942, 
    -8.686621, -8.390212, -8.09272, -7.794151, -7.494509, -7.193799, 
    -6.892026, -6.589197, -6.285317, -5.980393, -5.674431, -5.367437, 
    -5.059419, -4.750383, -4.440337, -4.129289, -3.817245, -3.504216, 
    -3.190208, -2.87523, -2.559292, -2.242402, -1.92457, -1.605805, 
    -1.286118, -0.9655175, -0.6440148, -0.3216203, 0.001655084, 0.3258002, 
    0.6508039, 0.9766544, 1.30334, 1.630848, 1.959167, 2.288284, 2.618186, 
    2.94886, 3.280293, 3.612472, 3.945381, 4.279009, 4.613339, 4.948359, 
    5.284052, 5.620406, 5.957403, 6.295029, 6.633269, 6.972106, 7.311525, 
    7.65151, 7.992044, 8.333111, 8.674694, 9.016777, 9.359342, 9.702372, 
    10.04585, 10.38976, 10.73408, 11.07879, 11.42389, 11.76934, 12.11513, 
    12.46124, 12.80766, 13.15437, 13.50134, 13.84855, 14.196, 14.54366, 
    14.89151, 15.23953, 15.5877, 15.93601, 16.28443, 16.63295, 16.98154, 
    17.33019, 17.67887, 18.02758, 18.37628, 18.72496, 19.07361, 19.42219, 
    19.77069, 20.1191, 20.46738, 20.81553, 21.16353, 21.51135, 21.85897, 
    22.20638, 22.55357, 22.9005, 23.24715, 23.59352, 23.93959, 24.28533, 
    24.63073, 24.97576, 25.32041, 25.66467, 26.00851, 26.35192, 26.69488, 
    27.03737, 27.37937, 27.72087, 28.06186, 28.40231, 28.7422, 29.08153, 
    29.42027, 29.75842, 30.09595, 30.43284, 30.76909, 31.10468, 31.43959, 
    31.77381, 32.10733, 32.44012, 32.77218, 33.1035, 33.43405, 33.76383, 
    34.09282, 34.42101, 34.74839, 35.07495, 35.40066, 35.72553, 36.04954, 
    36.37268, 36.69493, 37.01629, 37.33675, 37.65629, 37.97491, 38.29259, 
    38.60933, 38.92512, 39.23994, 39.5538, 39.86667, 40.17856, 40.48945, 
    40.79934, 41.10821, 41.41607, 41.7229, 42.0287, 42.33345, 42.63717, 
    42.93983, 43.24144, 43.54198, 43.84145, 44.13985, 44.43717, 44.73341, 
    45.02856, 45.32261, 45.61557, 45.90744, 46.19819, 46.48784, 46.77638, 
    47.0638, 47.35011, 47.6353, 47.91937, 48.20232, 48.48414, 48.76483, 
    49.0444, 49.32283, 49.60013, 49.8763, 50.15134, 50.42524, 50.69801, 
    50.96964, 51.24014, 51.50949, 51.77772, 52.04481, 52.31076, 52.57558, 
    52.83927, 53.10182, 53.36324, 53.62353, 53.88269, 54.14073, 54.39763, 
    54.65341, 54.90807, 55.16161, 55.41402, 55.66532, 55.9155, 56.16458, 
    56.41254, 56.65939, 56.90514, 57.14978, 57.39332, 57.63577, 57.87712, 
    58.11739, 58.35656, 58.59465, 58.83166, 59.06759, 59.30245, 59.53624, 
    59.76896, 60.00061, 60.2312, 60.46075, 60.68923, 60.91667, 61.14307, 
    61.36842, 61.59274, 61.81603, 62.03829, 62.25953, 62.47975, 62.69895, 
    62.91714, 63.13433, 63.35051, 63.5657, 63.7799, 63.9931, 64.20533, 
    64.41657, 64.62685, 64.83614, 65.04448, 65.25186, 65.45828, 65.66375, 
    65.86827, 66.07185, 66.27451, 66.47622, 66.677, 66.87687,
  -46.23638, -46.1021, -45.96729, -45.83197, -45.69613, -45.55976, -45.42286, 
    -45.28542, -45.14745, -45.00895, -44.86989, -44.73029, -44.59013, 
    -44.44942, -44.30815, -44.16632, -44.02392, -43.88095, -43.73741, 
    -43.59328, -43.44858, -43.30329, -43.15741, -43.01093, -42.86386, 
    -42.71618, -42.5679, -42.41901, -42.2695, -42.11938, -41.96863, 
    -41.81726, -41.66525, -41.51261, -41.35933, -41.20541, -41.05084, 
    -40.89561, -40.73973, -40.58319, -40.42599, -40.26811, -40.10956, 
    -39.95034, -39.79042, -39.62983, -39.46854, -39.30655, -39.14386, 
    -38.98047, -38.81637, -38.65155, -38.48602, -38.31976, -38.15277, 
    -37.98505, -37.81659, -37.64739, -37.47744, -37.30674, -37.13528, 
    -36.96306, -36.79008, -36.61632, -36.44179, -36.26648, -36.09038, 
    -35.91349, -35.73581, -35.55733, -35.37804, -35.19794, -35.01703, 
    -34.8353, -34.65274, -34.46936, -34.28514, -34.10008, -33.91418, 
    -33.72742, -33.53982, -33.35135, -33.16202, -32.97182, -32.78074, 
    -32.58879, -32.39595, -32.20222, -32.0076, -31.81208, -31.61566, 
    -31.41833, -31.22008, -31.02091, -30.82082, -30.6198, -30.41785, 
    -30.21496, -30.01112, -29.80634, -29.6006, -29.3939, -29.18624, 
    -28.97762, -28.76801, -28.55744, -28.34588, -28.13333, -27.91979, 
    -27.70526, -27.48972, -27.27318, -27.05562, -26.83706, -26.61747, 
    -26.39686, -26.17522, -25.95255, -25.72884, -25.50409, -25.27829, 
    -25.05145, -24.82355, -24.59459, -24.36457, -24.13349, -23.90133, 
    -23.6681, -23.43379, -23.19841, -22.96193, -22.72437, -22.48572, 
    -22.24597, -22.00512, -21.76317, -21.52011, -21.27595, -21.03067, 
    -20.78428, -20.53677, -20.28814, -20.03839, -19.78752, -19.53551, 
    -19.28238, -19.02812, -18.77272, -18.51618, -18.25851, -17.9997, 
    -17.73975, -17.47865, -17.21641, -16.95303, -16.6885, -16.42282, 
    -16.15599, -15.88802, -15.61889, -15.34862, -15.0772, -14.80463, 
    -14.53091, -14.25604, -13.98002, -13.70285, -13.42454, -13.14508, 
    -12.86448, -12.58273, -12.29984, -12.01582, -11.73065, -11.44435, 
    -11.15691, -10.86835, -10.57865, -10.28784, -9.995895, -9.702836, 
    -9.408663, -9.113378, -8.816986, -8.519492, -8.2209, -7.921214, -7.62044, 
    -7.318583, -7.015648, -6.711641, -6.406568, -6.100435, -5.793249, 
    -5.485015, -5.175742, -4.865436, -4.554104, -4.241755, -3.928396, 
    -3.614034, -3.29868, -2.982341, -2.665026, -2.346745, -2.027506, 
    -1.70732, -1.386197, -1.064146, -0.7411785, -0.4173047, -0.09253567, 
    0.2331173, 0.5596427, 0.8870288, 1.215264, 1.544335, 1.87423, 2.204937, 
    2.536442, 2.868732, 3.201794, 3.535613, 3.870177, 4.20547, 4.541478, 
    4.878187, 5.215582, 5.553648, 5.892368, 6.231729, 6.571714, 6.912307, 
    7.253492, 7.595252, 7.937572, 8.280434, 8.62382, 8.967715, 9.312101, 
    9.65696, 10.00228, 10.34803, 10.6942, 11.04078, 11.38774, 11.73506, 
    12.08273, 12.43073, 12.77904, 13.12764, 13.47651, 13.82563, 14.17498, 
    14.52455, 14.87432, 15.22426, 15.57435, 15.92458, 16.27493, 16.62538, 
    16.9759, 17.32648, 17.6771, 18.02773, 18.37837, 18.72898, 19.07955, 
    19.43006, 19.78049, 20.13083, 20.48104, 20.83111, 21.18102, 21.53076, 
    21.88029, 22.22961, 22.5787, 22.92752, 23.27608, 23.62434, 23.97229, 
    24.3199, 24.66717, 25.01407, 25.36058, 25.70669, 26.05238, 26.39762, 
    26.74241, 27.08672, 27.43053, 27.77384, 28.11661, 28.45885, 28.80052, 
    29.14161, 29.48211, 29.82199, 30.16125, 30.49987, 30.83783, 31.17512, 
    31.51172, 31.84762, 32.1828, 32.51724, 32.85094, 33.18388, 33.51605, 
    33.84743, 34.17801, 34.50777, 34.83671, 35.16481, 35.49207, 35.81845, 
    36.14397, 36.4686, 36.79233, 37.11515, 37.43705, 37.75803, 38.07807, 
    38.39716, 38.71529, 39.03244, 39.34863, 39.66383, 39.97803, 40.29123, 
    40.60342, 40.91459, 41.22473, 41.53384, 41.84191, 42.14893, 42.4549, 
    42.7598, 43.06364, 43.36641, 43.66809, 43.96869, 44.2682, 44.56662, 
    44.86395, 45.16016, 45.45527, 45.74927, 46.04215, 46.33391, 46.62455, 
    46.91407, 47.20246, 47.48971, 47.77583, 48.06082, 48.34467, 48.62738, 
    48.90894, 49.18936, 49.46864, 49.74677, 50.02375, 50.29959, 50.57428, 
    50.84782, 51.12021, 51.39145, 51.66154, 51.93048, 52.19828, 52.46492, 
    52.73042, 52.99477, 53.25797, 53.52003, 53.78094, 54.04071, 54.29935, 
    54.55684, 54.81319, 55.06841, 55.3225, 55.57545, 55.82728, 56.07797, 
    56.32755, 56.576, 56.82333, 57.06954, 57.31464, 57.55863, 57.80151, 
    58.04329, 58.28396, 58.52354, 58.76202, 58.99941, 59.23571, 59.47093, 
    59.70507, 59.93813, 60.17011, 60.40103, 60.63088, 60.85967, 61.0874, 
    61.31408, 61.53971, 61.7643, 61.98784, 62.21035, 62.43182, 62.65227, 
    62.8717, 63.0901, 63.3075, 63.52388, 63.73926, 63.95364, 64.16702, 
    64.37941, 64.59081, 64.80124, 65.01068, 65.21915, 65.42666, 65.63321, 
    65.83879, 66.04343, 66.24712, 66.44986, 66.65166, 66.85253, 67.05247,
  -46.40327, -46.26919, -46.13459, -45.99947, -45.86382, -45.72765, 
    -45.59095, -45.45371, -45.31593, -45.17762, -45.03876, -44.89935, 
    -44.75938, -44.61886, -44.47778, -44.33614, -44.19392, -44.05114, 
    -43.90778, -43.76384, -43.61931, -43.4742, -43.3285, -43.1822, -43.0353, 
    -42.88779, -42.73969, -42.59096, -42.44162, -42.29166, -42.14108, 
    -41.98987, -41.83803, -41.68554, -41.53242, -41.37865, -41.22424, 
    -41.06916, -40.91343, -40.75703, -40.59997, -40.44224, -40.28383, 
    -40.12474, -39.96496, -39.8045, -39.64334, -39.48148, -39.31891, 
    -39.15564, -38.99166, -38.82696, -38.66153, -38.49538, -38.3285, 
    -38.16088, -37.99253, -37.82343, -37.65357, -37.48296, -37.31159, 
    -37.13946, -36.96655, -36.79287, -36.61842, -36.44317, -36.26714, 
    -36.09032, -35.91269, -35.73426, -35.55503, -35.37497, -35.1941, 
    -35.01241, -34.82989, -34.64653, -34.46233, -34.27729, -34.0914, 
    -33.90466, -33.71706, -33.52859, -33.33925, -33.14904, -32.95795, 
    -32.76598, -32.57311, -32.37935, -32.1847, -31.98913, -31.79266, 
    -31.59527, -31.39696, -31.19773, -30.99756, -30.79646, -30.59443, 
    -30.39144, -30.18751, -29.98262, -29.77677, -29.56995, -29.36217, 
    -29.1534, -28.94366, -28.73294, -28.52122, -28.30851, -28.0948, 
    -27.88009, -27.66437, -27.44763, -27.22988, -27.0111, -26.79129, 
    -26.57046, -26.34858, -26.12567, -25.9017, -25.67669, -25.45063, 
    -25.2235, -24.99531, -24.76605, -24.53573, -24.30432, -24.07184, 
    -23.83827, -23.60362, -23.36787, -23.13103, -22.89309, -22.65405, 
    -22.4139, -22.17264, -21.93027, -21.68678, -21.44217, -21.19644, 
    -20.94958, -20.7016, -20.45248, -20.20223, -19.95084, -19.69831, 
    -19.44464, -19.18983, -18.93387, -18.67676, -18.4185, -18.15909, 
    -17.89852, -17.6368, -17.37392, -17.10988, -16.84469, -16.57833, 
    -16.31081, -16.04213, -15.77229, -15.50128, -15.22911, -14.95578, 
    -14.68128, -14.40562, -14.1288, -13.85082, -13.57167, -13.29137, 
    -13.0099, -12.72728, -12.4435, -12.15856, -11.87247, -11.58523, 
    -11.29685, -11.00731, -10.71664, -10.42482, -10.13186, -9.837777, 
    -9.542558, -9.246213, -8.948746, -8.65016, -8.35046, -8.049651, 
    -7.747739, -7.444727, -7.140623, -6.83543, -6.529155, -6.221805, 
    -5.913386, -5.603904, -5.293366, -4.98178, -4.669153, -4.355492, 
    -4.040806, -3.725103, -3.408391, -3.090678, -2.771975, -2.45229, 
    -2.131633, -1.810013, -1.48744, -1.163926, -0.8394794, -0.5141123, 
    -0.1878354, 0.13934, 0.4674021, 0.7963391, 1.126139, 1.456789, 1.788277, 
    2.12059, 2.453715, 2.787637, 3.122345, 3.457823, 3.794058, 4.131035, 
    4.46874, 4.807158, 5.146272, 5.48607, 5.826534, 6.167649, 6.509399, 
    6.851768, 7.194739, 7.538296, 7.882421, 8.227098, 8.572311, 8.91804, 
    9.26427, 9.61098, 9.958156, 10.30578, 10.65382, 11.00228, 11.35113, 
    11.70035, 12.04992, 12.39983, 12.75005, 13.10057, 13.45136, 13.80241, 
    14.1537, 14.50521, 14.85691, 15.20879, 15.56083, 15.91301, 16.26531, 
    16.61771, 16.97019, 17.32272, 17.67529, 18.02789, 18.38048, 18.73305, 
    19.08557, 19.43804, 19.79042, 20.1427, 20.49486, 20.84688, 21.19873, 
    21.55041, 21.90188, 22.25313, 22.60415, 22.9549, 23.30537, 23.65554, 
    24.0054, 24.35492, 24.70408, 25.05287, 25.40126, 25.74924, 26.09679, 
    26.4439, 26.79053, 27.13668, 27.48233, 27.82746, 28.17205, 28.51609, 
    28.85955, 29.20243, 29.5447, 29.88635, 30.22737, 30.56773, 30.90742, 
    31.24642, 31.58473, 31.92232, 32.25918, 32.59529, 32.93065, 33.26524, 
    33.59903, 33.93203, 34.26421, 34.59557, 34.92609, 35.25575, 35.58455, 
    35.91247, 36.23951, 36.56564, 36.89086, 37.21516, 37.53853, 37.86095, 
    38.18242, 38.50292, 38.82245, 39.141, 39.45856, 39.77511, 40.09065, 
    40.40518, 40.71867, 41.03114, 41.34256, 41.65293, 41.96224, 42.27049, 
    42.57767, 42.88378, 43.1888, 43.49273, 43.79557, 44.09731, 44.39794, 
    44.69746, 44.99587, 45.29316, 45.58933, 45.88437, 46.17828, 46.47105, 
    46.76269, 47.05319, 47.34254, 47.63075, 47.9178, 48.20371, 48.48846, 
    48.77206, 49.0545, 49.33578, 49.61591, 49.89487, 50.17267, 50.44931, 
    50.72478, 50.9991, 51.27224, 51.54423, 51.81505, 52.08471, 52.35321, 
    52.62054, 52.88671, 53.15173, 53.41558, 53.67828, 53.93982, 54.2002, 
    54.45943, 54.7175, 54.97443, 55.23021, 55.48484, 55.73833, 55.99068, 
    56.24189, 56.49196, 56.7409, 56.9887, 57.23538, 57.48093, 57.72536, 
    57.96868, 58.21087, 58.45196, 58.69193, 58.9308, 59.16857, 59.40524, 
    59.64081, 59.87529, 60.10869, 60.341, 60.57223, 60.80239, 61.03148, 
    61.2595, 61.48645, 61.71236, 61.9372, 62.161, 62.38375, 62.60546, 
    62.82613, 63.04578, 63.26439, 63.48198, 63.69856, 63.91412, 64.12868, 
    64.34222, 64.55478, 64.76633, 64.97691, 65.18649, 65.3951, 65.60273, 
    65.80939, 66.01509, 66.21983, 66.42361, 66.62645, 66.82834, 67.02929, 
    67.2293 ;

 lat =
  21.14534, 21.18575, 21.22604, 21.2662, 21.30622, 21.34612, 21.38589, 
    21.42553, 21.46503, 21.50441, 21.54366, 21.58277, 21.62175, 21.6606, 
    21.69932, 21.73791, 21.77636, 21.81468, 21.85287, 21.89092, 21.92884, 
    21.96663, 22.00429, 22.04181, 22.07919, 22.11644, 22.15356, 22.19054, 
    22.22739, 22.2641, 22.30067, 22.33711, 22.37342, 22.40958, 22.44561, 
    22.48151, 22.51726, 22.55288, 22.58836, 22.62371, 22.65891, 22.69398, 
    22.72891, 22.7637, 22.79836, 22.83287, 22.86724, 22.90148, 22.93557, 
    22.96953, 23.00334, 23.03702, 23.07055, 23.10394, 23.1372, 23.17031, 
    23.20328, 23.2361, 23.26879, 23.30133, 23.33374, 23.366, 23.39811, 
    23.43009, 23.46192, 23.4936, 23.52515, 23.55655, 23.5878, 23.61891, 
    23.64988, 23.6807, 23.71138, 23.74191, 23.7723, 23.80255, 23.83264, 
    23.86259, 23.8924, 23.92206, 23.95157, 23.98093, 24.01015, 24.03922, 
    24.06815, 24.09693, 24.12556, 24.15404, 24.18237, 24.21055, 24.23859, 
    24.26648, 24.29422, 24.32181, 24.34925, 24.37654, 24.40368, 24.43068, 
    24.45752, 24.48421, 24.51076, 24.53715, 24.56339, 24.58948, 24.61542, 
    24.6412, 24.66684, 24.69232, 24.71766, 24.74284, 24.76787, 24.79274, 
    24.81747, 24.84204, 24.86646, 24.89072, 24.91483, 24.93879, 24.96259, 
    24.98625, 25.00974, 25.03309, 25.05627, 25.07931, 25.10219, 25.12491, 
    25.14748, 25.1699, 25.19216, 25.21426, 25.23621, 25.258, 25.27964, 
    25.30112, 25.32245, 25.34361, 25.36463, 25.38548, 25.40618, 25.42672, 
    25.4471, 25.46733, 25.4874, 25.50731, 25.52706, 25.54666, 25.5661, 
    25.58538, 25.6045, 25.62346, 25.64226, 25.66091, 25.6794, 25.69772, 
    25.71589, 25.7339, 25.75175, 25.76944, 25.78697, 25.80434, 25.82154, 
    25.83859, 25.85548, 25.87221, 25.88878, 25.90519, 25.92143, 25.93752, 
    25.95345, 25.96921, 25.98481, 26.00025, 26.01553, 26.03065, 26.0456, 
    26.0604, 26.07503, 26.0895, 26.10381, 26.11795, 26.13194, 26.14576, 
    26.15941, 26.17291, 26.18624, 26.19941, 26.21242, 26.22526, 26.23794, 
    26.25045, 26.26281, 26.275, 26.28702, 26.29888, 26.31058, 26.32211, 
    26.33348, 26.34469, 26.35573, 26.36661, 26.37732, 26.38787, 26.39825, 
    26.40847, 26.41852, 26.42841, 26.43814, 26.4477, 26.45709, 26.46632, 
    26.47539, 26.48428, 26.49302, 26.50159, 26.50999, 26.51822, 26.5263, 
    26.5342, 26.54194, 26.54951, 26.55692, 26.56417, 26.57124, 26.57815, 
    26.5849, 26.59147, 26.59789, 26.60413, 26.61021, 26.61613, 26.62187, 
    26.62745, 26.63287, 26.63811, 26.64319, 26.64811, 26.65285, 26.65743, 
    26.66185, 26.6661, 26.67018, 26.67409, 26.67784, 26.68142, 26.68483, 
    26.68808, 26.69115, 26.69407, 26.69681, 26.69939, 26.7018, 26.70404, 
    26.70612, 26.70803, 26.70977, 26.71135, 26.71276, 26.71399, 26.71507, 
    26.71597, 26.71671, 26.71729, 26.71769, 26.71793, 26.718, 26.7179, 
    26.71764, 26.71721, 26.71661, 26.71584, 26.71491, 26.71381, 26.71254, 
    26.71111, 26.70951, 26.70774, 26.7058, 26.7037, 26.70143, 26.69899, 
    26.69639, 26.69362, 26.69068, 26.68757, 26.6843, 26.68086, 26.67726, 
    26.67348, 26.66954, 26.66544, 26.66116, 26.65672, 26.65211, 26.64734, 
    26.6424, 26.63729, 26.63202, 26.62658, 26.62097, 26.6152, 26.60926, 
    26.60316, 26.59688, 26.59045, 26.58384, 26.57707, 26.57014, 26.56303, 
    26.55576, 26.54833, 26.54073, 26.53296, 26.52503, 26.51693, 26.50867, 
    26.50024, 26.49165, 26.48289, 26.47396, 26.46487, 26.45562, 26.4462, 
    26.43661, 26.42686, 26.41694, 26.40686, 26.39662, 26.38621, 26.37564, 
    26.3649, 26.35399, 26.34293, 26.3317, 26.3203, 26.30874, 26.29702, 
    26.28513, 26.27308, 26.26086, 26.24849, 26.23594, 26.22324, 26.21037, 
    26.19734, 26.18414, 26.17079, 26.15726, 26.14358, 26.12974, 26.11573, 
    26.10156, 26.08722, 26.07273, 26.05807, 26.04325, 26.02827, 26.01313, 
    25.99782, 25.98236, 25.96673, 25.95094, 25.93499, 25.91888, 25.9026, 
    25.88617, 25.86958, 25.85282, 25.83591, 25.81883, 25.8016, 25.7842, 
    25.76665, 25.74893, 25.73106, 25.71303, 25.69483, 25.67648, 25.65797, 
    25.6393, 25.62047, 25.60148, 25.58234, 25.56303, 25.54357, 25.52395, 
    25.50417, 25.48424, 25.46414, 25.44389, 25.42348, 25.40291, 25.38219, 
    25.36131, 25.34028, 25.31908, 25.29773, 25.27623, 25.25457, 25.23275, 
    25.21078, 25.18865, 25.16636, 25.14392, 25.12133, 25.09858, 25.07568, 
    25.05262, 25.0294, 25.00604, 24.98252, 24.95884, 24.93501, 24.91103, 
    24.88689, 24.8626, 24.83816, 24.81357, 24.78882, 24.76392, 24.73886, 
    24.71366, 24.6883, 24.66279, 24.63713, 24.61132, 24.58536, 24.55925, 
    24.53298, 24.50657, 24.48, 24.45328, 24.42642, 24.3994, 24.37224, 
    24.34492, 24.31746,
  21.246, 21.28648, 21.32683, 21.36705, 21.40714, 21.4471, 21.48693, 
    21.52663, 21.5662, 21.60563, 21.64494, 21.68411, 21.72316, 21.76207, 
    21.80085, 21.83949, 21.87801, 21.91639, 21.95464, 21.99275, 22.03073, 
    22.06858, 22.10629, 22.14387, 22.18132, 22.21863, 22.2558, 22.29284, 
    22.32975, 22.36652, 22.40315, 22.43965, 22.47601, 22.51223, 22.54832, 
    22.58427, 22.62008, 22.65576, 22.6913, 22.7267, 22.76196, 22.79709, 
    22.83207, 22.86692, 22.90163, 22.9362, 22.97063, 23.00492, 23.03907, 
    23.07308, 23.10695, 23.14067, 23.17426, 23.20771, 23.24102, 23.27418, 
    23.30721, 23.34009, 23.37283, 23.40542, 23.43788, 23.47019, 23.50236, 
    23.53439, 23.56627, 23.59801, 23.62961, 23.66106, 23.69236, 23.72353, 
    23.75455, 23.78542, 23.81615, 23.84673, 23.87717, 23.90746, 23.93761, 
    23.96761, 23.99747, 24.02717, 24.05674, 24.08615, 24.11542, 24.14454, 
    24.17351, 24.20234, 24.23101, 24.25954, 24.28792, 24.31616, 24.34424, 
    24.37218, 24.39996, 24.4276, 24.45509, 24.48243, 24.50961, 24.53665, 
    24.56354, 24.59028, 24.61687, 24.6433, 24.66959, 24.69572, 24.7217, 
    24.74754, 24.77322, 24.79874, 24.82412, 24.84934, 24.87442, 24.89934, 
    24.9241, 24.94872, 24.97318, 24.99748, 25.02164, 25.04564, 25.06948, 
    25.09317, 25.11671, 25.14009, 25.16332, 25.1864, 25.20932, 25.23208, 
    25.25469, 25.27714, 25.29944, 25.32158, 25.34357, 25.3654, 25.38708, 
    25.40859, 25.42996, 25.45116, 25.47221, 25.4931, 25.51383, 25.53441, 
    25.55483, 25.57509, 25.5952, 25.61514, 25.63493, 25.65456, 25.67403, 
    25.69335, 25.7125, 25.7315, 25.75033, 25.76901, 25.78753, 25.80589, 
    25.82409, 25.84213, 25.86001, 25.87773, 25.89529, 25.91269, 25.92993, 
    25.94701, 25.96393, 25.98069, 25.99729, 26.01373, 26.03, 26.04611, 
    26.06207, 26.07786, 26.09349, 26.10896, 26.12426, 26.13941, 26.15439, 
    26.16921, 26.18387, 26.19837, 26.2127, 26.22687, 26.24088, 26.25472, 
    26.26841, 26.28192, 26.29528, 26.30847, 26.3215, 26.33437, 26.34707, 
    26.35961, 26.37198, 26.38419, 26.39624, 26.40812, 26.41984, 26.4314, 
    26.44279, 26.45401, 26.46507, 26.47597, 26.4867, 26.49727, 26.50767, 
    26.51791, 26.52798, 26.53789, 26.54763, 26.55721, 26.56662, 26.57586, 
    26.58494, 26.59386, 26.60261, 26.61119, 26.61961, 26.62786, 26.63595, 
    26.64387, 26.65162, 26.65921, 26.66663, 26.67389, 26.68097, 26.6879, 
    26.69465, 26.70124, 26.70767, 26.71393, 26.72002, 26.72594, 26.7317, 
    26.73729, 26.74271, 26.74797, 26.75306, 26.75798, 26.76274, 26.76732, 
    26.77175, 26.776, 26.78009, 26.78401, 26.78776, 26.79135, 26.79477, 
    26.79802, 26.80111, 26.80402, 26.80677, 26.80935, 26.81177, 26.81402, 
    26.8161, 26.81801, 26.81976, 26.82133, 26.82274, 26.82399, 26.82506, 
    26.82597, 26.82671, 26.82729, 26.82769, 26.82793, 26.828, 26.8279, 
    26.82764, 26.82721, 26.82661, 26.82584, 26.82491, 26.8238, 26.82253, 
    26.8211, 26.81949, 26.81772, 26.81578, 26.81367, 26.8114, 26.80896, 
    26.80635, 26.80357, 26.80063, 26.79752, 26.79424, 26.79079, 26.78718, 
    26.7834, 26.77945, 26.77534, 26.77106, 26.76661, 26.762, 26.75721, 
    26.75226, 26.74715, 26.74186, 26.73641, 26.7308, 26.72501, 26.71906, 
    26.71295, 26.70666, 26.70021, 26.6936, 26.68682, 26.67986, 26.67275, 
    26.66547, 26.65802, 26.65041, 26.64263, 26.63468, 26.62657, 26.61829, 
    26.60984, 26.60123, 26.59246, 26.58352, 26.57441, 26.56514, 26.5557, 
    26.5461, 26.53633, 26.5264, 26.5163, 26.50604, 26.49561, 26.48502, 
    26.47426, 26.46334, 26.45225, 26.441, 26.42958, 26.418, 26.40626, 
    26.39435, 26.38227, 26.37004, 26.35764, 26.34507, 26.33234, 26.31945, 
    26.3064, 26.29318, 26.2798, 26.26625, 26.25254, 26.23867, 26.22464, 
    26.21044, 26.19608, 26.18156, 26.16688, 26.15203, 26.13702, 26.12185, 
    26.10652, 26.09103, 26.07537, 26.05956, 26.04358, 26.02744, 26.01114, 
    25.99467, 25.97805, 25.96127, 25.94432, 25.92722, 25.90995, 25.89252, 
    25.87494, 25.85719, 25.83929, 25.82122, 25.803, 25.78461, 25.76607, 
    25.74737, 25.7285, 25.70948, 25.6903, 25.67097, 25.65147, 25.63181, 
    25.612, 25.59203, 25.5719, 25.55161, 25.53117, 25.51056, 25.48981, 
    25.46889, 25.44782, 25.42659, 25.4052, 25.38366, 25.36196, 25.3401, 
    25.31809, 25.29593, 25.2736, 25.25112, 25.22849, 25.2057, 25.18276, 
    25.15966, 25.1364, 25.113, 25.08944, 25.06572, 25.04185, 25.01782, 
    24.99365, 24.96932, 24.94483, 24.92019, 24.8954, 24.87046, 24.84537, 
    24.82012, 24.79472, 24.76917, 24.74346, 24.71761, 24.6916, 24.66544, 
    24.63913, 24.61267, 24.58606, 24.5593, 24.53238, 24.50532, 24.47811, 
    24.45075, 24.42324,
  21.34666, 21.3872, 21.42761, 21.46789, 21.50804, 21.54807, 21.58796, 
    21.62772, 21.66735, 21.70684, 21.74621, 21.78545, 21.82455, 21.86352, 
    21.90236, 21.94107, 21.97964, 22.01808, 22.05639, 22.09456, 22.13261, 
    22.17051, 22.20829, 22.24592, 22.28343, 22.3208, 22.35803, 22.39513, 
    22.43209, 22.46892, 22.50561, 22.54217, 22.57859, 22.61487, 22.65101, 
    22.68702, 22.72289, 22.75863, 22.79422, 22.82968, 22.865, 22.90018, 
    22.93522, 22.97013, 23.00489, 23.03951, 23.074, 23.10835, 23.14255, 
    23.17661, 23.21054, 23.24432, 23.27797, 23.31147, 23.34483, 23.37805, 
    23.41113, 23.44406, 23.47685, 23.50951, 23.54201, 23.57438, 23.6066, 
    23.63868, 23.67062, 23.70241, 23.73405, 23.76556, 23.79692, 23.82813, 
    23.8592, 23.89013, 23.92091, 23.95154, 23.98203, 24.01237, 24.04257, 
    24.07262, 24.10253, 24.13228, 24.16189, 24.19136, 24.22067, 24.24984, 
    24.27887, 24.30774, 24.33647, 24.36504, 24.39347, 24.42175, 24.44988, 
    24.47787, 24.5057, 24.53338, 24.56092, 24.5883, 24.61554, 24.64262, 
    24.66955, 24.69634, 24.72297, 24.74945, 24.77578, 24.80196, 24.82799, 
    24.85386, 24.87959, 24.90516, 24.93058, 24.95585, 24.98096, 25.00592, 
    25.03073, 25.05539, 25.07989, 25.10424, 25.12843, 25.15247, 25.17636, 
    25.20009, 25.22367, 25.2471, 25.27036, 25.29348, 25.31644, 25.33924, 
    25.36189, 25.38438, 25.40672, 25.4289, 25.45093, 25.47279, 25.49451, 
    25.51606, 25.53746, 25.5587, 25.57979, 25.60072, 25.62149, 25.6421, 
    25.66256, 25.68285, 25.70299, 25.72297, 25.7428, 25.76246, 25.78197, 
    25.80131, 25.8205, 25.83953, 25.8584, 25.87711, 25.89566, 25.91406, 
    25.93229, 25.95036, 25.96827, 25.98602, 26.00362, 26.02105, 26.03832, 
    26.05543, 26.07238, 26.08916, 26.10579, 26.12226, 26.13856, 26.15471, 
    26.17069, 26.18651, 26.20217, 26.21766, 26.23299, 26.24817, 26.26318, 
    26.27802, 26.29271, 26.30723, 26.32159, 26.33578, 26.34982, 26.36369, 
    26.37739, 26.39094, 26.40432, 26.41753, 26.43059, 26.44347, 26.4562, 
    26.46876, 26.48116, 26.49339, 26.50546, 26.51736, 26.5291, 26.54068, 
    26.55209, 26.56333, 26.57442, 26.58533, 26.59608, 26.60667, 26.61709, 
    26.62735, 26.63744, 26.64736, 26.65712, 26.66671, 26.67614, 26.68541, 
    26.6945, 26.70343, 26.7122, 26.7208, 26.72923, 26.7375, 26.7456, 
    26.75353, 26.7613, 26.7689, 26.77634, 26.78361, 26.79071, 26.79764, 
    26.80441, 26.81101, 26.81745, 26.82372, 26.82982, 26.83575, 26.84152, 
    26.84712, 26.85255, 26.85782, 26.86292, 26.86785, 26.87262, 26.87721, 
    26.88165, 26.88591, 26.89, 26.89393, 26.89769, 26.90128, 26.90471, 
    26.90797, 26.91106, 26.91398, 26.91673, 26.91932, 26.92174, 26.92399, 
    26.92608, 26.92799, 26.92974, 26.93132, 26.93274, 26.93398, 26.93506, 
    26.93597, 26.93671, 26.93728, 26.93769, 26.93793, 26.938, 26.9379, 
    26.93764, 26.9372, 26.9366, 26.93583, 26.9349, 26.93379, 26.93252, 
    26.93108, 26.92948, 26.9277, 26.92576, 26.92365, 26.92137, 26.91892, 
    26.91631, 26.91353, 26.91058, 26.90746, 26.90418, 26.90073, 26.89711, 
    26.89332, 26.88937, 26.88524, 26.88095, 26.8765, 26.87187, 26.86708, 
    26.86213, 26.857, 26.85171, 26.84625, 26.84062, 26.83483, 26.82887, 
    26.82274, 26.81644, 26.80998, 26.80335, 26.79656, 26.78959, 26.78247, 
    26.77517, 26.76771, 26.76008, 26.75229, 26.74433, 26.7362, 26.72791, 
    26.71945, 26.71082, 26.70203, 26.69308, 26.68395, 26.67466, 26.66521, 
    26.65559, 26.6458, 26.63585, 26.62573, 26.61545, 26.60501, 26.59439, 
    26.58362, 26.57267, 26.56157, 26.55029, 26.53886, 26.52726, 26.51549, 
    26.50356, 26.49147, 26.47921, 26.46678, 26.4542, 26.44145, 26.42853, 
    26.41545, 26.40221, 26.38881, 26.37524, 26.3615, 26.34761, 26.33355, 
    26.31933, 26.30494, 26.2904, 26.27568, 26.26081, 26.24578, 26.23058, 
    26.21522, 26.1997, 26.18402, 26.16817, 26.15216, 26.13599, 26.11967, 
    26.10317, 26.08652, 26.06971, 26.05273, 26.0356, 26.0183, 26.00084, 
    25.98323, 25.96545, 25.94751, 25.92941, 25.91116, 25.89274, 25.87416, 
    25.85543, 25.83653, 25.81748, 25.79826, 25.77889, 25.75936, 25.73967, 
    25.71982, 25.69982, 25.67965, 25.65933, 25.63885, 25.61821, 25.59742, 
    25.57646, 25.55535, 25.53409, 25.51266, 25.49108, 25.46935, 25.44745, 
    25.4254, 25.4032, 25.38083, 25.35832, 25.33564, 25.31282, 25.28983, 
    25.26669, 25.2434, 25.21995, 25.19635, 25.17259, 25.14868, 25.12461, 
    25.1004, 25.07602, 25.0515, 25.02682, 25.00198, 24.977, 24.95186, 
    24.92657, 24.90112, 24.87553, 24.84978, 24.82388, 24.79783, 24.77163, 
    24.74527, 24.71877, 24.69211, 24.6653, 24.63835, 24.61124, 24.58398, 
    24.55657, 24.52901,
  21.4473, 21.4879, 21.52838, 21.56872, 21.60893, 21.64902, 21.68897, 
    21.72879, 21.76848, 21.80804, 21.84747, 21.88677, 21.92593, 21.96496, 
    22.00386, 22.04263, 22.08126, 22.11977, 22.15813, 22.19637, 22.23447, 
    22.27243, 22.31027, 22.34797, 22.38553, 22.42296, 22.46025, 22.49741, 
    22.53443, 22.57131, 22.60806, 22.64468, 22.68115, 22.71749, 22.7537, 
    22.78976, 22.82569, 22.86148, 22.89713, 22.93265, 22.96803, 23.00326, 
    23.03836, 23.07332, 23.10814, 23.14282, 23.17736, 23.21176, 23.24602, 
    23.28014, 23.31412, 23.34796, 23.38166, 23.41522, 23.44863, 23.4819, 
    23.51504, 23.54803, 23.58087, 23.61358, 23.64614, 23.67856, 23.71083, 
    23.74296, 23.77495, 23.8068, 23.8385, 23.87005, 23.90146, 23.93273, 
    23.96385, 23.99483, 24.02566, 24.05634, 24.08688, 24.11728, 24.14752, 
    24.17762, 24.20758, 24.23738, 24.26705, 24.29656, 24.32592, 24.35514, 
    24.38421, 24.41314, 24.44191, 24.47054, 24.49901, 24.52734, 24.55552, 
    24.58355, 24.61143, 24.63916, 24.66674, 24.69417, 24.72145, 24.74858, 
    24.77556, 24.80239, 24.82907, 24.85559, 24.88197, 24.90819, 24.93427, 
    24.96018, 24.98595, 25.01157, 25.03703, 25.06234, 25.0875, 25.1125, 
    25.13735, 25.16205, 25.1866, 25.21099, 25.23522, 25.25931, 25.28323, 
    25.30701, 25.33063, 25.35409, 25.3774, 25.40055, 25.42355, 25.4464, 
    25.46908, 25.49162, 25.51399, 25.53621, 25.55828, 25.58018, 25.60193, 
    25.62353, 25.64496, 25.66624, 25.68736, 25.70833, 25.72913, 25.74978, 
    25.77028, 25.79061, 25.81078, 25.8308, 25.85066, 25.87036, 25.8899, 
    25.90928, 25.9285, 25.94756, 25.96646, 25.98521, 26.00379, 26.02222, 
    26.04048, 26.05859, 26.07653, 26.09431, 26.11194, 26.1294, 26.1467, 
    26.16384, 26.18082, 26.19764, 26.21429, 26.23079, 26.24712, 26.26329, 
    26.2793, 26.29515, 26.31084, 26.32636, 26.34172, 26.35692, 26.37196, 
    26.38683, 26.40154, 26.41609, 26.43047, 26.44469, 26.45875, 26.47265, 
    26.48638, 26.49995, 26.51335, 26.52659, 26.53967, 26.55258, 26.56533, 
    26.57791, 26.59033, 26.60258, 26.61468, 26.6266, 26.63836, 26.64996, 
    26.66139, 26.67266, 26.68376, 26.69469, 26.70546, 26.71607, 26.72651, 
    26.73678, 26.74689, 26.75683, 26.76661, 26.77622, 26.78567, 26.79495, 
    26.80406, 26.81301, 26.82179, 26.8304, 26.83885, 26.84713, 26.85525, 
    26.8632, 26.87098, 26.87859, 26.88604, 26.89332, 26.90044, 26.90739, 
    26.91417, 26.92078, 26.92723, 26.93351, 26.93962, 26.94557, 26.95135, 
    26.95696, 26.9624, 26.96768, 26.97278, 26.97772, 26.9825, 26.9871, 
    26.99154, 26.99581, 26.99991, 27.00385, 27.00762, 27.01122, 27.01465, 
    27.01791, 27.02101, 27.02394, 27.0267, 27.02929, 27.03171, 27.03397, 
    27.03605, 27.03798, 27.03973, 27.04131, 27.04273, 27.04397, 27.04505, 
    27.04597, 27.04671, 27.04728, 27.04769, 27.04793, 27.048, 27.0479, 
    27.04764, 27.0472, 27.0466, 27.04583, 27.04489, 27.04379, 27.04251, 
    27.04107, 27.03946, 27.03768, 27.03574, 27.03362, 27.03134, 27.02889, 
    27.02627, 27.02348, 27.02053, 27.01741, 27.01412, 27.01066, 27.00703, 
    27.00324, 26.99928, 26.99515, 26.99085, 26.98639, 26.98175, 26.97695, 
    26.97199, 26.96685, 26.96155, 26.95608, 26.95044, 26.94464, 26.93867, 
    26.93253, 26.92622, 26.91975, 26.91311, 26.9063, 26.89933, 26.89218, 
    26.88488, 26.8774, 26.86976, 26.86195, 26.85398, 26.84583, 26.83753, 
    26.82905, 26.82041, 26.8116, 26.80263, 26.79349, 26.78418, 26.77471, 
    26.76508, 26.75527, 26.7453, 26.73517, 26.72487, 26.7144, 26.70377, 
    26.69297, 26.68201, 26.67088, 26.65959, 26.64813, 26.63651, 26.62473, 
    26.61277, 26.60066, 26.58838, 26.57593, 26.56332, 26.55055, 26.53761, 
    26.52451, 26.51124, 26.49781, 26.48422, 26.47046, 26.45654, 26.44246, 
    26.42821, 26.4138, 26.39923, 26.38449, 26.36959, 26.35453, 26.3393, 
    26.32392, 26.30837, 26.29266, 26.27678, 26.26075, 26.24455, 26.22819, 
    26.21167, 26.19499, 26.17814, 26.16114, 26.14397, 26.12665, 26.10916, 
    26.09151, 26.0737, 26.05573, 26.0376, 26.01931, 26.00086, 25.98226, 
    25.96349, 25.94456, 25.92547, 25.90622, 25.88682, 25.86725, 25.84753, 
    25.82764, 25.8076, 25.7874, 25.76704, 25.74653, 25.72585, 25.70502, 
    25.68403, 25.66289, 25.64158, 25.62012, 25.5985, 25.57673, 25.5548, 
    25.53271, 25.51046, 25.48806, 25.46551, 25.44279, 25.41993, 25.3969, 
    25.37372, 25.35039, 25.3269, 25.30326, 25.27946, 25.25551, 25.2314, 
    25.20714, 25.18272, 25.15816, 25.13343, 25.10856, 25.08353, 25.05835, 
    25.03301, 25.00753, 24.98189, 24.95609, 24.93015, 24.90405, 24.87781, 
    24.85141, 24.82486, 24.79815, 24.7713, 24.7443, 24.71715, 24.68984, 
    24.66239, 24.63478,
  21.54793, 21.58859, 21.62913, 21.66953, 21.70981, 21.74996, 21.78997, 
    21.82985, 21.86961, 21.90923, 21.94872, 21.98807, 22.0273, 22.06639, 
    22.10535, 22.14418, 22.18287, 22.22144, 22.25986, 22.29816, 22.33632, 
    22.37434, 22.41224, 22.44999, 22.48762, 22.5251, 22.56245, 22.59967, 
    22.63675, 22.67369, 22.7105, 22.74718, 22.78371, 22.82011, 22.85637, 
    22.89249, 22.92848, 22.96432, 23.00003, 23.03561, 23.07104, 23.10633, 
    23.14149, 23.1765, 23.21138, 23.24612, 23.28071, 23.31517, 23.34949, 
    23.38366, 23.4177, 23.45159, 23.48534, 23.51896, 23.55243, 23.58575, 
    23.61894, 23.65198, 23.68488, 23.71764, 23.75025, 23.78272, 23.81505, 
    23.84724, 23.87928, 23.91117, 23.94293, 23.97453, 24.006, 24.03732, 
    24.06849, 24.09952, 24.1304, 24.16113, 24.19172, 24.22217, 24.25247, 
    24.28262, 24.31262, 24.34248, 24.37219, 24.40175, 24.43117, 24.46043, 
    24.48955, 24.51852, 24.54735, 24.57602, 24.60454, 24.63292, 24.66115, 
    24.68922, 24.71715, 24.74493, 24.77255, 24.80003, 24.82736, 24.85453, 
    24.88156, 24.90843, 24.93516, 24.96173, 24.98815, 25.01442, 25.04053, 
    25.0665, 25.09231, 25.11797, 25.14348, 25.16883, 25.19403, 25.21908, 
    25.24397, 25.26871, 25.2933, 25.31773, 25.34201, 25.36613, 25.3901, 
    25.41392, 25.43758, 25.46108, 25.48443, 25.50763, 25.53066, 25.55355, 
    25.57627, 25.59885, 25.62126, 25.64352, 25.66562, 25.68756, 25.70935, 
    25.73098, 25.75246, 25.77378, 25.79493, 25.81594, 25.83678, 25.85746, 
    25.87799, 25.89836, 25.91857, 25.93862, 25.95851, 25.97825, 25.99782, 
    26.01724, 26.03649, 26.05559, 26.07453, 26.0933, 26.11192, 26.13038, 
    26.14867, 26.16681, 26.18478, 26.2026, 26.22025, 26.23775, 26.25508, 
    26.27225, 26.28926, 26.30611, 26.32279, 26.33932, 26.35568, 26.37188, 
    26.38792, 26.4038, 26.41951, 26.43506, 26.45045, 26.46568, 26.48074, 
    26.49564, 26.51037, 26.52495, 26.53936, 26.5536, 26.56769, 26.58161, 
    26.59536, 26.60896, 26.62238, 26.63565, 26.64875, 26.66168, 26.67445, 
    26.68706, 26.6995, 26.71178, 26.72389, 26.73584, 26.74762, 26.75924, 
    26.77069, 26.78197, 26.79309, 26.80405, 26.81484, 26.82546, 26.83592, 
    26.84622, 26.85634, 26.8663, 26.8761, 26.88573, 26.89519, 26.90449, 
    26.91362, 26.92258, 26.93138, 26.94001, 26.94847, 26.95677, 26.9649, 
    26.97286, 26.98066, 26.98829, 26.99575, 27.00304, 27.01017, 27.01713, 
    27.02393, 27.03055, 27.03701, 27.0433, 27.04943, 27.05538, 27.06117, 
    27.06679, 27.07224, 27.07753, 27.08265, 27.0876, 27.09238, 27.09699, 
    27.10144, 27.10572, 27.10983, 27.11377, 27.11754, 27.12115, 27.12459, 
    27.12786, 27.13096, 27.13389, 27.13666, 27.13925, 27.14168, 27.14394, 
    27.14603, 27.14796, 27.14971, 27.1513, 27.15272, 27.15397, 27.15505, 
    27.15596, 27.15671, 27.15728, 27.15769, 27.15793, 27.158, 27.1579, 
    27.15764, 27.1572, 27.1566, 27.15583, 27.15489, 27.15378, 27.1525, 
    27.15106, 27.14944, 27.14766, 27.14571, 27.14359, 27.14131, 27.13885, 
    27.13623, 27.13344, 27.13048, 27.12735, 27.12405, 27.12059, 27.11696, 
    27.11316, 27.10919, 27.10505, 27.10075, 27.09627, 27.09163, 27.08682, 
    27.08185, 27.0767, 27.07139, 27.06591, 27.06026, 27.05445, 27.04847, 
    27.04232, 27.036, 27.02951, 27.02286, 27.01604, 27.00905, 27.0019, 
    26.99458, 26.98709, 26.97943, 26.97161, 26.96362, 26.95547, 26.94714, 
    26.93865, 26.93, 26.92117, 26.91218, 26.90303, 26.89371, 26.88422, 
    26.87456, 26.86474, 26.85475, 26.8446, 26.83428, 26.8238, 26.81314, 
    26.80233, 26.79135, 26.7802, 26.76889, 26.75741, 26.74577, 26.73396, 
    26.72198, 26.70985, 26.69754, 26.68508, 26.67244, 26.65965, 26.64668, 
    26.63356, 26.62027, 26.60682, 26.5932, 26.57942, 26.56547, 26.55136, 
    26.53709, 26.52265, 26.50805, 26.49329, 26.47836, 26.46328, 26.44802, 
    26.43261, 26.41703, 26.40129, 26.38539, 26.36933, 26.3531, 26.33671, 
    26.32016, 26.30345, 26.28658, 26.26954, 26.25235, 26.23499, 26.21747, 
    26.19979, 26.18195, 26.16395, 26.14579, 26.12747, 26.10899, 26.09034, 
    26.07154, 26.05258, 26.03346, 26.01418, 25.99474, 25.97514, 25.95538, 
    25.93546, 25.91538, 25.89515, 25.87475, 25.8542, 25.83349, 25.81262, 
    25.7916, 25.77041, 25.74907, 25.72757, 25.70592, 25.6841, 25.66213, 
    25.64001, 25.61773, 25.59529, 25.57269, 25.54994, 25.52703, 25.50397, 
    25.48075, 25.45737, 25.43385, 25.41016, 25.38632, 25.36233, 25.33818, 
    25.31388, 25.28942, 25.26481, 25.24004, 25.21513, 25.19005, 25.16483, 
    25.13945, 25.11392, 25.08824, 25.0624, 25.03641, 25.01027, 24.98398, 
    24.95754, 24.93094, 24.90419, 24.87729, 24.85025, 24.82305, 24.7957, 
    24.76819, 24.74054,
  21.64854, 21.68927, 21.72987, 21.77034, 21.81067, 21.85088, 21.89096, 
    21.9309, 21.97071, 22.0104, 22.04995, 22.08937, 22.12865, 22.16781, 
    22.20683, 22.24572, 22.28447, 22.32309, 22.36158, 22.39993, 22.43816, 
    22.47624, 22.51419, 22.55201, 22.58969, 22.62724, 22.66465, 22.70192, 
    22.73906, 22.77607, 22.81293, 22.84966, 22.88626, 22.92271, 22.95903, 
    22.99521, 23.03125, 23.06716, 23.10292, 23.13855, 23.17404, 23.20939, 
    23.24461, 23.27968, 23.31461, 23.3494, 23.38406, 23.41857, 23.45294, 
    23.48717, 23.52126, 23.55521, 23.58902, 23.62268, 23.65621, 23.68959, 
    23.72283, 23.75593, 23.78888, 23.82169, 23.85436, 23.88688, 23.91927, 
    23.9515, 23.98359, 24.01554, 24.04735, 24.07901, 24.11053, 24.14189, 
    24.17312, 24.2042, 24.23513, 24.26592, 24.29656, 24.32705, 24.3574, 
    24.3876, 24.41766, 24.44756, 24.47732, 24.50694, 24.5364, 24.56572, 
    24.59488, 24.6239, 24.65277, 24.6815, 24.71007, 24.73849, 24.76677, 
    24.79489, 24.82286, 24.85069, 24.87836, 24.90589, 24.93326, 24.96048, 
    24.98755, 25.01447, 25.04124, 25.06786, 25.09432, 25.12064, 25.1468, 
    25.17281, 25.19866, 25.22437, 25.24992, 25.27531, 25.30056, 25.32565, 
    25.35058, 25.37537, 25.39999, 25.42447, 25.44879, 25.47296, 25.49697, 
    25.52082, 25.54452, 25.56807, 25.59146, 25.61469, 25.63777, 25.66069, 
    25.68346, 25.70607, 25.72852, 25.75082, 25.77296, 25.79494, 25.81677, 
    25.83844, 25.85995, 25.8813, 25.9025, 25.92354, 25.94442, 25.96514, 
    25.9857, 26.00611, 26.02635, 26.04644, 26.06636, 26.08613, 26.10574, 
    26.12519, 26.14448, 26.16361, 26.18258, 26.20139, 26.22004, 26.23853, 
    26.25686, 26.27503, 26.29304, 26.31088, 26.32857, 26.34609, 26.36345, 
    26.38066, 26.3977, 26.41457, 26.43129, 26.44784, 26.46423, 26.48046, 
    26.49653, 26.51244, 26.52818, 26.54376, 26.55917, 26.57442, 26.58951, 
    26.60444, 26.6192, 26.6338, 26.64824, 26.66251, 26.67662, 26.69057, 
    26.70435, 26.71796, 26.73141, 26.7447, 26.75782, 26.77078, 26.78358, 
    26.79621, 26.80867, 26.82097, 26.8331, 26.84507, 26.85687, 26.86851, 
    26.87999, 26.89129, 26.90243, 26.91341, 26.92422, 26.93486, 26.94534, 
    26.95565, 26.9658, 26.97577, 26.98559, 26.99523, 27.00471, 27.01403, 
    27.02317, 27.03215, 27.04096, 27.04961, 27.05809, 27.0664, 27.07455, 
    27.08252, 27.09033, 27.09798, 27.10545, 27.11276, 27.1199, 27.12687, 
    27.13368, 27.14032, 27.14679, 27.15309, 27.15923, 27.16519, 27.17099, 
    27.17662, 27.18209, 27.18738, 27.19251, 27.19747, 27.20226, 27.20688, 
    27.21134, 27.21562, 27.21974, 27.22369, 27.22747, 27.23108, 27.23453, 
    27.2378, 27.24091, 27.24385, 27.24662, 27.24922, 27.25165, 27.25392, 
    27.25601, 27.25794, 27.2597, 27.26129, 27.26271, 27.26396, 27.26504, 
    27.26596, 27.2667, 27.26728, 27.26769, 27.26793, 27.268, 27.2679, 
    27.26764, 27.2672, 27.2666, 27.26582, 27.26488, 27.26377, 27.26249, 
    27.26105, 27.25943, 27.25764, 27.25569, 27.25357, 27.25128, 27.24882, 
    27.24619, 27.24339, 27.24043, 27.2373, 27.23399, 27.23052, 27.22688, 
    27.22307, 27.2191, 27.21495, 27.21064, 27.20616, 27.20151, 27.1967, 
    27.19171, 27.18656, 27.18123, 27.17575, 27.17009, 27.16426, 27.15827, 
    27.15211, 27.14578, 27.13928, 27.13262, 27.12578, 27.11878, 27.11162, 
    27.10428, 27.09678, 27.08911, 27.08127, 27.07327, 27.0651, 27.05676, 
    27.04825, 27.03958, 27.03074, 27.02174, 27.01256, 27.00322, 26.99372, 
    26.98405, 26.97421, 26.9642, 26.95403, 26.94369, 26.93319, 26.92252, 
    26.91168, 26.90068, 26.88951, 26.87818, 26.86668, 26.85502, 26.84319, 
    26.83119, 26.81903, 26.80671, 26.79422, 26.78156, 26.76874, 26.75576, 
    26.74261, 26.7293, 26.71582, 26.70218, 26.68837, 26.6744, 26.66026, 
    26.64597, 26.63151, 26.61688, 26.60209, 26.58714, 26.57202, 26.55674, 
    26.5413, 26.5257, 26.50993, 26.494, 26.47791, 26.46165, 26.44523, 
    26.42866, 26.41191, 26.39501, 26.37794, 26.36072, 26.34333, 26.32578, 
    26.30807, 26.2902, 26.27217, 26.25397, 26.23562, 26.2171, 26.19843, 
    26.17959, 26.1606, 26.14144, 26.12213, 26.10265, 26.08302, 26.06322, 
    26.04327, 26.02316, 26.00289, 25.98246, 25.96187, 25.94112, 25.92022, 
    25.89916, 25.87794, 25.85656, 25.83502, 25.81333, 25.79148, 25.76947, 
    25.7473, 25.72498, 25.7025, 25.67987, 25.65708, 25.63413, 25.61103, 
    25.58777, 25.56435, 25.54078, 25.51706, 25.49318, 25.46914, 25.44495, 
    25.42061, 25.39611, 25.37146, 25.34665, 25.32169, 25.29657, 25.27131, 
    25.24588, 25.22031, 25.19458, 25.1687, 25.14267, 25.11648, 25.09015, 
    25.06366, 25.03702, 25.01023, 24.98328, 24.95619, 24.92894, 24.90154, 
    24.87399, 24.8463,
  21.74915, 21.78994, 21.8306, 21.87112, 21.91152, 21.95179, 21.99193, 
    22.03194, 22.07181, 22.11156, 22.15117, 22.19065, 22.22999, 22.26921, 
    22.30829, 22.34724, 22.38605, 22.42474, 22.46329, 22.5017, 22.53998, 
    22.57813, 22.61614, 22.65401, 22.69175, 22.72936, 22.76683, 22.80416, 
    22.84136, 22.87842, 22.91535, 22.95214, 22.98879, 23.0253, 23.06168, 
    23.09792, 23.13402, 23.16998, 23.2058, 23.24149, 23.27703, 23.31244, 
    23.34771, 23.38284, 23.41783, 23.45268, 23.48739, 23.52195, 23.55638, 
    23.59067, 23.62481, 23.65882, 23.69268, 23.7264, 23.75998, 23.79342, 
    23.82671, 23.85986, 23.89287, 23.92573, 23.95845, 23.99103, 24.02347, 
    24.05576, 24.0879, 24.11991, 24.15176, 24.18347, 24.21504, 24.24646, 
    24.27774, 24.30887, 24.33985, 24.37069, 24.40138, 24.43193, 24.46233, 
    24.49258, 24.52268, 24.55264, 24.58245, 24.61211, 24.64162, 24.67099, 
    24.70021, 24.72927, 24.75819, 24.78696, 24.81558, 24.84406, 24.87238, 
    24.90055, 24.92857, 24.95644, 24.98416, 25.01173, 25.03915, 25.06642, 
    25.09354, 25.1205, 25.14732, 25.17398, 25.20049, 25.22685, 25.25305, 
    25.27911, 25.30501, 25.33075, 25.35635, 25.38179, 25.40708, 25.43221, 
    25.45719, 25.48201, 25.50669, 25.5312, 25.55556, 25.57977, 25.60382, 
    25.62772, 25.65146, 25.67505, 25.69848, 25.72175, 25.74487, 25.76783, 
    25.79064, 25.81329, 25.83578, 25.85812, 25.8803, 25.90232, 25.92418, 
    25.94589, 25.96744, 25.98883, 26.01006, 26.03114, 26.05205, 26.07281, 
    26.09341, 26.11385, 26.13413, 26.15425, 26.17421, 26.19402, 26.21366, 
    26.23314, 26.25247, 26.27163, 26.29063, 26.30948, 26.32816, 26.34668, 
    26.36504, 26.38324, 26.40128, 26.41916, 26.43688, 26.45443, 26.47183, 
    26.48906, 26.50613, 26.52304, 26.53978, 26.55636, 26.57279, 26.58904, 
    26.60514, 26.62107, 26.63684, 26.65245, 26.66789, 26.68317, 26.69829, 
    26.71324, 26.72803, 26.74266, 26.75712, 26.77142, 26.78555, 26.79952, 
    26.81333, 26.82697, 26.84044, 26.85375, 26.8669, 26.87988, 26.8927, 
    26.90535, 26.91784, 26.93016, 26.94231, 26.9543, 26.96613, 26.97779, 
    26.98928, 27.00061, 27.01177, 27.02276, 27.03359, 27.04426, 27.05475, 
    27.06508, 27.07525, 27.08524, 27.09507, 27.10474, 27.11423, 27.12356, 
    27.13273, 27.14172, 27.15055, 27.15921, 27.16771, 27.17603, 27.18419, 
    27.19219, 27.20001, 27.20767, 27.21516, 27.22248, 27.22963, 27.23662, 
    27.24344, 27.25009, 27.25657, 27.26288, 27.26903, 27.27501, 27.28082, 
    27.28646, 27.29193, 27.29724, 27.30237, 27.30734, 27.31214, 27.31677, 
    27.32123, 27.32553, 27.32965, 27.33361, 27.33739, 27.34101, 27.34447, 
    27.34775, 27.35086, 27.3538, 27.35658, 27.35918, 27.36162, 27.36389, 
    27.36599, 27.36792, 27.36968, 27.37127, 27.3727, 27.37395, 27.37504, 
    27.37595, 27.3767, 27.37728, 27.37769, 27.37793, 27.378, 27.3779, 
    27.37763, 27.3772, 27.37659, 27.37582, 27.37488, 27.37376, 27.37248, 
    27.37103, 27.36941, 27.36763, 27.36567, 27.36354, 27.36125, 27.35878, 
    27.35615, 27.35335, 27.35038, 27.34724, 27.34393, 27.34045, 27.33681, 
    27.33299, 27.32901, 27.32486, 27.32054, 27.31605, 27.31139, 27.30656, 
    27.30157, 27.29641, 27.29108, 27.28558, 27.27991, 27.27407, 27.26807, 
    27.2619, 27.25555, 27.24905, 27.24237, 27.23553, 27.22851, 27.22133, 
    27.21398, 27.20647, 27.19878, 27.19093, 27.18291, 27.17473, 27.16637, 
    27.15785, 27.14917, 27.14031, 27.13129, 27.1221, 27.11274, 27.10322, 
    27.09353, 27.08367, 27.07365, 27.06346, 27.0531, 27.04258, 27.03189, 
    27.02104, 27.01002, 26.99883, 26.98747, 26.97595, 26.96427, 26.95242, 
    26.9404, 26.92822, 26.91587, 26.90336, 26.89068, 26.87784, 26.86483, 
    26.85166, 26.83832, 26.82482, 26.81115, 26.79732, 26.78333, 26.76917, 
    26.75484, 26.74036, 26.7257, 26.71089, 26.69591, 26.68077, 26.66546, 
    26.64999, 26.63436, 26.61856, 26.6026, 26.58648, 26.5702, 26.55375, 
    26.53714, 26.52037, 26.50344, 26.48634, 26.46909, 26.45167, 26.43409, 
    26.41634, 26.39844, 26.38038, 26.36215, 26.34376, 26.32522, 26.30651, 
    26.28764, 26.26861, 26.24942, 26.23007, 26.21056, 26.1909, 26.17107, 
    26.15108, 26.13093, 26.11062, 26.09016, 26.06954, 26.04875, 26.02781, 
    26.00671, 25.98545, 25.96404, 25.94246, 25.92073, 25.89884, 25.8768, 
    25.8546, 25.83223, 25.80972, 25.78704, 25.76421, 25.74122, 25.71808, 
    25.69478, 25.67133, 25.64772, 25.62395, 25.60003, 25.57595, 25.55172, 
    25.52733, 25.50279, 25.4781, 25.45325, 25.42824, 25.40309, 25.37778, 
    25.35231, 25.32669, 25.30092, 25.275, 25.24892, 25.22269, 25.19631, 
    25.16977, 25.14309, 25.11625, 25.08926, 25.06212, 25.03483, 25.00738, 
    24.97979, 24.95204,
  21.84973, 21.89058, 21.93131, 21.9719, 22.01236, 22.05269, 22.09289, 
    22.13296, 22.1729, 22.2127, 22.25237, 22.29191, 22.33132, 22.3706, 
    22.40974, 22.44875, 22.48763, 22.52637, 22.56498, 22.60345, 22.64179, 
    22.68, 22.71807, 22.756, 22.79381, 22.83147, 22.869, 22.90639, 22.94365, 
    22.98077, 23.01775, 23.0546, 23.09131, 23.12788, 23.16431, 23.20061, 
    23.23677, 23.27279, 23.30867, 23.34441, 23.38002, 23.41548, 23.45081, 
    23.48599, 23.52104, 23.55594, 23.59071, 23.62533, 23.65981, 23.69415, 
    23.72836, 23.76241, 23.79633, 23.83011, 23.86374, 23.89723, 23.93058, 
    23.96379, 23.99685, 24.02977, 24.06254, 24.09517, 24.12766, 24.16, 
    24.1922, 24.22426, 24.25617, 24.28793, 24.31955, 24.35102, 24.38235, 
    24.41353, 24.44457, 24.47546, 24.5062, 24.5368, 24.56725, 24.59755, 
    24.6277, 24.65771, 24.68757, 24.71728, 24.74684, 24.77626, 24.80552, 
    24.83464, 24.86361, 24.89242, 24.92109, 24.94961, 24.97798, 25.0062, 
    25.03427, 25.06219, 25.08996, 25.11757, 25.14504, 25.17235, 25.19952, 
    25.22653, 25.25339, 25.2801, 25.30665, 25.33305, 25.3593, 25.3854, 
    25.41135, 25.43714, 25.46277, 25.48826, 25.51359, 25.53876, 25.56379, 
    25.58866, 25.61337, 25.63793, 25.66233, 25.68658, 25.71067, 25.73461, 
    25.7584, 25.78202, 25.80549, 25.82881, 25.85197, 25.87497, 25.89781, 
    25.9205, 25.94304, 25.96541, 25.98763, 26.00969, 26.03159, 26.05333, 
    26.07492, 26.09635, 26.11762, 26.13873, 26.15968, 26.18048, 26.20111, 
    26.22159, 26.2419, 26.26206, 26.28206, 26.3019, 26.32157, 26.34109, 
    26.36045, 26.37965, 26.39868, 26.41756, 26.43628, 26.45483, 26.47322, 
    26.49146, 26.50953, 26.52744, 26.54519, 26.56277, 26.5802, 26.59746, 
    26.61456, 26.6315, 26.64827, 26.66488, 26.68134, 26.69762, 26.71375, 
    26.72971, 26.7455, 26.76114, 26.77661, 26.79192, 26.80706, 26.82204, 
    26.83686, 26.85151, 26.866, 26.88032, 26.89448, 26.90848, 26.9223, 
    26.93597, 26.94947, 26.9628, 26.97598, 26.98898, 27.00182, 27.01449, 
    27.027, 27.03935, 27.05153, 27.06354, 27.07538, 27.08706, 27.09858, 
    27.10992, 27.12111, 27.13212, 27.14297, 27.15365, 27.16417, 27.17451, 
    27.1847, 27.19471, 27.20456, 27.21424, 27.22375, 27.2331, 27.24228, 
    27.25129, 27.26014, 27.26881, 27.27732, 27.28567, 27.29384, 27.30185, 
    27.30969, 27.31736, 27.32486, 27.3322, 27.33936, 27.34636, 27.35319, 
    27.35985, 27.36635, 27.37267, 27.37883, 27.38482, 27.39064, 27.39629, 
    27.40177, 27.40709, 27.41223, 27.41721, 27.42202, 27.42666, 27.43113, 
    27.43543, 27.43956, 27.44353, 27.44732, 27.45095, 27.4544, 27.45769, 
    27.46081, 27.46376, 27.46654, 27.46915, 27.47159, 27.47386, 27.47597, 
    27.4779, 27.47967, 27.48126, 27.48269, 27.48394, 27.48503, 27.48595, 
    27.4867, 27.48728, 27.48769, 27.48793, 27.488, 27.4879, 27.48763, 
    27.4872, 27.48659, 27.48582, 27.48487, 27.48376, 27.48247, 27.48102, 
    27.4794, 27.47761, 27.47565, 27.47352, 27.47122, 27.46875, 27.46611, 
    27.4633, 27.46033, 27.45718, 27.45387, 27.45038, 27.44673, 27.44291, 
    27.43892, 27.43476, 27.43043, 27.42594, 27.42127, 27.41644, 27.41143, 
    27.40626, 27.40092, 27.39541, 27.38973, 27.38388, 27.37787, 27.37168, 
    27.36533, 27.35881, 27.35212, 27.34526, 27.33824, 27.33105, 27.32368, 
    27.31615, 27.30846, 27.30059, 27.29256, 27.28436, 27.27599, 27.26745, 
    27.25875, 27.24988, 27.24084, 27.23163, 27.22226, 27.21272, 27.20301, 
    27.19314, 27.1831, 27.17289, 27.16251, 27.15197, 27.14126, 27.13039, 
    27.11935, 27.10814, 27.09677, 27.08523, 27.07352, 27.06165, 27.04961, 
    27.03741, 27.02504, 27.0125, 26.9998, 26.98693, 26.9739, 26.96071, 
    26.94735, 26.93382, 26.92013, 26.90627, 26.89225, 26.87807, 26.86372, 
    26.8492, 26.83453, 26.81968, 26.80468, 26.78951, 26.77417, 26.75868, 
    26.74302, 26.72719, 26.71121, 26.69506, 26.67874, 26.66227, 26.64563, 
    26.62883, 26.61186, 26.59474, 26.57745, 26.56, 26.54239, 26.52462, 
    26.50668, 26.48858, 26.47033, 26.45191, 26.43333, 26.41459, 26.39568, 
    26.37662, 26.3574, 26.33801, 26.31847, 26.29877, 26.27891, 26.25888, 
    26.2387, 26.21836, 26.19786, 26.1772, 26.15638, 26.1354, 26.11426, 
    26.09297, 26.07151, 26.0499, 26.02814, 26.00621, 25.98412, 25.96188, 
    25.93948, 25.91693, 25.89421, 25.87134, 25.84831, 25.82513, 25.80179, 
    25.7783, 25.75464, 25.73084, 25.70687, 25.68276, 25.65848, 25.63405, 
    25.60947, 25.58473, 25.55984, 25.53479, 25.50959, 25.48424, 25.45873, 
    25.43307, 25.40725, 25.38128, 25.35516, 25.32889, 25.30246, 25.27588, 
    25.24915, 25.22227, 25.19523, 25.16804, 25.14071, 25.11321, 25.08558, 
    25.05778,
  21.95031, 21.99122, 22.03201, 22.07266, 22.11318, 22.15358, 22.19384, 
    22.23397, 22.27397, 22.31383, 22.35357, 22.39317, 22.43264, 22.47198, 
    22.51118, 22.55025, 22.58919, 22.62799, 22.66666, 22.70519, 22.74359, 
    22.78186, 22.81999, 22.85798, 22.89584, 22.93357, 22.97116, 23.00861, 
    23.04592, 23.0831, 23.12015, 23.15705, 23.19382, 23.23045, 23.26694, 
    23.3033, 23.33951, 23.37559, 23.41153, 23.44733, 23.48299, 23.51851, 
    23.55389, 23.58913, 23.62423, 23.65919, 23.69402, 23.72869, 23.76323, 
    23.79763, 23.83189, 23.866, 23.89997, 23.9338, 23.96749, 24.00104, 
    24.03444, 24.0677, 24.10081, 24.13379, 24.16662, 24.1993, 24.23184, 
    24.26424, 24.29649, 24.3286, 24.36056, 24.39238, 24.42405, 24.45557, 
    24.48695, 24.51819, 24.54927, 24.58021, 24.61101, 24.64165, 24.67216, 
    24.70251, 24.73271, 24.76277, 24.79268, 24.82244, 24.85205, 24.88151, 
    24.91083, 24.93999, 24.96901, 24.99788, 25.02659, 25.05516, 25.08358, 
    25.11185, 25.13996, 25.16793, 25.19574, 25.22341, 25.25092, 25.27828, 
    25.30549, 25.33255, 25.35945, 25.3862, 25.4128, 25.43925, 25.46555, 
    25.49169, 25.51768, 25.54351, 25.56919, 25.59472, 25.6201, 25.64532, 
    25.67038, 25.69529, 25.72005, 25.74465, 25.76909, 25.79338, 25.81752, 
    25.8415, 25.86532, 25.88899, 25.9125, 25.93586, 25.95906, 25.9821, 
    26.00498, 26.02771, 26.05028, 26.0727, 26.09495, 26.11705, 26.13899, 
    26.16077, 26.1824, 26.20386, 26.22517, 26.24632, 26.26731, 26.28814, 
    26.30881, 26.32932, 26.34967, 26.36987, 26.3899, 26.40977, 26.42948, 
    26.44904, 26.46843, 26.48766, 26.50673, 26.52564, 26.54439, 26.56297, 
    26.5814, 26.59967, 26.61777, 26.63571, 26.65349, 26.67111, 26.68856, 
    26.70586, 26.72299, 26.73995, 26.75676, 26.7734, 26.78988, 26.8062, 
    26.82235, 26.83834, 26.85417, 26.86983, 26.88533, 26.90066, 26.91583, 
    26.93084, 26.94568, 26.96036, 26.97487, 26.98922, 27.00341, 27.01743, 
    27.03128, 27.04497, 27.05849, 27.07185, 27.08505, 27.09808, 27.11094, 
    27.12364, 27.13617, 27.14853, 27.16073, 27.17277, 27.18463, 27.19633, 
    27.20787, 27.21924, 27.23044, 27.24147, 27.25234, 27.26304, 27.27358, 
    27.28395, 27.29415, 27.30418, 27.31404, 27.32374, 27.33327, 27.34264, 
    27.35183, 27.36086, 27.36972, 27.37842, 27.38694, 27.3953, 27.40349, 
    27.41151, 27.41936, 27.42705, 27.43456, 27.44191, 27.44909, 27.4561, 
    27.46295, 27.46962, 27.47613, 27.48246, 27.48863, 27.49463, 27.50046, 
    27.50612, 27.51162, 27.51694, 27.52209, 27.52708, 27.5319, 27.53655, 
    27.54103, 27.54533, 27.54947, 27.55345, 27.55725, 27.56088, 27.56434, 
    27.56764, 27.57076, 27.57372, 27.5765, 27.57911, 27.58156, 27.58384, 
    27.58595, 27.58788, 27.58965, 27.59125, 27.59268, 27.59394, 27.59503, 
    27.59595, 27.59669, 27.59728, 27.59769, 27.59793, 27.598, 27.5979, 
    27.59763, 27.5972, 27.59659, 27.59581, 27.59487, 27.59375, 27.59246, 
    27.59101, 27.58938, 27.58759, 27.58562, 27.58349, 27.58119, 27.57871, 
    27.57607, 27.57326, 27.57028, 27.56713, 27.56381, 27.56032, 27.55666, 
    27.55283, 27.54883, 27.54466, 27.54033, 27.53582, 27.53115, 27.5263, 
    27.52129, 27.51611, 27.51076, 27.50524, 27.49955, 27.49369, 27.48767, 
    27.48147, 27.47511, 27.46857, 27.46187, 27.45501, 27.44797, 27.44076, 
    27.43339, 27.42584, 27.41813, 27.41025, 27.4022, 27.39399, 27.3856, 
    27.37705, 27.36833, 27.35945, 27.35039, 27.34117, 27.33178, 27.32222, 
    27.31249, 27.3026, 27.29254, 27.28232, 27.27192, 27.26136, 27.25063, 
    27.23974, 27.22868, 27.21745, 27.20606, 27.19449, 27.18277, 27.17087, 
    27.15881, 27.14659, 27.1342, 27.12164, 27.10892, 27.09603, 27.08297, 
    27.06975, 27.05637, 27.04282, 27.0291, 27.01522, 27.00117, 26.98696, 
    26.97259, 26.95805, 26.94334, 26.92848, 26.91344, 26.89825, 26.88289, 
    26.86736, 26.85167, 26.83582, 26.81981, 26.80363, 26.78728, 26.77078, 
    26.75411, 26.73728, 26.72029, 26.70313, 26.68581, 26.66833, 26.65069, 
    26.63288, 26.61492, 26.59679, 26.5785, 26.56005, 26.54143, 26.52266, 
    26.50372, 26.48463, 26.46537, 26.44595, 26.42638, 26.40664, 26.38674, 
    26.36668, 26.34646, 26.32609, 26.30555, 26.28485, 26.264, 26.24298, 
    26.22181, 26.20048, 26.17899, 26.15734, 26.13553, 26.11357, 26.09144, 
    26.06916, 26.04672, 26.02413, 26.00138, 25.97846, 25.9554, 25.93217, 
    25.90879, 25.88526, 25.86157, 25.83772, 25.81371, 25.78955, 25.76524, 
    25.74077, 25.71614, 25.69136, 25.66643, 25.64134, 25.61609, 25.59069, 
    25.56514, 25.53944, 25.51358, 25.48756, 25.4614, 25.43508, 25.40861, 
    25.38198, 25.35521, 25.32828, 25.3012, 25.27396, 25.24658, 25.21904, 
    25.19135, 25.16351,
  22.05087, 22.09184, 22.13269, 22.17341, 22.21399, 22.25445, 22.29477, 
    22.33496, 22.37502, 22.41495, 22.45475, 22.49441, 22.53394, 22.57334, 
    22.6126, 22.65174, 22.69073, 22.7296, 22.76832, 22.80692, 22.84538, 
    22.88371, 22.9219, 22.95995, 22.99787, 23.03565, 23.0733, 23.11081, 
    23.14819, 23.18542, 23.22252, 23.25949, 23.29631, 23.333, 23.36955, 
    23.40597, 23.44224, 23.47837, 23.51437, 23.55023, 23.58595, 23.62152, 
    23.65696, 23.69226, 23.72742, 23.76244, 23.79731, 23.83205, 23.86664, 
    23.9011, 23.93541, 23.96958, 24.0036, 24.03749, 24.07123, 24.10483, 
    24.13829, 24.1716, 24.20477, 24.2378, 24.27068, 24.30342, 24.33602, 
    24.36847, 24.40077, 24.43293, 24.46494, 24.49681, 24.52854, 24.56011, 
    24.59155, 24.62283, 24.65397, 24.68496, 24.71581, 24.7465, 24.77706, 
    24.80746, 24.83771, 24.86782, 24.89778, 24.92759, 24.95725, 24.98676, 
    25.01613, 25.04534, 25.07441, 25.10332, 25.13209, 25.1607, 25.18917, 
    25.21748, 25.24565, 25.27366, 25.30152, 25.32923, 25.35679, 25.3842, 
    25.41145, 25.43856, 25.46551, 25.49231, 25.51895, 25.54544, 25.57178, 
    25.59797, 25.624, 25.64988, 25.67561, 25.70118, 25.7266, 25.75186, 
    25.77697, 25.80192, 25.82672, 25.85136, 25.87585, 25.90018, 25.92436, 
    25.94838, 25.97225, 25.99595, 26.01951, 26.0429, 26.06614, 26.08922, 
    26.11215, 26.13492, 26.15753, 26.17998, 26.20227, 26.22441, 26.24639, 
    26.26821, 26.28987, 26.31137, 26.33272, 26.3539, 26.37493, 26.3958, 
    26.4165, 26.43705, 26.45744, 26.47767, 26.49773, 26.51764, 26.53739, 
    26.55698, 26.5764, 26.59567, 26.61477, 26.63371, 26.6525, 26.67112, 
    26.68958, 26.70787, 26.72601, 26.74398, 26.76179, 26.77944, 26.79693, 
    26.81425, 26.83141, 26.84841, 26.86524, 26.88192, 26.89842, 26.91477, 
    26.93095, 26.94697, 26.96282, 26.97851, 26.99404, 27.0094, 27.0246, 
    27.03963, 27.0545, 27.06921, 27.08375, 27.09812, 27.11233, 27.12638, 
    27.14025, 27.15397, 27.16752, 27.1809, 27.19412, 27.20717, 27.22006, 
    27.23278, 27.24533, 27.25772, 27.26994, 27.282, 27.29388, 27.3056, 
    27.31716, 27.32855, 27.33977, 27.35083, 27.36171, 27.37243, 27.38299, 
    27.39337, 27.40359, 27.41364, 27.42353, 27.43324, 27.44279, 27.45217, 
    27.46139, 27.47043, 27.47931, 27.48802, 27.49656, 27.50493, 27.51313, 
    27.52117, 27.52904, 27.53674, 27.54427, 27.55163, 27.55882, 27.56584, 
    27.5727, 27.57939, 27.5859, 27.59225, 27.59843, 27.60444, 27.61028, 
    27.61596, 27.62146, 27.62679, 27.63196, 27.63695, 27.64178, 27.64643, 
    27.65092, 27.65524, 27.65939, 27.66336, 27.66717, 27.67081, 27.67428, 
    27.67758, 27.68071, 27.68367, 27.68646, 27.68908, 27.69153, 27.69381, 
    27.69592, 27.69786, 27.69963, 27.70124, 27.70267, 27.70393, 27.70502, 
    27.70594, 27.70669, 27.70728, 27.70769, 27.70793, 27.708, 27.7079, 
    27.70763, 27.70719, 27.70659, 27.70581, 27.70486, 27.70374, 27.70245, 
    27.70099, 27.69937, 27.69757, 27.6956, 27.69346, 27.69115, 27.68868, 
    27.68603, 27.68321, 27.68023, 27.67707, 27.67374, 27.67025, 27.66658, 
    27.66275, 27.65874, 27.65457, 27.65022, 27.64571, 27.64103, 27.63617, 
    27.63115, 27.62596, 27.6206, 27.61507, 27.60937, 27.6035, 27.59747, 
    27.59126, 27.58488, 27.57834, 27.57163, 27.56474, 27.55769, 27.55047, 
    27.54309, 27.53553, 27.5278, 27.51991, 27.51185, 27.50362, 27.49522, 
    27.48665, 27.47791, 27.46901, 27.45994, 27.4507, 27.44129, 27.43172, 
    27.42198, 27.41207, 27.40199, 27.39174, 27.38133, 27.37075, 27.36, 
    27.34909, 27.33801, 27.32676, 27.31534, 27.30376, 27.29202, 27.2801, 
    27.26802, 27.25577, 27.24336, 27.23078, 27.21803, 27.20512, 27.19204, 
    27.1788, 27.16539, 27.15181, 27.13807, 27.12417, 27.11009, 27.09586, 
    27.08146, 27.06689, 27.05216, 27.03727, 27.02221, 27.00698, 26.99159, 
    26.97604, 26.96033, 26.94445, 26.9284, 26.9122, 26.89582, 26.87929, 
    26.86259, 26.84573, 26.82871, 26.81152, 26.79417, 26.77666, 26.75899, 
    26.74115, 26.72315, 26.70499, 26.68667, 26.66818, 26.64954, 26.63073, 
    26.61176, 26.59263, 26.57334, 26.55389, 26.53428, 26.5145, 26.49457, 
    26.47448, 26.45422, 26.43381, 26.41324, 26.39251, 26.37161, 26.35056, 
    26.32935, 26.30798, 26.28645, 26.26477, 26.24292, 26.22092, 26.19876, 
    26.17644, 26.15396, 26.13132, 26.10853, 26.08558, 26.06248, 26.03921, 
    26.01579, 25.99221, 25.96848, 25.94459, 25.92055, 25.89635, 25.87199, 
    25.84748, 25.82281, 25.79799, 25.77301, 25.74787, 25.72259, 25.69715, 
    25.67155, 25.6458, 25.6199, 25.59384, 25.56763, 25.54126, 25.51475, 
    25.48808, 25.46125, 25.43428, 25.40715, 25.37987, 25.35244, 25.32486, 
    25.29712, 25.26924,
  22.15141, 22.19245, 22.23336, 22.27414, 22.31479, 22.3553, 22.39569, 
    22.43594, 22.47606, 22.51606, 22.55591, 22.59564, 22.63523, 22.67469, 
    22.71401, 22.75321, 22.79226, 22.83119, 22.86998, 22.90863, 22.94715, 
    22.98554, 23.02379, 23.0619, 23.09988, 23.13773, 23.17543, 23.213, 
    23.25044, 23.28773, 23.32489, 23.36192, 23.3988, 23.43555, 23.47215, 
    23.50863, 23.54496, 23.58115, 23.6172, 23.65312, 23.68889, 23.72453, 
    23.76002, 23.79538, 23.83059, 23.86567, 23.9006, 23.93539, 23.97004, 
    24.00455, 24.03892, 24.07314, 24.10723, 24.14117, 24.17496, 24.20862, 
    24.24213, 24.2755, 24.30872, 24.3418, 24.37474, 24.40753, 24.44018, 
    24.47268, 24.50504, 24.53725, 24.56932, 24.60124, 24.63302, 24.66465, 
    24.69613, 24.72747, 24.75866, 24.7897, 24.8206, 24.85135, 24.88195, 
    24.9124, 24.94271, 24.97286, 25.00287, 25.03273, 25.06244, 25.092, 
    25.12142, 25.15068, 25.17979, 25.20876, 25.23757, 25.26624, 25.29475, 
    25.32311, 25.35132, 25.37938, 25.40729, 25.43505, 25.46265, 25.49011, 
    25.51741, 25.54456, 25.57156, 25.5984, 25.62509, 25.65163, 25.67801, 
    25.70424, 25.73032, 25.75624, 25.78201, 25.80763, 25.83309, 25.8584, 
    25.88355, 25.90854, 25.93339, 25.95807, 25.9826, 26.00698, 26.03119, 
    26.05526, 26.07916, 26.10291, 26.1265, 26.14994, 26.17322, 26.19634, 
    26.21931, 26.24212, 26.26476, 26.28725, 26.30959, 26.33176, 26.35378, 
    26.37564, 26.39734, 26.41888, 26.44026, 26.46148, 26.48255, 26.50345, 
    26.52419, 26.54478, 26.5652, 26.58546, 26.60557, 26.62551, 26.64529, 
    26.66491, 26.68437, 26.70367, 26.72281, 26.74179, 26.7606, 26.77925, 
    26.79774, 26.81607, 26.83424, 26.85225, 26.87009, 26.88777, 26.90529, 
    26.92264, 26.93983, 26.95686, 26.97372, 26.99043, 27.00696, 27.02334, 
    27.03955, 27.0556, 27.07148, 27.0872, 27.10275, 27.11814, 27.13337, 
    27.14843, 27.16332, 27.17805, 27.19262, 27.20702, 27.22125, 27.23532, 
    27.24923, 27.26297, 27.27654, 27.28995, 27.30319, 27.31626, 27.32917, 
    27.34192, 27.35449, 27.3669, 27.37914, 27.39122, 27.40313, 27.41488, 
    27.42645, 27.43786, 27.4491, 27.46018, 27.47108, 27.48182, 27.4924, 
    27.5028, 27.51304, 27.52311, 27.53301, 27.54275, 27.55231, 27.56171, 
    27.57094, 27.58, 27.58889, 27.59762, 27.60617, 27.61456, 27.62278, 
    27.63083, 27.63871, 27.64642, 27.65397, 27.66134, 27.66855, 27.67558, 
    27.68245, 27.68915, 27.69568, 27.70204, 27.70823, 27.71425, 27.72011, 
    27.72579, 27.7313, 27.73664, 27.74182, 27.74682, 27.75166, 27.75632, 
    27.76082, 27.76514, 27.7693, 27.77328, 27.7771, 27.78074, 27.78422, 
    27.78753, 27.79066, 27.79362, 27.79642, 27.79905, 27.8015, 27.80379, 
    27.8059, 27.80785, 27.80962, 27.81122, 27.81266, 27.81392, 27.81502, 
    27.81594, 27.81669, 27.81727, 27.81769, 27.81793, 27.818, 27.8179, 
    27.81763, 27.81719, 27.81658, 27.8158, 27.81485, 27.81373, 27.81244, 
    27.81098, 27.80935, 27.80755, 27.80558, 27.80344, 27.80112, 27.79864, 
    27.79599, 27.79317, 27.79018, 27.78701, 27.78368, 27.78018, 27.77651, 
    27.77266, 27.76865, 27.76447, 27.76012, 27.75559, 27.7509, 27.74604, 
    27.74101, 27.73581, 27.73044, 27.7249, 27.71919, 27.71331, 27.70726, 
    27.70105, 27.69466, 27.6881, 27.68138, 27.67448, 27.66742, 27.66019, 
    27.65278, 27.64521, 27.63748, 27.62957, 27.62149, 27.61325, 27.60483, 
    27.59625, 27.5875, 27.57858, 27.56949, 27.56023, 27.55081, 27.54122, 
    27.53146, 27.52153, 27.51143, 27.50117, 27.49074, 27.48014, 27.46937, 
    27.45844, 27.44734, 27.43607, 27.42463, 27.41303, 27.40126, 27.38932, 
    27.37722, 27.36495, 27.35251, 27.33991, 27.32714, 27.31421, 27.30111, 
    27.28784, 27.2744, 27.26081, 27.24704, 27.23311, 27.21901, 27.20475, 
    27.19032, 27.17573, 27.16098, 27.14606, 27.13097, 27.11572, 27.1003, 
    27.08472, 27.06898, 27.05307, 27.037, 27.02076, 27.00436, 26.98779, 
    26.97107, 26.95418, 26.93712, 26.91991, 26.90253, 26.88498, 26.86728, 
    26.84941, 26.83138, 26.81319, 26.79483, 26.77631, 26.75764, 26.73879, 
    26.71979, 26.70063, 26.6813, 26.66182, 26.64217, 26.62237, 26.6024, 
    26.58227, 26.56198, 26.54153, 26.52092, 26.50015, 26.47922, 26.45814, 
    26.43689, 26.41548, 26.39392, 26.37219, 26.35031, 26.32827, 26.30607, 
    26.28371, 26.26119, 26.23852, 26.21568, 26.1927, 26.16955, 26.14625, 
    26.12278, 26.09917, 26.07539, 26.05146, 26.02737, 26.00313, 25.97873, 
    25.95418, 25.92947, 25.9046, 25.87958, 25.8544, 25.82907, 25.80359, 
    25.77795, 25.75216, 25.72621, 25.70011, 25.67385, 25.64744, 25.62088, 
    25.59416, 25.5673, 25.54027, 25.5131, 25.48577, 25.4583, 25.43067, 
    25.40289, 25.37495,
  22.25194, 22.29305, 22.33402, 22.37486, 22.41557, 22.45615, 22.4966, 
    22.53691, 22.5771, 22.61715, 22.65707, 22.69685, 22.73651, 22.77603, 
    22.81541, 22.85467, 22.89378, 22.93277, 22.97162, 23.01034, 23.04892, 
    23.08736, 23.12567, 23.16385, 23.20189, 23.23979, 23.27755, 23.31518, 
    23.35268, 23.39003, 23.42725, 23.46433, 23.50127, 23.53808, 23.57475, 
    23.61127, 23.64766, 23.68391, 23.72002, 23.756, 23.79183, 23.82752, 
    23.86307, 23.89849, 23.93376, 23.96889, 24.00388, 24.03872, 24.07343, 
    24.10799, 24.14242, 24.1767, 24.21084, 24.24483, 24.27868, 24.31239, 
    24.34596, 24.37938, 24.41266, 24.4458, 24.47878, 24.51163, 24.54433, 
    24.57689, 24.6093, 24.64157, 24.67369, 24.70566, 24.73749, 24.76917, 
    24.8007, 24.83209, 24.86333, 24.89443, 24.92538, 24.95618, 24.98683, 
    25.01733, 25.04769, 25.0779, 25.10796, 25.13787, 25.16763, 25.19724, 
    25.2267, 25.25601, 25.28518, 25.31419, 25.34305, 25.37176, 25.40032, 
    25.42873, 25.45699, 25.4851, 25.51305, 25.54086, 25.56851, 25.59601, 
    25.62336, 25.65055, 25.6776, 25.70449, 25.73122, 25.75781, 25.78424, 
    25.81051, 25.83663, 25.8626, 25.88841, 25.91407, 25.93958, 25.96493, 
    25.99012, 26.01516, 26.04005, 26.06477, 26.08935, 26.11376, 26.13802, 
    26.16213, 26.18608, 26.20987, 26.2335, 26.25698, 26.28029, 26.30346, 
    26.32646, 26.34931, 26.372, 26.39453, 26.4169, 26.43911, 26.46117, 
    26.48306, 26.5048, 26.52638, 26.5478, 26.56906, 26.59016, 26.6111, 
    26.63188, 26.6525, 26.67296, 26.69326, 26.71339, 26.73337, 26.75319, 
    26.77284, 26.79234, 26.81167, 26.83084, 26.84985, 26.8687, 26.88739, 
    26.90591, 26.92427, 26.94247, 26.96051, 26.97838, 26.9961, 27.01364, 
    27.03103, 27.04825, 27.06531, 27.0822, 27.09893, 27.1155, 27.1319, 
    27.14815, 27.16422, 27.18013, 27.19588, 27.21146, 27.22688, 27.24213, 
    27.25722, 27.27214, 27.2869, 27.30149, 27.31591, 27.33017, 27.34427, 
    27.3582, 27.37196, 27.38556, 27.39899, 27.41226, 27.42535, 27.43829, 
    27.45105, 27.46365, 27.47608, 27.48835, 27.50045, 27.51238, 27.52414, 
    27.53574, 27.54717, 27.55843, 27.56953, 27.58045, 27.59122, 27.60181, 
    27.61223, 27.62249, 27.63257, 27.64249, 27.65224, 27.66183, 27.67124, 
    27.68049, 27.68957, 27.69847, 27.70721, 27.71579, 27.72419, 27.73242, 
    27.74049, 27.74838, 27.75611, 27.76367, 27.77106, 27.77828, 27.78533, 
    27.79221, 27.79892, 27.80546, 27.81183, 27.81803, 27.82406, 27.82993, 
    27.83562, 27.84114, 27.8465, 27.85168, 27.85669, 27.86154, 27.86621, 
    27.87071, 27.87505, 27.87921, 27.8832, 27.88702, 27.89068, 27.89416, 
    27.89747, 27.90061, 27.90358, 27.90638, 27.90901, 27.91147, 27.91376, 
    27.91588, 27.91783, 27.91961, 27.92121, 27.92265, 27.92391, 27.92501, 
    27.92593, 27.92669, 27.92727, 27.92768, 27.92793, 27.928, 27.9279, 
    27.92763, 27.92719, 27.92658, 27.9258, 27.92485, 27.92373, 27.92243, 
    27.92097, 27.91933, 27.91753, 27.91556, 27.91341, 27.91109, 27.90861, 
    27.90595, 27.90312, 27.90013, 27.89696, 27.89362, 27.89011, 27.88643, 
    27.88258, 27.87856, 27.87437, 27.87001, 27.86548, 27.86078, 27.85591, 
    27.85087, 27.84566, 27.84028, 27.83473, 27.82901, 27.82312, 27.81706, 
    27.81083, 27.80443, 27.79787, 27.79113, 27.78422, 27.77715, 27.7699, 
    27.76248, 27.7549, 27.74715, 27.73922, 27.73113, 27.72287, 27.71444, 
    27.70584, 27.69708, 27.68814, 27.67904, 27.66976, 27.66032, 27.65071, 
    27.64093, 27.63099, 27.62087, 27.61059, 27.60014, 27.58952, 27.57874, 
    27.56778, 27.55666, 27.54537, 27.53392, 27.52229, 27.5105, 27.49854, 
    27.48642, 27.47413, 27.46167, 27.44905, 27.43625, 27.42329, 27.41017, 
    27.39688, 27.38342, 27.3698, 27.35601, 27.34205, 27.32793, 27.31364, 
    27.29919, 27.28457, 27.26979, 27.25484, 27.23973, 27.22445, 27.20901, 
    27.1934, 27.17763, 27.16169, 27.14559, 27.12932, 27.11289, 27.0963, 
    27.07954, 27.06262, 27.04554, 27.02829, 27.01088, 26.99331, 26.97557, 
    26.95767, 26.93961, 26.92138, 26.90299, 26.88444, 26.86573, 26.84686, 
    26.82782, 26.80862, 26.78927, 26.76975, 26.75006, 26.73022, 26.71022, 
    26.69006, 26.66973, 26.64925, 26.6286, 26.6078, 26.58683, 26.56571, 
    26.54442, 26.52298, 26.50137, 26.47961, 26.45769, 26.43561, 26.41337, 
    26.39097, 26.36842, 26.34571, 26.32283, 26.2998, 26.27662, 26.25327, 
    26.22977, 26.20611, 26.1823, 26.15833, 26.1342, 26.10991, 26.08547, 
    26.06087, 26.03612, 26.01121, 25.98615, 25.96093, 25.93555, 25.91003, 
    25.88434, 25.8585, 25.83251, 25.80637, 25.78007, 25.75361, 25.72701, 
    25.70024, 25.67333, 25.64626, 25.61904, 25.59167, 25.56415, 25.53647, 
    25.50864, 25.48066,
  22.35246, 22.39362, 22.43466, 22.47556, 22.51634, 22.55698, 22.59749, 
    22.63787, 22.67811, 22.71822, 22.75821, 22.79805, 22.83777, 22.87735, 
    22.9168, 22.95611, 22.99529, 23.03434, 23.07325, 23.11202, 23.15066, 
    23.18917, 23.22754, 23.26577, 23.30387, 23.34184, 23.37966, 23.41735, 
    23.4549, 23.49232, 23.52959, 23.56673, 23.60373, 23.6406, 23.67732, 
    23.71391, 23.75036, 23.78666, 23.82283, 23.85886, 23.89475, 23.9305, 
    23.96611, 24.00158, 24.03691, 24.07209, 24.10714, 24.14204, 24.17681, 
    24.21143, 24.24591, 24.28024, 24.31444, 24.34849, 24.38239, 24.41616, 
    24.44978, 24.48326, 24.51659, 24.54978, 24.58282, 24.61572, 24.64848, 
    24.68108, 24.71355, 24.74587, 24.77804, 24.81007, 24.84195, 24.87368, 
    24.90527, 24.93671, 24.968, 24.99915, 25.03015, 25.061, 25.0917, 
    25.12226, 25.15266, 25.18292, 25.21303, 25.24299, 25.2728, 25.30246, 
    25.33197, 25.36134, 25.39055, 25.41961, 25.44852, 25.47728, 25.50589, 
    25.53435, 25.56265, 25.59081, 25.61881, 25.64666, 25.67436, 25.70191, 
    25.7293, 25.75654, 25.78363, 25.81057, 25.83735, 25.86398, 25.89045, 
    25.91677, 25.94294, 25.96895, 25.99481, 26.02051, 26.04606, 26.07145, 
    26.09669, 26.12177, 26.1467, 26.17147, 26.19608, 26.22054, 26.24485, 
    26.26899, 26.29298, 26.31681, 26.34049, 26.364, 26.38736, 26.41056, 
    26.43361, 26.4565, 26.47922, 26.50179, 26.5242, 26.54646, 26.56855, 
    26.59048, 26.61226, 26.63388, 26.65533, 26.67663, 26.69777, 26.71874, 
    26.73956, 26.76021, 26.78071, 26.80104, 26.82122, 26.84123, 26.86108, 
    26.88077, 26.9003, 26.91967, 26.93888, 26.95792, 26.9768, 26.99552, 
    27.01407, 27.03247, 27.0507, 27.06877, 27.08668, 27.10442, 27.122, 
    27.13941, 27.15667, 27.17375, 27.19068, 27.20744, 27.22404, 27.24047, 
    27.25674, 27.27284, 27.28878, 27.30456, 27.32017, 27.33561, 27.35089, 
    27.366, 27.38095, 27.39574, 27.41035, 27.42481, 27.43909, 27.45321, 
    27.46717, 27.48096, 27.49458, 27.50803, 27.52132, 27.53444, 27.5474, 
    27.56019, 27.57281, 27.58526, 27.59755, 27.60967, 27.62163, 27.63341, 
    27.64503, 27.65648, 27.66776, 27.67888, 27.68982, 27.7006, 27.71121, 
    27.72165, 27.73193, 27.74203, 27.75197, 27.76174, 27.77134, 27.78078, 
    27.79004, 27.79913, 27.80806, 27.81681, 27.8254, 27.83382, 27.84207, 
    27.85015, 27.85806, 27.8658, 27.87337, 27.88077, 27.888, 27.89507, 
    27.90196, 27.90868, 27.91523, 27.92162, 27.92783, 27.93387, 27.93975, 
    27.94545, 27.95098, 27.95635, 27.96154, 27.96656, 27.97141, 27.9761, 
    27.98061, 27.98495, 27.98912, 27.99312, 27.99695, 28.00061, 28.0041, 
    28.00741, 28.01056, 28.01354, 28.01634, 28.01898, 28.02144, 28.02374, 
    28.02586, 28.02781, 28.02959, 28.0312, 28.03264, 28.03391, 28.035, 
    28.03593, 28.03669, 28.03727, 28.03769, 28.03793, 28.038, 28.0379, 
    28.03763, 28.03719, 28.03658, 28.0358, 28.03484, 28.03372, 28.03242, 
    28.03096, 28.02932, 28.02751, 28.02553, 28.02338, 28.02106, 28.01857, 
    28.01591, 28.01308, 28.01007, 28.0069, 28.00356, 28.00004, 27.99636, 
    27.9925, 27.98847, 27.98427, 27.97991, 27.97537, 27.97066, 27.96578, 
    27.96073, 27.95551, 27.95012, 27.94456, 27.93883, 27.93293, 27.92686, 
    27.92062, 27.91421, 27.90763, 27.90088, 27.89396, 27.88687, 27.87961, 
    27.87218, 27.86458, 27.85682, 27.84888, 27.84077, 27.8325, 27.82405, 
    27.81544, 27.80666, 27.7977, 27.78858, 27.77929, 27.76983, 27.76021, 
    27.75041, 27.74045, 27.73032, 27.72001, 27.70955, 27.69891, 27.6881, 
    27.67713, 27.66599, 27.65468, 27.6432, 27.63156, 27.61975, 27.60777, 
    27.59562, 27.58331, 27.57082, 27.55818, 27.54536, 27.53238, 27.51923, 
    27.50591, 27.49243, 27.47878, 27.46497, 27.45099, 27.43684, 27.42253, 
    27.40805, 27.39341, 27.3786, 27.36362, 27.34848, 27.33318, 27.31771, 
    27.30207, 27.28627, 27.27031, 27.25418, 27.23788, 27.22142, 27.2048, 
    27.18801, 27.17106, 27.15395, 27.13667, 27.11923, 27.10162, 27.08385, 
    27.06592, 27.04783, 27.02957, 27.01115, 26.99257, 26.97382, 26.95492, 
    26.93585, 26.91662, 26.89722, 26.87767, 26.85795, 26.83808, 26.81804, 
    26.79784, 26.77748, 26.75696, 26.73628, 26.71544, 26.69443, 26.67327, 
    26.65195, 26.63047, 26.60883, 26.58703, 26.56507, 26.54295, 26.52067, 
    26.49823, 26.47564, 26.45289, 26.42998, 26.40691, 26.38368, 26.36029, 
    26.33675, 26.31305, 26.2892, 26.26518, 26.24101, 26.21668, 26.1922, 
    26.16756, 26.14277, 26.11782, 26.09271, 26.06745, 26.04203, 26.01646, 
    25.99073, 25.96485, 25.93881, 25.91262, 25.88627, 25.85978, 25.83312, 
    25.80632, 25.77936, 25.75224, 25.72498, 25.69756, 25.66999, 25.64227, 
    25.61439, 25.58636,
  22.45296, 22.49419, 22.53529, 22.57625, 22.61709, 22.65779, 22.69836, 
    22.73881, 22.77911, 22.81929, 22.85933, 22.89924, 22.93902, 22.97866, 
    23.01817, 23.05754, 23.09678, 23.13589, 23.17486, 23.2137, 23.2524, 
    23.29097, 23.3294, 23.36769, 23.40585, 23.44387, 23.48176, 23.5195, 
    23.55712, 23.59459, 23.63193, 23.66912, 23.70618, 23.7431, 23.77989, 
    23.81653, 23.85304, 23.8894, 23.92563, 23.96172, 23.99767, 24.03347, 
    24.06914, 24.10466, 24.14005, 24.17529, 24.21039, 24.24535, 24.28017, 
    24.31485, 24.34938, 24.38378, 24.41802, 24.45213, 24.48609, 24.51991, 
    24.55359, 24.58712, 24.6205, 24.65375, 24.68685, 24.7198, 24.75261, 
    24.78527, 24.81779, 24.85016, 24.88239, 24.91446, 24.9464, 24.97819, 
    25.00982, 25.04132, 25.07266, 25.10386, 25.13491, 25.16581, 25.19657, 
    25.22717, 25.25763, 25.28794, 25.3181, 25.34811, 25.37797, 25.40768, 
    25.43724, 25.46665, 25.49591, 25.52502, 25.55398, 25.58279, 25.61144, 
    25.63995, 25.6683, 25.69651, 25.72456, 25.75246, 25.7802, 25.8078, 
    25.83524, 25.86252, 25.88966, 25.91664, 25.94347, 25.97014, 25.99666, 
    26.02303, 26.04924, 26.07529, 26.1012, 26.12694, 26.15253, 26.17797, 
    26.20325, 26.22838, 26.25335, 26.27816, 26.30282, 26.32732, 26.35166, 
    26.37585, 26.39988, 26.42375, 26.44747, 26.47103, 26.49443, 26.51767, 
    26.54075, 26.56368, 26.58645, 26.60905, 26.6315, 26.6538, 26.67593, 
    26.6979, 26.71971, 26.74137, 26.76286, 26.78419, 26.80537, 26.82638, 
    26.84723, 26.86793, 26.88846, 26.90883, 26.92904, 26.94909, 26.96897, 
    26.9887, 27.00826, 27.02766, 27.0469, 27.06598, 27.08489, 27.10365, 
    27.12223, 27.14066, 27.15893, 27.17702, 27.19496, 27.21274, 27.23035, 
    27.2478, 27.26508, 27.2822, 27.29915, 27.31594, 27.33257, 27.34903, 
    27.36533, 27.38146, 27.39743, 27.41323, 27.42887, 27.44434, 27.45965, 
    27.47479, 27.48977, 27.50457, 27.51922, 27.5337, 27.54801, 27.56215, 
    27.57613, 27.58995, 27.60359, 27.61707, 27.63038, 27.64353, 27.65651, 
    27.66932, 27.68196, 27.69444, 27.70675, 27.71889, 27.73087, 27.74268, 
    27.75431, 27.76579, 27.77709, 27.78822, 27.79919, 27.80999, 27.82062, 
    27.83108, 27.84137, 27.8515, 27.86145, 27.87124, 27.88086, 27.89031, 
    27.89959, 27.9087, 27.91764, 27.92641, 27.93501, 27.94345, 27.95171, 
    27.9598, 27.96773, 27.97548, 27.98307, 27.99048, 27.99773, 28.0048, 
    28.01171, 28.01845, 28.02501, 28.0314, 28.03763, 28.04368, 28.04957, 
    28.05528, 28.06083, 28.0662, 28.0714, 28.07643, 28.08129, 28.08598, 
    28.0905, 28.09485, 28.09903, 28.10304, 28.10687, 28.11054, 28.11403, 
    28.11736, 28.12051, 28.12349, 28.1263, 28.12894, 28.13141, 28.13371, 
    28.13583, 28.13779, 28.13957, 28.14119, 28.14263, 28.1439, 28.145, 
    28.14593, 28.14668, 28.14727, 28.14768, 28.14793, 28.148, 28.1479, 
    28.14763, 28.14719, 28.14658, 28.14579, 28.14484, 28.14371, 28.14241, 
    28.14094, 28.1393, 28.13749, 28.13551, 28.13336, 28.13103, 28.12854, 
    28.12587, 28.12303, 28.12002, 28.11684, 28.11349, 28.10997, 28.10628, 
    28.10242, 28.09838, 28.09418, 28.0898, 28.08525, 28.08054, 28.07565, 
    28.07059, 28.06536, 28.05996, 28.05439, 28.04865, 28.04274, 28.03666, 
    28.03041, 28.02398, 28.01739, 28.01063, 28.0037, 27.9966, 27.98932, 
    27.98188, 27.97427, 27.96649, 27.95853, 27.95041, 27.94212, 27.93366, 
    27.92503, 27.91623, 27.90727, 27.89813, 27.88882, 27.87935, 27.8697, 
    27.85989, 27.84991, 27.83976, 27.82944, 27.81895, 27.80829, 27.79747, 
    27.78647, 27.77531, 27.76398, 27.75249, 27.74082, 27.72899, 27.71699, 
    27.70482, 27.69248, 27.67998, 27.6673, 27.65447, 27.64146, 27.62829, 
    27.61495, 27.60144, 27.58777, 27.57393, 27.55993, 27.54576, 27.53142, 
    27.51691, 27.50224, 27.48741, 27.4724, 27.45724, 27.4419, 27.4264, 
    27.41074, 27.39491, 27.37892, 27.36276, 27.34644, 27.32995, 27.3133, 
    27.29648, 27.2795, 27.26235, 27.24504, 27.22757, 27.20994, 27.19214, 
    27.17417, 27.15605, 27.13776, 27.1193, 27.10069, 27.08191, 27.06297, 
    27.04387, 27.0246, 27.00518, 26.98559, 26.96584, 26.94592, 26.92585, 
    26.90562, 26.88522, 26.86466, 26.84395, 26.82307, 26.80203, 26.78083, 
    26.75947, 26.73795, 26.71627, 26.69444, 26.67244, 26.65028, 26.62796, 
    26.60549, 26.58286, 26.56006, 26.53711, 26.514, 26.49073, 26.46731, 
    26.44373, 26.41999, 26.39609, 26.37203, 26.34782, 26.32345, 26.29893, 
    26.27425, 26.24941, 26.22441, 26.19926, 26.17396, 26.1485, 26.12288, 
    26.09711, 26.07118, 26.0451, 26.01887, 25.99248, 25.96593, 25.93923, 
    25.91238, 25.88538, 25.85822, 25.83091, 25.80344, 25.77582, 25.74805, 
    25.72013, 25.69206,
  22.55345, 22.59474, 22.6359, 22.67693, 22.71783, 22.75859, 22.79923, 
    22.83973, 22.8801, 22.92034, 22.96044, 23.00041, 23.04025, 23.07995, 
    23.11953, 23.15896, 23.19826, 23.23743, 23.27646, 23.31536, 23.35412, 
    23.39275, 23.43124, 23.46959, 23.50781, 23.54589, 23.58384, 23.62164, 
    23.65932, 23.69685, 23.73424, 23.7715, 23.80862, 23.8456, 23.88244, 
    23.91915, 23.95571, 23.99213, 24.02842, 24.06456, 24.10057, 24.13643, 
    24.17215, 24.20774, 24.24318, 24.27848, 24.31364, 24.34865, 24.38353, 
    24.41826, 24.45285, 24.4873, 24.5216, 24.55576, 24.58978, 24.62366, 
    24.65738, 24.69097, 24.72441, 24.75771, 24.79086, 24.82387, 24.85673, 
    24.88945, 24.92202, 24.95444, 24.98672, 25.01885, 25.05084, 25.08268, 
    25.11437, 25.14592, 25.17731, 25.20856, 25.23966, 25.27062, 25.30142, 
    25.33208, 25.36259, 25.39294, 25.42315, 25.45321, 25.48313, 25.51289, 
    25.5425, 25.57196, 25.60126, 25.63042, 25.65943, 25.68829, 25.71699, 
    25.74555, 25.77395, 25.8022, 25.8303, 25.85824, 25.88604, 25.91368, 
    25.94116, 25.9685, 25.99568, 26.02271, 26.04958, 26.0763, 26.10286, 
    26.12927, 26.15553, 26.18163, 26.20758, 26.23337, 26.259, 26.28448, 
    26.30981, 26.33498, 26.35999, 26.38484, 26.40954, 26.43409, 26.45847, 
    26.4827, 26.50677, 26.53069, 26.55444, 26.57804, 26.60148, 26.62477, 
    26.64789, 26.67086, 26.69366, 26.71631, 26.7388, 26.76113, 26.7833, 
    26.80531, 26.82716, 26.84885, 26.87039, 26.89176, 26.91297, 26.93402, 
    26.95491, 26.97564, 26.9962, 27.01661, 27.03685, 27.05694, 27.07686, 
    27.09662, 27.11621, 27.13565, 27.15492, 27.17403, 27.19298, 27.21177, 
    27.23039, 27.24885, 27.26715, 27.28528, 27.30325, 27.32105, 27.3387, 
    27.35617, 27.37349, 27.39064, 27.40762, 27.42444, 27.4411, 27.45759, 
    27.47392, 27.49008, 27.50607, 27.5219, 27.53757, 27.55307, 27.5684, 
    27.58357, 27.59857, 27.61341, 27.62808, 27.64258, 27.65692, 27.67109, 
    27.6851, 27.69893, 27.71261, 27.72611, 27.73945, 27.75261, 27.76562, 
    27.77845, 27.79112, 27.80362, 27.81595, 27.82812, 27.84011, 27.85194, 
    27.8636, 27.87509, 27.88642, 27.89757, 27.90856, 27.91937, 27.93002, 
    27.9405, 27.95082, 27.96096, 27.97093, 27.98074, 27.99037, 27.99984, 
    28.00913, 28.01826, 28.02722, 28.03601, 28.04462, 28.05307, 28.06135, 
    28.06946, 28.0774, 28.08517, 28.09277, 28.1002, 28.10745, 28.11454, 
    28.12146, 28.12821, 28.13479, 28.14119, 28.14743, 28.15349, 28.15939, 
    28.16511, 28.17067, 28.17605, 28.18126, 28.1863, 28.19117, 28.19587, 
    28.2004, 28.20475, 28.20894, 28.21296, 28.2168, 28.22047, 28.22397, 
    28.2273, 28.23046, 28.23345, 28.23626, 28.23891, 28.24138, 28.24368, 
    28.24581, 28.24777, 28.24956, 28.25117, 28.25262, 28.25389, 28.25499, 
    28.25592, 28.25668, 28.25727, 28.25768, 28.25793, 28.258, 28.2579, 
    28.25763, 28.25719, 28.25657, 28.25579, 28.25483, 28.2537, 28.2524, 
    28.25093, 28.24929, 28.24747, 28.24549, 28.24333, 28.241, 28.2385, 
    28.23583, 28.23299, 28.22997, 28.22679, 28.22343, 28.2199, 28.2162, 
    28.21233, 28.20829, 28.20408, 28.19969, 28.19514, 28.19041, 28.18551, 
    28.18045, 28.17521, 28.1698, 28.16422, 28.15847, 28.15255, 28.14645, 
    28.14019, 28.13376, 28.12715, 28.12038, 28.11343, 28.10632, 28.09903, 
    28.09158, 28.08395, 28.07615, 28.06819, 28.06005, 28.05175, 28.04327, 
    28.03463, 28.02581, 28.01683, 28.00768, 27.99835, 27.98886, 27.9792, 
    27.96937, 27.95936, 27.9492, 27.93886, 27.92835, 27.91768, 27.90683, 
    27.89582, 27.88464, 27.87329, 27.86177, 27.85008, 27.83822, 27.8262, 
    27.81401, 27.80165, 27.78913, 27.77643, 27.76357, 27.75054, 27.73735, 
    27.72398, 27.71045, 27.69676, 27.68289, 27.66886, 27.65466, 27.6403, 
    27.62577, 27.61107, 27.59621, 27.58118, 27.56599, 27.55063, 27.5351, 
    27.51941, 27.50355, 27.48753, 27.47134, 27.45499, 27.43847, 27.42179, 
    27.40495, 27.38793, 27.37076, 27.35342, 27.33591, 27.31825, 27.30042, 
    27.28242, 27.26426, 27.24594, 27.22746, 27.20881, 27.19, 27.17102, 
    27.15189, 27.13259, 27.11313, 27.0935, 27.07372, 27.05377, 27.03366, 
    27.01339, 26.99296, 26.97237, 26.95161, 26.9307, 26.90962, 26.88839, 
    26.86699, 26.84543, 26.82372, 26.80184, 26.7798, 26.75761, 26.73525, 
    26.71274, 26.69007, 26.66723, 26.64424, 26.62109, 26.59779, 26.57432, 
    26.5507, 26.52691, 26.50298, 26.47888, 26.45463, 26.43022, 26.40565, 
    26.38092, 26.35604, 26.33101, 26.30581, 26.28046, 26.25496, 26.2293, 
    26.20348, 26.17751, 26.15139, 26.12511, 26.09867, 26.07208, 26.04534, 
    26.01844, 25.99139, 25.96418, 25.93683, 25.90932, 25.88165, 25.85383, 
    25.82586, 25.79774,
  22.65392, 22.69528, 22.7365, 22.77759, 22.81855, 22.85938, 22.90008, 
    22.94064, 22.98108, 23.02137, 23.06154, 23.10157, 23.14147, 23.18124, 
    23.22087, 23.26037, 23.29973, 23.33896, 23.37805, 23.41701, 23.45583, 
    23.49452, 23.53307, 23.57148, 23.60976, 23.6479, 23.68591, 23.72377, 
    23.7615, 23.7991, 23.83655, 23.87387, 23.91105, 23.94808, 23.98498, 
    24.02174, 24.05837, 24.09485, 24.13119, 24.16739, 24.20345, 24.23938, 
    24.27516, 24.3108, 24.34629, 24.38165, 24.41687, 24.45194, 24.48687, 
    24.52166, 24.5563, 24.59081, 24.62517, 24.65939, 24.69346, 24.72739, 
    24.76117, 24.79481, 24.82831, 24.86166, 24.89487, 24.92793, 24.96084, 
    24.99361, 25.02624, 25.05872, 25.09105, 25.12323, 25.15527, 25.18716, 
    25.21891, 25.2505, 25.28195, 25.31326, 25.34441, 25.37541, 25.40627, 
    25.43698, 25.46754, 25.49794, 25.5282, 25.55831, 25.58827, 25.61808, 
    25.64774, 25.67725, 25.70661, 25.73582, 25.76488, 25.79378, 25.82254, 
    25.85114, 25.87959, 25.90788, 25.93603, 25.96402, 25.99186, 26.01955, 
    26.04708, 26.07446, 26.10169, 26.12876, 26.15568, 26.18245, 26.20906, 
    26.23551, 26.26181, 26.28796, 26.31395, 26.33979, 26.36547, 26.39099, 
    26.41636, 26.44157, 26.46662, 26.49152, 26.51626, 26.54085, 26.56528, 
    26.58955, 26.61366, 26.63762, 26.66141, 26.68505, 26.70853, 26.73186, 
    26.75502, 26.77803, 26.80087, 26.82356, 26.84609, 26.86846, 26.89067, 
    26.91272, 26.93461, 26.95634, 26.97791, 26.99931, 27.02056, 27.04165, 
    27.06257, 27.08334, 27.10394, 27.12438, 27.14466, 27.16478, 27.18474, 
    27.20453, 27.22417, 27.24364, 27.26294, 27.28209, 27.30107, 27.31989, 
    27.33854, 27.35703, 27.37536, 27.39353, 27.41153, 27.42937, 27.44704, 
    27.46455, 27.48189, 27.49907, 27.51609, 27.53294, 27.54962, 27.56614, 
    27.5825, 27.59869, 27.61471, 27.63057, 27.64627, 27.66179, 27.67716, 
    27.69235, 27.70738, 27.72224, 27.73694, 27.75147, 27.76583, 27.78003, 
    27.79406, 27.80792, 27.82162, 27.83515, 27.84851, 27.8617, 27.87473, 
    27.88758, 27.90027, 27.91279, 27.92515, 27.93734, 27.94935, 27.9612, 
    27.97288, 27.9844, 27.99574, 28.00691, 28.01792, 28.02876, 28.03943, 
    28.04993, 28.06026, 28.07042, 28.08041, 28.09023, 28.09988, 28.10937, 
    28.11868, 28.12782, 28.1368, 28.1456, 28.15424, 28.1627, 28.17099, 
    28.17912, 28.18707, 28.19485, 28.20247, 28.20991, 28.21718, 28.22428, 
    28.23121, 28.23797, 28.24456, 28.25098, 28.25723, 28.2633, 28.26921, 
    28.27494, 28.28051, 28.2859, 28.29112, 28.29617, 28.30105, 28.30576, 
    28.31029, 28.31466, 28.31885, 28.32287, 28.32672, 28.3304, 28.33391, 
    28.33725, 28.34041, 28.3434, 28.34622, 28.34887, 28.35135, 28.35366, 
    28.35579, 28.35775, 28.35954, 28.36116, 28.36261, 28.36388, 28.36499, 
    28.36592, 28.36668, 28.36727, 28.36768, 28.36793, 28.368, 28.3679, 
    28.36763, 28.36719, 28.36657, 28.36578, 28.36482, 28.36369, 28.36239, 
    28.36092, 28.35927, 28.35745, 28.35546, 28.3533, 28.35097, 28.34846, 
    28.34579, 28.34294, 28.33992, 28.33673, 28.33337, 28.32983, 28.32613, 
    28.32225, 28.3182, 28.31398, 28.30959, 28.30502, 28.30029, 28.29538, 
    28.29031, 28.28506, 28.27964, 28.27405, 28.26829, 28.26235, 28.25625, 
    28.24998, 28.24353, 28.23691, 28.23013, 28.22317, 28.21604, 28.20874, 
    28.20127, 28.19363, 28.18582, 28.17784, 28.16969, 28.16137, 28.15288, 
    28.14422, 28.13539, 28.12639, 28.11722, 28.10788, 28.09837, 28.08869, 
    28.07884, 28.06882, 28.05863, 28.04828, 28.03775, 28.02706, 28.01619, 
    28.00516, 27.99396, 27.98259, 27.97105, 27.95934, 27.94746, 27.93542, 
    27.92321, 27.91083, 27.89828, 27.88556, 27.87267, 27.85962, 27.8464, 
    27.83302, 27.81946, 27.80574, 27.79185, 27.7778, 27.76357, 27.74918, 
    27.73463, 27.7199, 27.70502, 27.68996, 27.67474, 27.65935, 27.6438, 
    27.62808, 27.61219, 27.59614, 27.57992, 27.56354, 27.547, 27.53028, 
    27.51341, 27.49637, 27.47916, 27.46179, 27.44425, 27.42656, 27.40869, 
    27.39067, 27.37247, 27.35412, 27.3356, 27.31692, 27.29808, 27.27907, 
    27.2599, 27.24057, 27.22107, 27.20141, 27.18159, 27.16161, 27.14147, 
    27.12116, 27.10069, 27.08006, 27.05927, 27.03832, 27.01721, 26.99594, 
    26.9745, 26.95291, 26.93115, 26.90924, 26.88717, 26.86493, 26.84254, 
    26.81998, 26.79727, 26.7744, 26.75137, 26.72818, 26.70483, 26.68132, 
    26.65766, 26.63384, 26.60986, 26.58572, 26.56142, 26.53697, 26.51236, 
    26.48759, 26.46267, 26.43759, 26.41235, 26.38696, 26.36141, 26.33571, 
    26.30985, 26.28383, 26.25766, 26.23134, 26.20486, 26.17822, 26.15144, 
    26.12449, 26.09739, 26.07014, 26.04274, 26.01518, 25.98747, 25.95961, 
    25.93159, 25.90342,
  22.75438, 22.7958, 22.83709, 22.87824, 22.91926, 22.96015, 23.00091, 
    23.04154, 23.08204, 23.12239, 23.16262, 23.20272, 23.24268, 23.28251, 
    23.3222, 23.36176, 23.40118, 23.44047, 23.47963, 23.51864, 23.55753, 
    23.59627, 23.63489, 23.67336, 23.7117, 23.7499, 23.78796, 23.82589, 
    23.86368, 23.90133, 23.93884, 23.97622, 24.01346, 24.05055, 24.08751, 
    24.12433, 24.16101, 24.19755, 24.23395, 24.27021, 24.30633, 24.34231, 
    24.37815, 24.41385, 24.4494, 24.48482, 24.52009, 24.55522, 24.5902, 
    24.62505, 24.65975, 24.69431, 24.72872, 24.763, 24.79712, 24.83111, 
    24.86495, 24.89864, 24.9322, 24.9656, 24.99886, 25.03198, 25.06495, 
    25.09777, 25.13045, 25.16298, 25.19536, 25.2276, 25.25969, 25.29164, 
    25.32343, 25.35508, 25.38659, 25.41794, 25.44914, 25.4802, 25.51111, 
    25.54186, 25.57247, 25.60293, 25.63324, 25.6634, 25.69341, 25.72327, 
    25.75298, 25.78254, 25.81195, 25.84121, 25.87031, 25.89927, 25.92807, 
    25.95672, 25.98522, 26.01356, 26.04176, 26.0698, 26.09768, 26.12542, 
    26.153, 26.18042, 26.2077, 26.23482, 26.26178, 26.28859, 26.31524, 
    26.34175, 26.36809, 26.39428, 26.42032, 26.4462, 26.47192, 26.49749, 
    26.5229, 26.54815, 26.57325, 26.59819, 26.62298, 26.64761, 26.67208, 
    26.69639, 26.72054, 26.74454, 26.76838, 26.79206, 26.81558, 26.83894, 
    26.86215, 26.88519, 26.90808, 26.93081, 26.95337, 26.97578, 26.99803, 
    27.02012, 27.04205, 27.06381, 27.08542, 27.10686, 27.12815, 27.14927, 
    27.17024, 27.19104, 27.21168, 27.23215, 27.25247, 27.27262, 27.29262, 
    27.31245, 27.33211, 27.35162, 27.37096, 27.39014, 27.40915, 27.428, 
    27.44669, 27.46522, 27.48358, 27.50177, 27.51981, 27.53768, 27.55538, 
    27.57292, 27.5903, 27.60751, 27.62455, 27.64143, 27.65815, 27.6747, 
    27.69108, 27.7073, 27.72335, 27.73924, 27.75496, 27.77052, 27.78591, 
    27.80113, 27.81618, 27.83108, 27.8458, 27.86035, 27.87474, 27.88897, 
    27.90302, 27.91691, 27.93063, 27.94418, 27.95756, 27.97078, 27.98383, 
    27.99671, 28.00942, 28.02197, 28.03435, 28.04655, 28.05859, 28.07046, 
    28.08216, 28.0937, 28.10506, 28.11626, 28.12729, 28.13814, 28.14883, 
    28.15935, 28.1697, 28.17988, 28.18989, 28.19973, 28.2094, 28.2189, 
    28.22823, 28.23739, 28.24638, 28.2552, 28.26385, 28.27233, 28.28063, 
    28.28877, 28.29674, 28.30454, 28.31216, 28.31962, 28.32691, 28.33402, 
    28.34096, 28.34773, 28.35434, 28.36077, 28.36703, 28.37311, 28.37903, 
    28.38477, 28.39035, 28.39575, 28.40098, 28.40604, 28.41093, 28.41564, 
    28.42019, 28.42456, 28.42876, 28.43279, 28.43665, 28.44033, 28.44385, 
    28.44719, 28.45036, 28.45336, 28.45618, 28.45884, 28.46132, 28.46363, 
    28.46577, 28.46773, 28.46953, 28.47115, 28.4726, 28.47388, 28.47498, 
    28.47592, 28.47668, 28.47727, 28.47768, 28.47793, 28.478, 28.4779, 
    28.47763, 28.47718, 28.47657, 28.47578, 28.47482, 28.47369, 28.47238, 
    28.47091, 28.46926, 28.46743, 28.46544, 28.46328, 28.46094, 28.45843, 
    28.45575, 28.45289, 28.44987, 28.44667, 28.4433, 28.43976, 28.43605, 
    28.43217, 28.42811, 28.42388, 28.41948, 28.41491, 28.41017, 28.40525, 
    28.40016, 28.39491, 28.38948, 28.38388, 28.3781, 28.37216, 28.36605, 
    28.35976, 28.3533, 28.34668, 28.33988, 28.3329, 28.32576, 28.31845, 
    28.31097, 28.30332, 28.29549, 28.2875, 28.27933, 28.271, 28.26249, 
    28.25381, 28.24497, 28.23595, 28.22676, 28.21741, 28.20788, 28.19818, 
    28.18831, 28.17828, 28.16807, 28.1577, 28.14715, 28.13643, 28.12555, 
    28.1145, 28.10328, 28.09188, 28.08033, 28.0686, 28.0567, 28.04463, 
    28.0324, 28.01999, 28.00742, 27.99468, 27.98178, 27.9687, 27.95546, 
    27.94205, 27.92847, 27.91472, 27.90081, 27.88673, 27.87248, 27.85806, 
    27.84348, 27.82873, 27.81382, 27.79873, 27.78348, 27.76807, 27.75249, 
    27.73674, 27.72083, 27.70475, 27.6885, 27.67209, 27.65551, 27.63877, 
    27.62187, 27.60479, 27.58756, 27.57016, 27.55259, 27.53486, 27.51697, 
    27.49891, 27.48068, 27.4623, 27.44375, 27.42503, 27.40615, 27.38711, 
    27.36791, 27.34854, 27.32901, 27.30932, 27.28946, 27.26945, 27.24927, 
    27.22893, 27.20842, 27.18776, 27.16693, 27.14594, 27.12479, 27.10348, 
    27.08201, 27.06038, 27.03859, 27.01664, 26.99452, 26.97225, 26.94982, 
    26.92722, 26.90447, 26.88156, 26.85849, 26.83526, 26.81187, 26.78832, 
    26.76462, 26.74076, 26.71673, 26.69255, 26.66821, 26.64372, 26.61907, 
    26.59426, 26.56929, 26.54417, 26.51889, 26.49345, 26.46786, 26.44211, 
    26.41621, 26.39015, 26.36394, 26.33756, 26.31104, 26.28436, 26.25752, 
    26.23054, 26.20339, 26.1761, 26.14864, 26.12104, 26.09328, 26.06537, 
    26.03731, 26.00909,
  22.85483, 22.89631, 22.93765, 22.97887, 23.01996, 23.06091, 23.10173, 
    23.14242, 23.18298, 23.2234, 23.26369, 23.30385, 23.34387, 23.38376, 
    23.42352, 23.46313, 23.50262, 23.54197, 23.58119, 23.62027, 23.65921, 
    23.69802, 23.73669, 23.77522, 23.81362, 23.85188, 23.89001, 23.92799, 
    23.96584, 24.00355, 24.04113, 24.07856, 24.11585, 24.15301, 24.19003, 
    24.22691, 24.26365, 24.30024, 24.3367, 24.37302, 24.4092, 24.44523, 
    24.48113, 24.51688, 24.5525, 24.58797, 24.62329, 24.65848, 24.69352, 
    24.72843, 24.76318, 24.7978, 24.83227, 24.8666, 24.90078, 24.93482, 
    24.96871, 25.00246, 25.03607, 25.06953, 25.10285, 25.13601, 25.16904, 
    25.20192, 25.23465, 25.26723, 25.29967, 25.33196, 25.36411, 25.3961, 
    25.42795, 25.45965, 25.49121, 25.52261, 25.55387, 25.58497, 25.61593, 
    25.64674, 25.6774, 25.70791, 25.73828, 25.76849, 25.79855, 25.82845, 
    25.85822, 25.88782, 25.91728, 25.94659, 25.97574, 26.00474, 26.03359, 
    26.06229, 26.09084, 26.11923, 26.14747, 26.17556, 26.20349, 26.23127, 
    26.2589, 26.28638, 26.31369, 26.34086, 26.36787, 26.39473, 26.42143, 
    26.44797, 26.47436, 26.5006, 26.52668, 26.5526, 26.57837, 26.60398, 
    26.62943, 26.65473, 26.67987, 26.70486, 26.72969, 26.75436, 26.77887, 
    26.80322, 26.82742, 26.85146, 26.87534, 26.89906, 26.92262, 26.94603, 
    26.96927, 26.99236, 27.01528, 27.03805, 27.06066, 27.0831, 27.10539, 
    27.12751, 27.14948, 27.17129, 27.19293, 27.21441, 27.23573, 27.2569, 
    27.27789, 27.29873, 27.31941, 27.33992, 27.36027, 27.38046, 27.40049, 
    27.42035, 27.44006, 27.45959, 27.47897, 27.49818, 27.51723, 27.53612, 
    27.55484, 27.57339, 27.59179, 27.61002, 27.62808, 27.64598, 27.66372, 
    27.68129, 27.69869, 27.71593, 27.73301, 27.74992, 27.76667, 27.78325, 
    27.79966, 27.81591, 27.83199, 27.84791, 27.86366, 27.87924, 27.89466, 
    27.9099, 27.92499, 27.93991, 27.95465, 27.96924, 27.98365, 27.9979, 
    28.01198, 28.02589, 28.03963, 28.05321, 28.06662, 28.07986, 28.09293, 
    28.10584, 28.11857, 28.13114, 28.14354, 28.15577, 28.16783, 28.17972, 
    28.19145, 28.203, 28.21438, 28.2256, 28.23665, 28.24752, 28.25823, 
    28.26877, 28.27913, 28.28933, 28.29936, 28.30922, 28.31891, 28.32842, 
    28.33777, 28.34695, 28.35596, 28.36479, 28.37346, 28.38195, 28.39027, 
    28.39843, 28.40641, 28.41422, 28.42186, 28.42933, 28.43663, 28.44376, 
    28.45071, 28.4575, 28.46411, 28.47055, 28.47682, 28.48292, 28.48885, 
    28.4946, 28.50019, 28.5056, 28.51084, 28.51591, 28.5208, 28.52553, 
    28.53008, 28.53446, 28.53867, 28.54271, 28.54657, 28.55026, 28.55379, 
    28.55713, 28.56031, 28.56331, 28.56614, 28.5688, 28.57129, 28.5736, 
    28.57574, 28.57771, 28.57951, 28.58114, 28.58259, 28.58387, 28.58498, 
    28.58591, 28.58667, 28.58727, 28.58768, 28.58793, 28.588, 28.5879, 
    28.58763, 28.58718, 28.58657, 28.58578, 28.58481, 28.58368, 28.58237, 
    28.58089, 28.57924, 28.57742, 28.57542, 28.57325, 28.57091, 28.56839, 
    28.56571, 28.56285, 28.55982, 28.55661, 28.55324, 28.54969, 28.54597, 
    28.54208, 28.53802, 28.53378, 28.52937, 28.52479, 28.52004, 28.51512, 
    28.51002, 28.50476, 28.49932, 28.4937, 28.48792, 28.48197, 28.47584, 
    28.46954, 28.46308, 28.45643, 28.44962, 28.44264, 28.43549, 28.42816, 
    28.42067, 28.413, 28.40516, 28.39715, 28.38897, 28.38062, 28.3721, 
    28.3634, 28.35454, 28.34551, 28.3363, 28.32693, 28.31738, 28.30767, 
    28.29779, 28.28773, 28.27751, 28.26711, 28.25655, 28.24581, 28.23491, 
    28.22384, 28.21259, 28.20118, 28.1896, 28.17785, 28.16593, 28.15384, 
    28.14159, 28.12916, 28.11657, 28.10381, 28.09088, 28.07778, 28.06451, 
    28.05107, 28.03747, 28.0237, 28.00976, 27.99566, 27.98138, 27.96694, 
    27.95233, 27.93756, 27.92261, 27.9075, 27.89223, 27.87679, 27.86118, 
    27.8454, 27.82946, 27.81335, 27.79708, 27.78064, 27.76403, 27.74726, 
    27.73032, 27.71322, 27.69595, 27.67852, 27.66092, 27.64316, 27.62523, 
    27.60714, 27.58889, 27.57047, 27.55189, 27.53314, 27.51423, 27.49515, 
    27.47592, 27.45651, 27.43695, 27.41722, 27.39733, 27.37728, 27.35707, 
    27.33669, 27.31615, 27.29545, 27.27458, 27.25356, 27.23237, 27.21103, 
    27.18952, 27.16785, 27.14602, 27.12403, 27.10187, 27.07956, 27.05709, 
    27.03446, 27.01167, 26.98871, 26.9656, 26.94233, 26.91891, 26.89532, 
    26.87157, 26.84767, 26.8236, 26.79938, 26.775, 26.75046, 26.72577, 
    26.70092, 26.67591, 26.65074, 26.62542, 26.59994, 26.5743, 26.54851, 
    26.52256, 26.49646, 26.4702, 26.44378, 26.41721, 26.39049, 26.36361, 
    26.33657, 26.30938, 26.28204, 26.25454, 26.22689, 26.19909, 26.17113, 
    26.14301, 26.11475,
  22.95526, 22.9968, 23.03821, 23.07949, 23.12064, 23.16166, 23.20254, 
    23.24329, 23.28391, 23.3244, 23.36475, 23.40497, 23.44505, 23.485, 
    23.52482, 23.5645, 23.60405, 23.64346, 23.68273, 23.72187, 23.76088, 
    23.79975, 23.83848, 23.87707, 23.91553, 23.95385, 23.99204, 24.03008, 
    24.06799, 24.10576, 24.14339, 24.18089, 24.21824, 24.25546, 24.29253, 
    24.32947, 24.36627, 24.40292, 24.43944, 24.47581, 24.51205, 24.54815, 
    24.5841, 24.61991, 24.65558, 24.6911, 24.72649, 24.76173, 24.79683, 
    24.83179, 24.86661, 24.90128, 24.9358, 24.97019, 25.00443, 25.03852, 
    25.07247, 25.10627, 25.13993, 25.17345, 25.20682, 25.24004, 25.27312, 
    25.30605, 25.33884, 25.37148, 25.40397, 25.43631, 25.46851, 25.50056, 
    25.53246, 25.56421, 25.59582, 25.62728, 25.65858, 25.68974, 25.72075, 
    25.75161, 25.78232, 25.81289, 25.8433, 25.87356, 25.90367, 25.93363, 
    25.96344, 25.9931, 26.0226, 26.05196, 26.08116, 26.11021, 26.13911, 
    26.16786, 26.19645, 26.22489, 26.25318, 26.28131, 26.3093, 26.33713, 
    26.3648, 26.39232, 26.41968, 26.4469, 26.47395, 26.50085, 26.5276, 
    26.55419, 26.58063, 26.60691, 26.63303, 26.659, 26.68481, 26.71047, 
    26.73596, 26.76131, 26.78649, 26.81152, 26.83639, 26.8611, 26.88565, 
    26.91005, 26.93429, 26.95837, 26.98229, 27.00605, 27.02966, 27.0531, 
    27.07639, 27.09951, 27.12248, 27.14528, 27.16793, 27.19041, 27.21274, 
    27.23491, 27.25691, 27.27875, 27.30043, 27.32195, 27.34332, 27.36451, 
    27.38555, 27.40642, 27.42714, 27.44769, 27.46807, 27.4883, 27.50836, 
    27.52826, 27.54799, 27.56757, 27.58698, 27.60622, 27.62531, 27.64422, 
    27.66298, 27.68157, 27.69999, 27.71826, 27.73635, 27.75428, 27.77205, 
    27.78965, 27.80709, 27.82436, 27.84147, 27.85841, 27.87519, 27.89179, 
    27.90824, 27.92451, 27.94062, 27.95657, 27.97235, 27.98796, 28.0034, 
    28.01868, 28.03379, 28.04873, 28.06351, 28.07812, 28.09256, 28.10683, 
    28.12093, 28.13487, 28.14864, 28.16224, 28.17567, 28.18894, 28.20203, 
    28.21496, 28.22772, 28.24031, 28.25273, 28.26498, 28.27707, 28.28898, 
    28.30072, 28.3123, 28.32371, 28.33494, 28.34601, 28.3569, 28.36763, 
    28.37819, 28.38857, 28.39879, 28.40883, 28.41871, 28.42842, 28.43795, 
    28.44732, 28.45651, 28.46553, 28.47438, 28.48306, 28.49158, 28.49991, 
    28.50808, 28.51608, 28.5239, 28.53156, 28.53904, 28.54635, 28.55349, 
    28.56046, 28.56726, 28.57388, 28.58034, 28.58662, 28.59273, 28.59867, 
    28.60443, 28.61003, 28.61545, 28.6207, 28.62578, 28.63068, 28.63541, 
    28.63998, 28.64437, 28.64858, 28.65262, 28.6565, 28.6602, 28.66372, 
    28.66708, 28.67026, 28.67327, 28.6761, 28.67877, 28.68126, 28.68358, 
    28.68572, 28.6877, 28.6895, 28.69112, 28.69258, 28.69386, 28.69497, 
    28.69591, 28.69667, 28.69726, 28.69768, 28.69793, 28.698, 28.6979, 
    28.69763, 28.69718, 28.69656, 28.69577, 28.69481, 28.69367, 28.69236, 
    28.69088, 28.68922, 28.6874, 28.68539, 28.68322, 28.68088, 28.67836, 
    28.67567, 28.6728, 28.66977, 28.66656, 28.66318, 28.65962, 28.6559, 
    28.652, 28.64792, 28.64368, 28.63927, 28.63468, 28.62992, 28.62498, 
    28.61988, 28.6146, 28.60915, 28.60353, 28.59774, 28.59177, 28.58564, 
    28.57933, 28.57285, 28.56619, 28.55937, 28.55238, 28.54521, 28.53787, 
    28.53036, 28.52268, 28.51483, 28.5068, 28.49861, 28.49024, 28.4817, 
    28.47299, 28.46412, 28.45507, 28.44584, 28.43645, 28.42689, 28.41716, 
    28.40726, 28.39718, 28.38694, 28.37653, 28.36594, 28.35519, 28.34427, 
    28.33318, 28.32191, 28.31048, 28.29888, 28.28711, 28.27517, 28.26306, 
    28.25078, 28.23833, 28.22571, 28.21293, 28.19997, 28.18685, 28.17356, 
    28.1601, 28.14647, 28.13268, 28.11871, 28.10458, 28.09028, 28.07582, 
    28.06118, 28.04638, 28.03141, 28.01627, 28.00097, 27.9855, 27.96986, 
    27.95406, 27.93809, 27.92195, 27.90565, 27.88918, 27.87254, 27.85574, 
    27.83877, 27.82164, 27.80434, 27.78688, 27.76925, 27.75146, 27.7335, 
    27.71538, 27.69709, 27.67864, 27.66002, 27.64124, 27.6223, 27.60319, 
    27.58392, 27.56448, 27.54488, 27.52512, 27.5052, 27.48511, 27.46486, 
    27.44444, 27.42387, 27.40313, 27.38223, 27.36117, 27.33995, 27.31856, 
    27.29702, 27.27531, 27.25344, 27.23141, 27.20922, 27.18687, 27.16436, 
    27.14169, 27.11885, 27.09586, 27.07271, 27.0494, 27.02593, 27.0023, 
    26.97852, 26.95457, 26.93047, 26.9062, 26.88178, 26.8572, 26.83246, 
    26.80757, 26.78252, 26.75731, 26.73194, 26.70642, 26.68074, 26.6549, 
    26.62891, 26.60276, 26.57646, 26.55, 26.52338, 26.49661, 26.46968, 
    26.4426, 26.41537, 26.38798, 26.36043, 26.33273, 26.30488, 26.27687, 
    26.24872, 26.2204,
  23.05567, 23.09728, 23.13875, 23.1801, 23.22131, 23.26239, 23.30333, 
    23.34415, 23.38483, 23.42537, 23.46579, 23.50607, 23.54622, 23.58623, 
    23.62611, 23.66585, 23.70546, 23.74493, 23.78427, 23.82347, 23.86253, 
    23.90146, 23.94025, 23.97891, 24.01743, 24.05581, 24.09405, 24.13216, 
    24.17013, 24.20796, 24.24565, 24.2832, 24.32062, 24.35789, 24.39503, 
    24.43202, 24.46888, 24.50559, 24.54216, 24.5786, 24.61489, 24.65104, 
    24.68705, 24.72292, 24.75865, 24.79423, 24.82968, 24.86497, 24.90013, 
    24.93514, 24.97001, 25.00474, 25.03933, 25.07376, 25.10806, 25.14221, 
    25.17621, 25.21007, 25.24379, 25.27736, 25.31078, 25.34406, 25.37719, 
    25.41018, 25.44302, 25.47571, 25.50825, 25.54065, 25.5729, 25.605, 
    25.63696, 25.66876, 25.70042, 25.73193, 25.76329, 25.7945, 25.82556, 
    25.85647, 25.88724, 25.91785, 25.94831, 25.97862, 26.00878, 26.03879, 
    26.06865, 26.09836, 26.12791, 26.15732, 26.18657, 26.21567, 26.24462, 
    26.27341, 26.30206, 26.33055, 26.35888, 26.38706, 26.41509, 26.44297, 
    26.47069, 26.49825, 26.52567, 26.55293, 26.58003, 26.60697, 26.63377, 
    26.6604, 26.68688, 26.71321, 26.73938, 26.76539, 26.79124, 26.81694, 
    26.84249, 26.86787, 26.8931, 26.91817, 26.94308, 26.96784, 26.99244, 
    27.01687, 27.04115, 27.06528, 27.08924, 27.11304, 27.13668, 27.16017, 
    27.1835, 27.20666, 27.22967, 27.25251, 27.2752, 27.29772, 27.32009, 
    27.34229, 27.36433, 27.38622, 27.40793, 27.42949, 27.45089, 27.47212, 
    27.4932, 27.51411, 27.53486, 27.55544, 27.57587, 27.59613, 27.61622, 
    27.63616, 27.65593, 27.67554, 27.69498, 27.71426, 27.73338, 27.75233, 
    27.77111, 27.78974, 27.8082, 27.82649, 27.84462, 27.86258, 27.88038, 
    27.89802, 27.91548, 27.93279, 27.94992, 27.96689, 27.9837, 28.00034, 
    28.01681, 28.03312, 28.04926, 28.06523, 28.08103, 28.09667, 28.11214, 
    28.12745, 28.14259, 28.15755, 28.17236, 28.18699, 28.20146, 28.21576, 
    28.22989, 28.24385, 28.25764, 28.27127, 28.28473, 28.29801, 28.31113, 
    28.32409, 28.33687, 28.34948, 28.36192, 28.3742, 28.3863, 28.39824, 
    28.41, 28.4216, 28.43302, 28.44428, 28.45537, 28.46628, 28.47703, 
    28.4876, 28.49801, 28.50824, 28.51831, 28.5282, 28.53793, 28.54748, 
    28.55686, 28.56607, 28.57511, 28.58397, 28.59267, 28.6012, 28.60955, 
    28.61773, 28.62575, 28.63359, 28.64125, 28.64875, 28.65608, 28.66323, 
    28.67021, 28.67702, 28.68366, 28.69012, 28.69641, 28.70254, 28.70848, 
    28.71426, 28.71987, 28.7253, 28.73056, 28.73564, 28.74056, 28.7453, 
    28.74987, 28.75427, 28.75849, 28.76254, 28.76642, 28.77013, 28.77366, 
    28.77702, 28.78021, 28.78322, 28.78606, 28.78873, 28.79123, 28.79355, 
    28.7957, 28.79768, 28.79948, 28.80111, 28.80257, 28.80385, 28.80497, 
    28.8059, 28.80667, 28.80726, 28.80768, 28.80793, 28.808, 28.8079, 
    28.80763, 28.80718, 28.80656, 28.80577, 28.8048, 28.80366, 28.80235, 
    28.80087, 28.79921, 28.79738, 28.79537, 28.7932, 28.79084, 28.78832, 
    28.78563, 28.78276, 28.77971, 28.7765, 28.77311, 28.76955, 28.76582, 
    28.76191, 28.75783, 28.75358, 28.74916, 28.74456, 28.73979, 28.73485, 
    28.72974, 28.72445, 28.71899, 28.71336, 28.70756, 28.70158, 28.69543, 
    28.68911, 28.68262, 28.67595, 28.66912, 28.66211, 28.65493, 28.64758, 
    28.64005, 28.63236, 28.62449, 28.61645, 28.60824, 28.59986, 28.59131, 
    28.58258, 28.57369, 28.56462, 28.55539, 28.54598, 28.5364, 28.52665, 
    28.51673, 28.50664, 28.49637, 28.48594, 28.47534, 28.46457, 28.45362, 
    28.44251, 28.43123, 28.41978, 28.40815, 28.39636, 28.3844, 28.37227, 
    28.35997, 28.3475, 28.33486, 28.32205, 28.30907, 28.29592, 28.28261, 
    28.26912, 28.25547, 28.24165, 28.22766, 28.21351, 28.19918, 28.18469, 
    28.17003, 28.1552, 28.1402, 28.12504, 28.10971, 28.09421, 28.07854, 
    28.06271, 28.04671, 28.03055, 28.01422, 27.99772, 27.98105, 27.96422, 
    27.94722, 27.93006, 27.91273, 27.89524, 27.87758, 27.85975, 27.84176, 
    27.82361, 27.80529, 27.7868, 27.76815, 27.74934, 27.73036, 27.71122, 
    27.69192, 27.67245, 27.65281, 27.63302, 27.61306, 27.59293, 27.57265, 
    27.5522, 27.53159, 27.51081, 27.48988, 27.46878, 27.44752, 27.42609, 
    27.40451, 27.38276, 27.36086, 27.33879, 27.31656, 27.29417, 27.27162, 
    27.24891, 27.22604, 27.20301, 27.17982, 27.15647, 27.13296, 27.10929, 
    27.08546, 27.06147, 27.03732, 27.01302, 26.98855, 26.96393, 26.93915, 
    26.91422, 26.88912, 26.86387, 26.83846, 26.81289, 26.78717, 26.76129, 
    26.73525, 26.70905, 26.6827, 26.6562, 26.62954, 26.60272, 26.57575, 
    26.54862, 26.52134, 26.4939, 26.46631, 26.43857, 26.41067, 26.38262, 
    26.35441, 26.32605,
  23.15607, 23.19774, 23.23928, 23.28068, 23.32196, 23.3631, 23.40411, 
    23.44499, 23.48573, 23.52634, 23.56682, 23.60716, 23.64737, 23.68744, 
    23.72738, 23.76719, 23.80685, 23.84639, 23.88579, 23.92505, 23.96417, 
    24.00316, 24.04202, 24.08073, 24.11931, 24.15775, 24.19606, 24.23422, 
    24.27225, 24.31014, 24.34789, 24.3855, 24.42298, 24.46031, 24.4975, 
    24.53456, 24.57147, 24.60824, 24.64488, 24.68137, 24.71772, 24.75393, 
    24.79, 24.82592, 24.86171, 24.89735, 24.93285, 24.9682, 25.00342, 
    25.03849, 25.07341, 25.1082, 25.14284, 25.17733, 25.21168, 25.24589, 
    25.27995, 25.31386, 25.34763, 25.38126, 25.41473, 25.44807, 25.48125, 
    25.51429, 25.54718, 25.57993, 25.61253, 25.64498, 25.67728, 25.70944, 
    25.74144, 25.7733, 25.80501, 25.83657, 25.86799, 25.89925, 25.93036, 
    25.96132, 25.99214, 26.0228, 26.05331, 26.08368, 26.11389, 26.14395, 
    26.17386, 26.20361, 26.23322, 26.26267, 26.29197, 26.32112, 26.35012, 
    26.37896, 26.40765, 26.43619, 26.46457, 26.4928, 26.52088, 26.5488, 
    26.57657, 26.60418, 26.63164, 26.65895, 26.68609, 26.71309, 26.73993, 
    26.76661, 26.79313, 26.8195, 26.84572, 26.87177, 26.89767, 26.92342, 
    26.949, 26.97443, 26.9997, 27.02482, 27.04977, 27.07457, 27.09921, 
    27.12369, 27.14801, 27.17217, 27.19618, 27.22002, 27.24371, 27.26723, 
    27.2906, 27.31381, 27.33685, 27.35974, 27.38246, 27.40503, 27.42743, 
    27.44967, 27.47175, 27.49367, 27.51543, 27.53703, 27.55846, 27.57973, 
    27.60084, 27.62179, 27.64257, 27.6632, 27.68365, 27.70395, 27.72408, 
    27.74405, 27.76386, 27.7835, 27.80298, 27.82229, 27.84144, 27.86043, 
    27.87925, 27.89791, 27.9164, 27.93472, 27.95288, 27.97088, 27.98871, 
    28.00637, 28.02387, 28.04121, 28.05837, 28.07537, 28.09221, 28.10888, 
    28.12538, 28.14171, 28.15788, 28.17388, 28.18972, 28.20539, 28.22088, 
    28.23622, 28.25138, 28.26638, 28.28121, 28.29587, 28.31036, 28.32468, 
    28.33884, 28.35283, 28.36665, 28.38029, 28.39378, 28.40709, 28.42023, 
    28.43321, 28.44601, 28.45865, 28.47111, 28.48341, 28.49553, 28.50749, 
    28.51928, 28.5309, 28.54234, 28.55362, 28.56472, 28.57566, 28.58643, 
    28.59702, 28.60744, 28.6177, 28.62778, 28.63769, 28.64743, 28.657, 
    28.6664, 28.67563, 28.68468, 28.69357, 28.70228, 28.71082, 28.71919, 
    28.72739, 28.73541, 28.74327, 28.75095, 28.75846, 28.7658, 28.77296, 
    28.77996, 28.78678, 28.79343, 28.79991, 28.80621, 28.81234, 28.8183, 
    28.82409, 28.8297, 28.83515, 28.84042, 28.84551, 28.85044, 28.85518, 
    28.85976, 28.86417, 28.8684, 28.87246, 28.87634, 28.88006, 28.8836, 
    28.88696, 28.89016, 28.89318, 28.89602, 28.8987, 28.9012, 28.90352, 
    28.90568, 28.90766, 28.90947, 28.9111, 28.91256, 28.91385, 28.91496, 
    28.9159, 28.91667, 28.91726, 28.91768, 28.91793, 28.918, 28.9179, 
    28.91763, 28.91718, 28.91656, 28.91576, 28.91479, 28.91365, 28.91234, 
    28.91085, 28.90919, 28.90736, 28.90535, 28.90317, 28.90081, 28.89828, 
    28.89558, 28.89271, 28.88966, 28.88644, 28.88305, 28.87948, 28.87574, 
    28.87183, 28.86774, 28.86348, 28.85905, 28.85445, 28.84967, 28.84472, 
    28.83959, 28.8343, 28.82883, 28.82319, 28.81737, 28.81138, 28.80523, 
    28.79889, 28.79239, 28.78571, 28.77886, 28.77184, 28.76465, 28.75728, 
    28.74975, 28.74204, 28.73416, 28.7261, 28.71788, 28.70948, 28.70091, 
    28.69217, 28.68326, 28.67418, 28.66492, 28.6555, 28.6459, 28.63614, 
    28.6262, 28.61609, 28.60581, 28.59536, 28.58473, 28.57394, 28.56298, 
    28.55185, 28.54054, 28.52907, 28.51743, 28.50561, 28.49363, 28.48147, 
    28.46915, 28.45666, 28.444, 28.43117, 28.41816, 28.40499, 28.39165, 
    28.37815, 28.36447, 28.35062, 28.33661, 28.32243, 28.30808, 28.29356, 
    28.27887, 28.26402, 28.24899, 28.2338, 28.21844, 28.20292, 28.18722, 
    28.17136, 28.15534, 28.13914, 28.12278, 28.10625, 28.08956, 28.0727, 
    28.05567, 28.03848, 28.02112, 28.00359, 27.9859, 27.96804, 27.95002, 
    27.93184, 27.91348, 27.89496, 27.87628, 27.85744, 27.83842, 27.81925, 
    27.79991, 27.78041, 27.76074, 27.74091, 27.72091, 27.70075, 27.68043, 
    27.65994, 27.6393, 27.61849, 27.59751, 27.57638, 27.55508, 27.53362, 
    27.512, 27.49022, 27.46827, 27.44616, 27.4239, 27.40147, 27.37888, 
    27.35613, 27.33322, 27.31015, 27.28691, 27.26352, 27.23997, 27.21626, 
    27.19239, 27.16836, 27.14417, 27.11983, 27.09532, 27.07066, 27.04584, 
    27.02085, 26.99572, 26.97042, 26.94497, 26.91936, 26.89359, 26.86766, 
    26.84158, 26.81534, 26.78895, 26.7624, 26.73569, 26.70883, 26.68181, 
    26.65464, 26.62731, 26.59983, 26.57219, 26.5444, 26.51645, 26.48835, 
    26.46009, 26.43169,
  23.25645, 23.29819, 23.33979, 23.38126, 23.4226, 23.4638, 23.50487, 
    23.54581, 23.58662, 23.62729, 23.66783, 23.70823, 23.7485, 23.78864, 
    23.82864, 23.86851, 23.90824, 23.94783, 23.98729, 24.02662, 24.0658, 
    24.10485, 24.14377, 24.18254, 24.22118, 24.25969, 24.29805, 24.33628, 
    24.37436, 24.41231, 24.45012, 24.48779, 24.52533, 24.56272, 24.59997, 
    24.63708, 24.67406, 24.71089, 24.74758, 24.78413, 24.82054, 24.8568, 
    24.89293, 24.92891, 24.96475, 25.00045, 25.03601, 25.07142, 25.10669, 
    25.14182, 25.1768, 25.21164, 25.24634, 25.28089, 25.31529, 25.34955, 
    25.38367, 25.41764, 25.45146, 25.48514, 25.51868, 25.55206, 25.5853, 
    25.6184, 25.65134, 25.68414, 25.71679, 25.7493, 25.78165, 25.81386, 
    25.84592, 25.87783, 25.9096, 25.94121, 25.97267, 26.00399, 26.03515, 
    26.06617, 26.09703, 26.12774, 26.15831, 26.18872, 26.21898, 26.24909, 
    26.27905, 26.30886, 26.33851, 26.36802, 26.39737, 26.42657, 26.45561, 
    26.4845, 26.51324, 26.54183, 26.57026, 26.59854, 26.62666, 26.65463, 
    26.68245, 26.7101, 26.73761, 26.76496, 26.79215, 26.81919, 26.84608, 
    26.8728, 26.89938, 26.92579, 26.95205, 26.97815, 27.0041, 27.02988, 
    27.05551, 27.08098, 27.1063, 27.13146, 27.15645, 27.1813, 27.20598, 
    27.2305, 27.25486, 27.27907, 27.30311, 27.327, 27.35073, 27.37429, 
    27.3977, 27.42094, 27.44403, 27.46696, 27.48972, 27.51232, 27.53477, 
    27.55705, 27.57917, 27.60112, 27.62292, 27.64455, 27.66603, 27.68734, 
    27.70848, 27.72947, 27.75029, 27.77095, 27.79144, 27.81177, 27.83194, 
    27.85195, 27.87179, 27.89146, 27.91097, 27.93032, 27.94951, 27.96852, 
    27.98738, 28.00607, 28.02459, 28.04295, 28.06114, 28.07917, 28.09703, 
    28.11473, 28.13226, 28.14962, 28.16682, 28.18385, 28.20072, 28.21741, 
    28.23395, 28.25031, 28.26651, 28.28254, 28.2984, 28.31409, 28.32962, 
    28.34498, 28.36017, 28.3752, 28.39005, 28.40474, 28.41926, 28.43361, 
    28.44779, 28.4618, 28.47565, 28.48932, 28.50282, 28.51616, 28.52933, 
    28.54232, 28.55515, 28.56781, 28.5803, 28.59262, 28.60477, 28.61674, 
    28.62855, 28.64019, 28.65166, 28.66295, 28.67408, 28.68504, 28.69582, 
    28.70644, 28.71688, 28.72715, 28.73725, 28.74718, 28.75694, 28.76653, 
    28.77594, 28.78518, 28.79426, 28.80316, 28.81189, 28.82044, 28.82883, 
    28.83704, 28.84508, 28.85295, 28.86065, 28.86817, 28.87552, 28.8827, 
    28.88971, 28.89654, 28.9032, 28.90969, 28.91601, 28.92215, 28.92812, 
    28.93392, 28.93954, 28.94499, 28.95027, 28.95538, 28.96031, 28.96507, 
    28.96966, 28.97407, 28.97831, 28.98238, 28.98627, 28.98999, 28.99353, 
    28.99691, 29.0001, 29.00313, 29.00598, 29.00866, 29.01117, 29.0135, 
    29.01566, 29.01764, 29.01945, 29.02109, 29.02255, 29.02384, 29.02495, 
    29.0259, 29.02666, 29.02726, 29.02768, 29.02793, 29.028, 29.0279, 
    29.02762, 29.02718, 29.02655, 29.02576, 29.02479, 29.02365, 29.02233, 
    29.02084, 29.01917, 29.01734, 29.01533, 29.01314, 29.01078, 29.00825, 
    29.00554, 29.00266, 28.99961, 28.99638, 28.99298, 28.98941, 28.98566, 
    28.98174, 28.97765, 28.97338, 28.96894, 28.96433, 28.95954, 28.95458, 
    28.94945, 28.94414, 28.93867, 28.93301, 28.92719, 28.92119, 28.91502, 
    28.90868, 28.90216, 28.89547, 28.88861, 28.88158, 28.87437, 28.86699, 
    28.85944, 28.85172, 28.84382, 28.83575, 28.82751, 28.8191, 28.81052, 
    28.80176, 28.79283, 28.78373, 28.77446, 28.76502, 28.75541, 28.74562, 
    28.73566, 28.72554, 28.71524, 28.70477, 28.69413, 28.68332, 28.67233, 
    28.66118, 28.64985, 28.63836, 28.6267, 28.61486, 28.60286, 28.59068, 
    28.57833, 28.56582, 28.55313, 28.54028, 28.52726, 28.51406, 28.5007, 
    28.48717, 28.47346, 28.45959, 28.44556, 28.43135, 28.41697, 28.40243, 
    28.38771, 28.37283, 28.35778, 28.34256, 28.32718, 28.31162, 28.2959, 
    28.28001, 28.26396, 28.24773, 28.23134, 28.21478, 28.19806, 28.18117, 
    28.16411, 28.14689, 28.1295, 28.11194, 28.09422, 28.07633, 28.05828, 
    28.04006, 28.02167, 28.00312, 27.98441, 27.96553, 27.94648, 27.92727, 
    27.9079, 27.88836, 27.86866, 27.84879, 27.82876, 27.80857, 27.78821, 
    27.76769, 27.74701, 27.72616, 27.70515, 27.68398, 27.66264, 27.64114, 
    27.61948, 27.59766, 27.57568, 27.55353, 27.53123, 27.50876, 27.48613, 
    27.46334, 27.44039, 27.41728, 27.39401, 27.37057, 27.34698, 27.32323, 
    27.29932, 27.27525, 27.25102, 27.22663, 27.20208, 27.17738, 27.15251, 
    27.12749, 27.1023, 27.07697, 27.05147, 27.02581, 27, 26.97403, 26.94791, 
    26.92162, 26.89518, 26.86859, 26.84184, 26.81493, 26.78786, 26.76064, 
    26.73327, 26.70574, 26.67805, 26.65022, 26.62222, 26.59407, 26.56577, 
    26.53732,
  23.35682, 23.39862, 23.44028, 23.48182, 23.52322, 23.56449, 23.60562, 
    23.64662, 23.68749, 23.72823, 23.76883, 23.80929, 23.84963, 23.88982, 
    23.92989, 23.96981, 24.00961, 24.04926, 24.08879, 24.12817, 24.16742, 
    24.20653, 24.2455, 24.28434, 24.32304, 24.3616, 24.40003, 24.43831, 
    24.47646, 24.51447, 24.55234, 24.59007, 24.62766, 24.66511, 24.70242, 
    24.7396, 24.77663, 24.81352, 24.85027, 24.88687, 24.92334, 24.95967, 
    24.99585, 25.03189, 25.06779, 25.10355, 25.13916, 25.17463, 25.20996, 
    25.24514, 25.28018, 25.31507, 25.34982, 25.38443, 25.41889, 25.45321, 
    25.48738, 25.52141, 25.55528, 25.58902, 25.62261, 25.65605, 25.68934, 
    25.72249, 25.75549, 25.78834, 25.82105, 25.85361, 25.88602, 25.91828, 
    25.95039, 25.98235, 26.01417, 26.04583, 26.07735, 26.10872, 26.13993, 
    26.171, 26.20192, 26.23268, 26.26329, 26.29376, 26.32407, 26.35423, 
    26.38424, 26.4141, 26.4438, 26.47335, 26.50275, 26.532, 26.56109, 
    26.59003, 26.61882, 26.64746, 26.67594, 26.70426, 26.73243, 26.76045, 
    26.78831, 26.81602, 26.84357, 26.87097, 26.89821, 26.92529, 26.95222, 
    26.97899, 27.00561, 27.03207, 27.05837, 27.08452, 27.11051, 27.13634, 
    27.16201, 27.18753, 27.21289, 27.23809, 27.26313, 27.28801, 27.31274, 
    27.3373, 27.36171, 27.38596, 27.41004, 27.43397, 27.45774, 27.48134, 
    27.50479, 27.52808, 27.5512, 27.57417, 27.59697, 27.61962, 27.6421, 
    27.66442, 27.68657, 27.70857, 27.73041, 27.75208, 27.77359, 27.79493, 
    27.81612, 27.83714, 27.858, 27.87869, 27.89922, 27.91959, 27.93979, 
    27.95983, 27.97971, 27.99942, 28.01897, 28.03835, 28.05757, 28.07662, 
    28.0955, 28.11423, 28.13278, 28.15117, 28.1694, 28.18746, 28.20535, 
    28.22308, 28.24064, 28.25804, 28.27527, 28.29233, 28.30922, 28.32595, 
    28.34251, 28.3589, 28.37513, 28.39119, 28.40708, 28.4228, 28.43836, 
    28.45374, 28.46896, 28.48401, 28.4989, 28.51361, 28.52815, 28.54253, 
    28.55674, 28.57077, 28.58464, 28.59834, 28.61187, 28.62523, 28.63842, 
    28.65144, 28.66429, 28.67698, 28.68949, 28.70183, 28.714, 28.726, 
    28.73783, 28.74949, 28.76097, 28.77229, 28.78344, 28.79441, 28.80522, 
    28.81585, 28.82631, 28.8366, 28.84672, 28.85667, 28.86645, 28.87605, 
    28.88548, 28.89474, 28.90383, 28.91275, 28.92149, 28.93006, 28.93846, 
    28.94669, 28.95475, 28.96263, 28.97034, 28.97788, 28.98524, 28.99243, 
    28.99945, 29.0063, 29.01297, 29.01947, 29.0258, 29.03196, 29.03794, 
    29.04375, 29.04938, 29.05484, 29.06013, 29.06525, 29.07019, 29.07495, 
    29.07955, 29.08397, 29.08822, 29.09229, 29.09619, 29.09992, 29.10347, 
    29.10685, 29.11005, 29.11308, 29.11594, 29.11863, 29.12114, 29.12347, 
    29.12563, 29.12762, 29.12943, 29.13107, 29.13254, 29.13383, 29.13495, 
    29.13589, 29.13666, 29.13726, 29.13768, 29.13793, 29.138, 29.1379, 
    29.13762, 29.13717, 29.13655, 29.13576, 29.13478, 29.13364, 29.13232, 
    29.13083, 29.12916, 29.12732, 29.1253, 29.12311, 29.12075, 29.11821, 
    29.1155, 29.11262, 29.10956, 29.10633, 29.10292, 29.09934, 29.09559, 
    29.09166, 29.08756, 29.08328, 29.07883, 29.07421, 29.06942, 29.06445, 
    29.05931, 29.05399, 29.0485, 29.04284, 29.037, 29.03099, 29.02481, 
    29.01846, 29.01193, 29.00523, 28.99836, 28.99131, 28.98409, 28.9767, 
    28.96913, 28.96139, 28.95348, 28.9454, 28.93715, 28.92872, 28.92012, 
    28.91135, 28.9024, 28.89329, 28.884, 28.87454, 28.86491, 28.85511, 
    28.84513, 28.83499, 28.82467, 28.81418, 28.80352, 28.79269, 28.78168, 
    28.77051, 28.75917, 28.74765, 28.73597, 28.72411, 28.71208, 28.69988, 
    28.68752, 28.67498, 28.66227, 28.64939, 28.63635, 28.62313, 28.60974, 
    28.59619, 28.58246, 28.56856, 28.5545, 28.54027, 28.52586, 28.51129, 
    28.49655, 28.48164, 28.46657, 28.45132, 28.43591, 28.42033, 28.40458, 
    28.38866, 28.37258, 28.35632, 28.3399, 28.32332, 28.30656, 28.28964, 
    28.27255, 28.2553, 28.23788, 28.22029, 28.20254, 28.18461, 28.16653, 
    28.14828, 28.12986, 28.11128, 28.09253, 28.07361, 28.05454, 28.03529, 
    28.01588, 27.99631, 27.97657, 27.95667, 27.93661, 27.91638, 27.89598, 
    27.87543, 27.85471, 27.83382, 27.81278, 27.79157, 27.7702, 27.74866, 
    27.72696, 27.7051, 27.68308, 27.6609, 27.63855, 27.61604, 27.59338, 
    27.57055, 27.54756, 27.5244, 27.50109, 27.47762, 27.45399, 27.43019, 
    27.40624, 27.38213, 27.35786, 27.33343, 27.30884, 27.28409, 27.25918, 
    27.23411, 27.20889, 27.18351, 27.15796, 27.13227, 27.10641, 27.08039, 
    27.05422, 27.0279, 27.00141, 26.97477, 26.94797, 26.92102, 26.89391, 
    26.86664, 26.83922, 26.81165, 26.78391, 26.75603, 26.72799, 26.69979, 
    26.67144, 26.64294,
  23.45718, 23.49904, 23.54077, 23.58236, 23.62383, 23.66516, 23.70635, 
    23.74742, 23.78835, 23.82915, 23.86981, 23.91034, 23.95074, 23.99099, 
    24.03112, 24.07111, 24.11096, 24.15068, 24.19026, 24.22971, 24.26902, 
    24.30819, 24.34723, 24.38612, 24.42488, 24.4635, 24.50199, 24.54034, 
    24.57854, 24.61661, 24.65454, 24.69233, 24.72998, 24.76749, 24.80486, 
    24.84209, 24.87918, 24.91613, 24.95294, 24.98961, 25.02613, 25.06252, 
    25.09876, 25.13486, 25.17081, 25.20662, 25.2423, 25.27782, 25.31321, 
    25.34845, 25.38354, 25.41849, 25.4533, 25.48796, 25.52248, 25.55685, 
    25.59108, 25.62516, 25.6591, 25.69288, 25.72653, 25.76002, 25.79337, 
    25.82657, 25.85963, 25.89253, 25.92529, 25.9579, 25.99037, 26.02268, 
    26.05485, 26.08686, 26.11873, 26.15045, 26.18202, 26.21344, 26.2447, 
    26.27582, 26.30679, 26.3376, 26.36827, 26.39878, 26.42915, 26.45936, 
    26.48942, 26.51933, 26.54908, 26.57868, 26.60813, 26.63743, 26.66657, 
    26.69556, 26.72439, 26.75308, 26.7816, 26.80998, 26.8382, 26.86626, 
    26.89417, 26.92192, 26.94952, 26.97696, 27.00425, 27.03138, 27.05836, 
    27.08518, 27.11184, 27.13834, 27.16469, 27.19088, 27.21692, 27.24279, 
    27.26851, 27.29407, 27.31947, 27.34472, 27.3698, 27.39473, 27.41949, 
    27.4441, 27.46855, 27.49284, 27.51697, 27.54093, 27.56474, 27.58839, 
    27.61188, 27.63521, 27.65837, 27.68138, 27.70422, 27.7269, 27.74942, 
    27.77178, 27.79398, 27.81601, 27.83788, 27.8596, 27.88114, 27.90253, 
    27.92375, 27.94481, 27.9657, 27.98643, 28.007, 28.0274, 28.04764, 
    28.06771, 28.08763, 28.10737, 28.12695, 28.14637, 28.16562, 28.18471, 
    28.20363, 28.22238, 28.24097, 28.2594, 28.27765, 28.29575, 28.31367, 
    28.33143, 28.34902, 28.36645, 28.38371, 28.4008, 28.41772, 28.43448, 
    28.45107, 28.46749, 28.48375, 28.49984, 28.51576, 28.53151, 28.54709, 
    28.5625, 28.57775, 28.59283, 28.60774, 28.62248, 28.63705, 28.65145, 
    28.66568, 28.67974, 28.69364, 28.70736, 28.72091, 28.7343, 28.74751, 
    28.76056, 28.77343, 28.78614, 28.79867, 28.81103, 28.82323, 28.83525, 
    28.8471, 28.85878, 28.87029, 28.88162, 28.89279, 28.90379, 28.91461, 
    28.92526, 28.93574, 28.94605, 28.95619, 28.96616, 28.97595, 28.98557, 
    28.99502, 29.0043, 29.0134, 29.02234, 29.0311, 29.03968, 29.0481, 
    29.05634, 29.06441, 29.07231, 29.08003, 29.08759, 29.09496, 29.10217, 
    29.1092, 29.11606, 29.12275, 29.12926, 29.1356, 29.14176, 29.14775, 
    29.15357, 29.15922, 29.16469, 29.16999, 29.17511, 29.18006, 29.18484, 
    29.18944, 29.19387, 29.19813, 29.20221, 29.20612, 29.20985, 29.21341, 
    29.21679, 29.22, 29.22304, 29.2259, 29.22859, 29.2311, 29.23344, 
    29.23561, 29.2376, 29.23942, 29.24106, 29.24253, 29.24382, 29.24494, 
    29.24589, 29.24666, 29.24726, 29.24768, 29.24793, 29.248, 29.2479, 
    29.24762, 29.24717, 29.24655, 29.24575, 29.24478, 29.24363, 29.24231, 
    29.24081, 29.23914, 29.2373, 29.23528, 29.23309, 29.23072, 29.22818, 
    29.22546, 29.22257, 29.21951, 29.21627, 29.21286, 29.20927, 29.20551, 
    29.20157, 29.19747, 29.19318, 29.18873, 29.1841, 29.17929, 29.17431, 
    29.16916, 29.16384, 29.15834, 29.15266, 29.14682, 29.1408, 29.13461, 
    29.12824, 29.1217, 29.11499, 29.1081, 29.10104, 29.09381, 29.0864, 
    29.07882, 29.07107, 29.06315, 29.05505, 29.04678, 29.03834, 29.02972, 
    29.02094, 29.01197, 29.00284, 28.99354, 28.98406, 28.97441, 28.96459, 
    28.9546, 28.94443, 28.9341, 28.92359, 28.91291, 28.90206, 28.89104, 
    28.87984, 28.86848, 28.85694, 28.84523, 28.83336, 28.82131, 28.80909, 
    28.7967, 28.78414, 28.77141, 28.75851, 28.74543, 28.73219, 28.71878, 
    28.7052, 28.69145, 28.67753, 28.66344, 28.64918, 28.63475, 28.62016, 
    28.60539, 28.59045, 28.57535, 28.56008, 28.54464, 28.52903, 28.51325, 
    28.4973, 28.48119, 28.46491, 28.44846, 28.43184, 28.41506, 28.39811, 
    28.38099, 28.3637, 28.34625, 28.32863, 28.31085, 28.2929, 28.27478, 
    28.25649, 28.23804, 28.21943, 28.20065, 28.1817, 28.16259, 28.14331, 
    28.12387, 28.10426, 28.08449, 28.06455, 28.04445, 28.02419, 28.00376, 
    27.98316, 27.96241, 27.94148, 27.9204, 27.89915, 27.87774, 27.85617, 
    27.83444, 27.81254, 27.79048, 27.76826, 27.74587, 27.72333, 27.70062, 
    27.67775, 27.65472, 27.63153, 27.60817, 27.58466, 27.56099, 27.53715, 
    27.51316, 27.48901, 27.46469, 27.44022, 27.41558, 27.39079, 27.36584, 
    27.34073, 27.31546, 27.29004, 27.26445, 27.23871, 27.21281, 27.18675, 
    27.16054, 27.13416, 27.10763, 27.08095, 27.0541, 27.0271, 26.99995, 
    26.97264, 26.94517, 26.91754, 26.88976, 26.86183, 26.83374, 26.8055, 
    26.7771, 26.74855,
  23.55752, 23.59944, 23.64123, 23.68289, 23.72442, 23.76581, 23.80707, 
    23.8482, 23.88919, 23.93005, 23.97078, 24.01137, 24.05183, 24.09215, 
    24.13234, 24.17239, 24.2123, 24.25208, 24.29173, 24.33123, 24.3706, 
    24.40984, 24.44893, 24.48789, 24.52671, 24.5654, 24.60394, 24.64235, 
    24.68061, 24.71874, 24.75673, 24.79458, 24.83229, 24.86986, 24.90729, 
    24.94458, 24.98173, 25.01874, 25.0556, 25.09233, 25.12891, 25.16535, 
    25.20165, 25.23781, 25.27382, 25.30969, 25.34542, 25.381, 25.41644, 
    25.45174, 25.48689, 25.5219, 25.55677, 25.59148, 25.62606, 25.66049, 
    25.69477, 25.7289, 25.76289, 25.79674, 25.83044, 25.86399, 25.89739, 
    25.93065, 25.96375, 25.99672, 26.02953, 26.06219, 26.09471, 26.12708, 
    26.15929, 26.19136, 26.22328, 26.25505, 26.28667, 26.31815, 26.34947, 
    26.38063, 26.41165, 26.44252, 26.47324, 26.5038, 26.53422, 26.56448, 
    26.59459, 26.62454, 26.65435, 26.684, 26.7135, 26.74284, 26.77204, 
    26.80107, 26.82996, 26.85869, 26.88726, 26.91569, 26.94395, 26.97206, 
    27.00002, 27.02782, 27.05547, 27.08296, 27.11029, 27.13747, 27.16449, 
    27.19135, 27.21806, 27.24461, 27.271, 27.29724, 27.32332, 27.34924, 
    27.375, 27.4006, 27.42605, 27.45134, 27.47646, 27.50143, 27.52624, 
    27.55089, 27.57538, 27.59971, 27.62388, 27.64789, 27.67174, 27.69543, 
    27.71896, 27.74233, 27.76553, 27.78858, 27.81146, 27.83418, 27.85674, 
    27.87914, 27.90138, 27.92345, 27.94536, 27.96711, 27.98869, 28.01011, 
    28.03137, 28.05247, 28.0734, 28.09417, 28.11477, 28.13521, 28.15548, 
    28.17559, 28.19554, 28.21532, 28.23494, 28.25439, 28.27367, 28.29279, 
    28.31175, 28.33053, 28.34916, 28.36761, 28.3859, 28.40403, 28.42199, 
    28.43978, 28.4574, 28.47486, 28.49215, 28.50927, 28.52622, 28.54301, 
    28.55963, 28.57608, 28.59237, 28.60848, 28.62443, 28.64021, 28.65582, 
    28.67126, 28.68653, 28.70164, 28.71658, 28.73134, 28.74594, 28.76036, 
    28.77462, 28.78871, 28.80263, 28.81638, 28.82996, 28.84336, 28.8566, 
    28.86967, 28.88257, 28.8953, 28.90785, 28.92024, 28.93245, 28.94449, 
    28.95637, 28.96807, 28.9796, 28.99096, 29.00214, 29.01316, 29.024, 
    29.03467, 29.04517, 29.0555, 29.06566, 29.07564, 29.08545, 29.09509, 
    29.10456, 29.11385, 29.12297, 29.13192, 29.1407, 29.1493, 29.15773, 
    29.16599, 29.17408, 29.18199, 29.18973, 29.19729, 29.20468, 29.2119, 
    29.21895, 29.22582, 29.23252, 29.23904, 29.24539, 29.25157, 29.25757, 
    29.2634, 29.26906, 29.27454, 29.27985, 29.28498, 29.28994, 29.29472, 
    29.29934, 29.30377, 29.30803, 29.31212, 29.31604, 29.31978, 29.32334, 
    29.32673, 29.32995, 29.33299, 29.33586, 29.33855, 29.34107, 29.34342, 
    29.34559, 29.34758, 29.3494, 29.35105, 29.35252, 29.35382, 29.35494, 
    29.35588, 29.35666, 29.35725, 29.35768, 29.35793, 29.358, 29.3579, 
    29.35762, 29.35717, 29.35655, 29.35575, 29.35477, 29.35362, 29.3523, 
    29.3508, 29.34913, 29.34728, 29.34526, 29.34306, 29.34069, 29.33814, 
    29.33542, 29.33253, 29.32945, 29.32621, 29.32279, 29.3192, 29.31543, 
    29.31149, 29.30737, 29.30308, 29.29862, 29.29398, 29.28917, 29.28418, 
    29.27902, 29.27368, 29.26817, 29.26249, 29.25663, 29.2506, 29.2444, 
    29.23802, 29.23147, 29.22474, 29.21784, 29.21077, 29.20353, 29.19611, 
    29.18851, 29.18075, 29.17281, 29.1647, 29.15641, 29.14795, 29.13932, 
    29.13052, 29.12154, 29.11239, 29.10307, 29.09358, 29.08391, 29.07407, 
    29.06406, 29.05388, 29.04352, 29.033, 29.0223, 29.01143, 29.00039, 
    28.98917, 28.97779, 28.96623, 28.9545, 28.9426, 28.93053, 28.91829, 
    28.90588, 28.89329, 28.88054, 28.86762, 28.85452, 28.84126, 28.82782, 
    28.81421, 28.80044, 28.7865, 28.77238, 28.75809, 28.74364, 28.72902, 
    28.71422, 28.69926, 28.68413, 28.66883, 28.65336, 28.63772, 28.62192, 
    28.60595, 28.5898, 28.57349, 28.55701, 28.54037, 28.52355, 28.50657, 
    28.48942, 28.47211, 28.45462, 28.43697, 28.41916, 28.40117, 28.38302, 
    28.36471, 28.34622, 28.32757, 28.30876, 28.28978, 28.27063, 28.25132, 
    28.23184, 28.2122, 28.1924, 28.17242, 28.15229, 28.13199, 28.11152, 
    28.09089, 28.0701, 28.04914, 28.02802, 28.00674, 27.98529, 27.96368, 
    27.94191, 27.91997, 27.89787, 27.87561, 27.85319, 27.8306, 27.80785, 
    27.78494, 27.76187, 27.73864, 27.71525, 27.6917, 27.66798, 27.64411, 
    27.62007, 27.59587, 27.57152, 27.547, 27.52233, 27.49749, 27.4725, 
    27.44735, 27.42203, 27.39656, 27.37094, 27.34515, 27.3192, 27.2931, 
    27.26684, 27.24042, 27.21385, 27.18711, 27.16022, 27.13318, 27.10598, 
    27.07862, 27.0511, 27.02343, 26.99561, 26.96763, 26.93949, 26.9112, 
    26.88275, 26.85415,
  23.65784, 23.69983, 23.74168, 23.78341, 23.825, 23.86645, 23.90778, 
    23.94897, 23.99002, 24.03094, 24.07173, 24.11239, 24.15291, 24.19329, 
    24.23354, 24.27365, 24.31363, 24.35347, 24.39318, 24.43274, 24.47218, 
    24.51147, 24.55063, 24.58965, 24.62853, 24.66727, 24.70588, 24.74434, 
    24.78267, 24.82086, 24.85891, 24.89682, 24.93459, 24.97222, 25.00971, 
    25.04705, 25.08426, 25.12133, 25.15825, 25.19504, 25.23168, 25.26818, 
    25.30453, 25.34075, 25.37682, 25.41275, 25.44853, 25.48417, 25.51967, 
    25.55503, 25.59023, 25.6253, 25.66022, 25.69499, 25.72962, 25.76411, 
    25.79844, 25.83264, 25.86668, 25.90058, 25.93433, 25.96794, 26.0014, 
    26.03471, 26.06787, 26.10089, 26.13375, 26.16647, 26.19904, 26.23146, 
    26.26373, 26.29585, 26.32783, 26.35965, 26.39132, 26.42285, 26.45422, 
    26.48544, 26.51651, 26.54743, 26.5782, 26.60881, 26.63927, 26.66959, 
    26.69975, 26.72975, 26.75961, 26.78931, 26.81886, 26.84825, 26.87749, 
    26.90658, 26.93551, 26.96429, 26.99292, 27.02139, 27.0497, 27.07786, 
    27.10586, 27.13371, 27.1614, 27.18894, 27.21632, 27.24354, 27.27061, 
    27.29752, 27.32427, 27.35087, 27.37731, 27.40359, 27.42971, 27.45568, 
    27.48148, 27.50713, 27.53262, 27.55795, 27.58312, 27.60813, 27.63298, 
    27.65768, 27.68221, 27.70658, 27.73079, 27.75484, 27.77874, 27.80247, 
    27.82604, 27.84944, 27.87269, 27.89577, 27.9187, 27.94146, 27.96406, 
    27.9865, 28.00877, 28.03088, 28.05283, 28.07462, 28.09624, 28.1177, 
    28.13899, 28.16013, 28.18109, 28.2019, 28.22254, 28.24301, 28.26332, 
    28.28347, 28.30345, 28.32327, 28.34291, 28.3624, 28.38172, 28.40087, 
    28.41986, 28.43868, 28.45734, 28.47583, 28.49415, 28.51231, 28.5303, 
    28.54812, 28.56577, 28.58326, 28.60058, 28.61773, 28.63472, 28.65154, 
    28.66819, 28.68467, 28.70098, 28.71712, 28.7331, 28.74891, 28.76455, 
    28.78002, 28.79532, 28.81045, 28.82541, 28.8402, 28.85483, 28.86928, 
    28.88356, 28.89768, 28.91162, 28.92539, 28.939, 28.95243, 28.96569, 
    28.97878, 28.9917, 29.00445, 29.01703, 29.02944, 29.04168, 29.05374, 
    29.06564, 29.07736, 29.08891, 29.10029, 29.11149, 29.12253, 29.13339, 
    29.14408, 29.1546, 29.16495, 29.17513, 29.18513, 29.19496, 29.20461, 
    29.2141, 29.22341, 29.23255, 29.24151, 29.2503, 29.25892, 29.26737, 
    29.27564, 29.28374, 29.29167, 29.29942, 29.307, 29.3144, 29.32163, 
    29.32869, 29.33558, 29.34229, 29.34882, 29.35518, 29.36137, 29.36739, 
    29.37323, 29.37889, 29.38439, 29.3897, 29.39485, 29.39981, 29.40461, 
    29.40923, 29.41367, 29.41794, 29.42204, 29.42596, 29.42971, 29.43328, 
    29.43668, 29.4399, 29.44295, 29.44582, 29.44852, 29.45104, 29.45339, 
    29.45556, 29.45756, 29.45939, 29.46104, 29.46251, 29.46381, 29.46493, 
    29.46588, 29.46665, 29.46725, 29.46768, 29.46793, 29.468, 29.4679, 
    29.46762, 29.46717, 29.46654, 29.46574, 29.46477, 29.46362, 29.46229, 
    29.46079, 29.45911, 29.45726, 29.45523, 29.45303, 29.45065, 29.4481, 
    29.44538, 29.44248, 29.4394, 29.43615, 29.43273, 29.42913, 29.42535, 
    29.4214, 29.41728, 29.41298, 29.40851, 29.40386, 29.39904, 29.39404, 
    29.38887, 29.38353, 29.37801, 29.37232, 29.36645, 29.36041, 29.35419, 
    29.3478, 29.34124, 29.3345, 29.32759, 29.3205, 29.31324, 29.30581, 
    29.2982, 29.29042, 29.28247, 29.27434, 29.26604, 29.25757, 29.24892, 
    29.2401, 29.23111, 29.22194, 29.21261, 29.2031, 29.19341, 29.18356, 
    29.17353, 29.16332, 29.15295, 29.1424, 29.13169, 29.1208, 29.10973, 
    29.0985, 29.08709, 29.07552, 29.06377, 29.05185, 29.03975, 29.02749, 
    29.01505, 29.00245, 28.98967, 28.97672, 28.96361, 28.95032, 28.93686, 
    28.92323, 28.90943, 28.89546, 28.88132, 28.86701, 28.85253, 28.83788, 
    28.82306, 28.80807, 28.79291, 28.77758, 28.76208, 28.74642, 28.73059, 
    28.71458, 28.69841, 28.68207, 28.66556, 28.64889, 28.63204, 28.61503, 
    28.59785, 28.58051, 28.56299, 28.54531, 28.52746, 28.50945, 28.49126, 
    28.47291, 28.4544, 28.43572, 28.41687, 28.39785, 28.37868, 28.35933, 
    28.33982, 28.32014, 28.3003, 28.28029, 28.26012, 28.23978, 28.21928, 
    28.19862, 28.17779, 28.15679, 28.13564, 28.11432, 28.09283, 28.07118, 
    28.04937, 28.0274, 28.00526, 27.98296, 27.96049, 27.93787, 27.91508, 
    27.89214, 27.86902, 27.84575, 27.82232, 27.79872, 27.77497, 27.75105, 
    27.72697, 27.70274, 27.67834, 27.65378, 27.62906, 27.60419, 27.57915, 
    27.55395, 27.5286, 27.50308, 27.47741, 27.45158, 27.42559, 27.39944, 
    27.37314, 27.34667, 27.32005, 27.29327, 27.26634, 27.23925, 27.212, 
    27.1846, 27.15703, 27.12932, 27.10144, 27.07342, 27.04523, 27.01689, 
    26.9884, 26.95975,
  23.75815, 23.8002, 23.84212, 23.8839, 23.92556, 23.96708, 24.00846, 
    24.04972, 24.09084, 24.13182, 24.17267, 24.21339, 24.25397, 24.29442, 
    24.33473, 24.3749, 24.41494, 24.45485, 24.49461, 24.53424, 24.57373, 
    24.61309, 24.65231, 24.69139, 24.73033, 24.76913, 24.8078, 24.84633, 
    24.88471, 24.92296, 24.96107, 24.99904, 25.03687, 25.07456, 25.11211, 
    25.14952, 25.18678, 25.22391, 25.26089, 25.29773, 25.33443, 25.37099, 
    25.40741, 25.44368, 25.47981, 25.51579, 25.55164, 25.58733, 25.62289, 
    25.6583, 25.69356, 25.72869, 25.76366, 25.79849, 25.83318, 25.86772, 
    25.90211, 25.93636, 25.97046, 26.00441, 26.03822, 26.07188, 26.10539, 
    26.13876, 26.17198, 26.20504, 26.23796, 26.27074, 26.30336, 26.33583, 
    26.36816, 26.40034, 26.43236, 26.46424, 26.49596, 26.52753, 26.55896, 
    26.59023, 26.62135, 26.65232, 26.68314, 26.71381, 26.74433, 26.77469, 
    26.8049, 26.83496, 26.86486, 26.89461, 26.92421, 26.95365, 26.98294, 
    27.01208, 27.04106, 27.06989, 27.09856, 27.12708, 27.15544, 27.18365, 
    27.2117, 27.23959, 27.26733, 27.29492, 27.32234, 27.34961, 27.37672, 
    27.40368, 27.43048, 27.45712, 27.4836, 27.50993, 27.5361, 27.56211, 
    27.58796, 27.61365, 27.63918, 27.66455, 27.68977, 27.71482, 27.73972, 
    27.76445, 27.78903, 27.81344, 27.8377, 27.86179, 27.88573, 27.9095, 
    27.93311, 27.95655, 27.97984, 28.00297, 28.02593, 28.04873, 28.07137, 
    28.09385, 28.11616, 28.13831, 28.1603, 28.18212, 28.20378, 28.22528, 
    28.24661, 28.26778, 28.28878, 28.30962, 28.3303, 28.35081, 28.37116, 
    28.39134, 28.41135, 28.4312, 28.45089, 28.47041, 28.48976, 28.50895, 
    28.52797, 28.54683, 28.56552, 28.58404, 28.60239, 28.62058, 28.6386, 
    28.65646, 28.67414, 28.69166, 28.70901, 28.7262, 28.74321, 28.76006, 
    28.77674, 28.79325, 28.80959, 28.82577, 28.84177, 28.8576, 28.87327, 
    28.88877, 28.9041, 28.91926, 28.93425, 28.94906, 28.96371, 28.97819, 
    28.9925, 29.00664, 29.02061, 29.03441, 29.04803, 29.06149, 29.07478, 
    29.08789, 29.10084, 29.11361, 29.12621, 29.13864, 29.1509, 29.16299, 
    29.1749, 29.18665, 29.19822, 29.20962, 29.22084, 29.2319, 29.24278, 
    29.25349, 29.26403, 29.2744, 29.28459, 29.29461, 29.30446, 29.31413, 
    29.32363, 29.33296, 29.34212, 29.3511, 29.35991, 29.36854, 29.377, 
    29.38529, 29.3934, 29.40134, 29.40911, 29.4167, 29.42412, 29.43137, 
    29.43844, 29.44533, 29.45206, 29.4586, 29.46498, 29.47118, 29.4772, 
    29.48305, 29.48873, 29.49423, 29.49956, 29.50471, 29.50969, 29.51449, 
    29.51912, 29.52357, 29.52785, 29.53196, 29.53588, 29.53964, 29.54322, 
    29.54662, 29.54985, 29.5529, 29.55578, 29.55848, 29.56101, 29.56336, 
    29.56554, 29.56754, 29.56937, 29.57102, 29.5725, 29.5738, 29.57493, 
    29.57588, 29.57665, 29.57725, 29.57768, 29.57793, 29.578, 29.5779, 
    29.57762, 29.57717, 29.57654, 29.57574, 29.57476, 29.57361, 29.57228, 
    29.57077, 29.56909, 29.56724, 29.56521, 29.563, 29.56062, 29.55807, 
    29.55534, 29.55243, 29.54935, 29.54609, 29.54266, 29.53906, 29.53527, 
    29.53132, 29.52719, 29.52288, 29.5184, 29.51374, 29.50891, 29.50391, 
    29.49873, 29.49337, 29.48784, 29.48214, 29.47626, 29.47021, 29.46398, 
    29.45758, 29.451, 29.44425, 29.43733, 29.43023, 29.42296, 29.41551, 
    29.40789, 29.4001, 29.39213, 29.38399, 29.37568, 29.36719, 29.35852, 
    29.34969, 29.34068, 29.3315, 29.32214, 29.31261, 29.30291, 29.29304, 
    29.28299, 29.27277, 29.26238, 29.25181, 29.24107, 29.23016, 29.21908, 
    29.20782, 29.1964, 29.1848, 29.17303, 29.16109, 29.14897, 29.13669, 
    29.12423, 29.1116, 29.0988, 29.08583, 29.07269, 29.05938, 29.04589, 
    29.03224, 29.01841, 29.00442, 28.99025, 28.97591, 28.96141, 28.94673, 
    28.93188, 28.91687, 28.90168, 28.88633, 28.87081, 28.85511, 28.83925, 
    28.82322, 28.80702, 28.79065, 28.77411, 28.75741, 28.74053, 28.72349, 
    28.70628, 28.6889, 28.67136, 28.65364, 28.63576, 28.61772, 28.5995, 
    28.58112, 28.56257, 28.54386, 28.52497, 28.50593, 28.48671, 28.46733, 
    28.44779, 28.42808, 28.4082, 28.38816, 28.36795, 28.34758, 28.32704, 
    28.30634, 28.28547, 28.26444, 28.24325, 28.22189, 28.20037, 28.17868, 
    28.15683, 28.13482, 28.11264, 28.0903, 28.0678, 28.04514, 28.02231, 
    27.99932, 27.97617, 27.95286, 27.92938, 27.90575, 27.88195, 27.85799, 
    27.83387, 27.80959, 27.78515, 27.76055, 27.73579, 27.71087, 27.68579, 
    27.66055, 27.63515, 27.60959, 27.58388, 27.558, 27.53197, 27.50578, 
    27.47943, 27.45292, 27.42625, 27.39943, 27.37245, 27.34531, 27.31801, 
    27.29056, 27.26295, 27.23519, 27.20727, 27.1792, 27.15096, 27.12258, 
    27.09403, 27.06534,
  23.85844, 23.90055, 23.94254, 23.98438, 24.0261, 24.06769, 24.10914, 
    24.15045, 24.19164, 24.23268, 24.2736, 24.31437, 24.35502, 24.39553, 
    24.4359, 24.47614, 24.51624, 24.5562, 24.59603, 24.63572, 24.67528, 
    24.71469, 24.75397, 24.79311, 24.83212, 24.87098, 24.90971, 24.9483, 
    24.98674, 25.02505, 25.06322, 25.10125, 25.13914, 25.17689, 25.21449, 
    25.25196, 25.28929, 25.32647, 25.36351, 25.40042, 25.43717, 25.47379, 
    25.51026, 25.54659, 25.58278, 25.61882, 25.65472, 25.69048, 25.72609, 
    25.76156, 25.79688, 25.83206, 25.86709, 25.90198, 25.93672, 25.97132, 
    26.00577, 26.04007, 26.07422, 26.10823, 26.1421, 26.17581, 26.20938, 
    26.2428, 26.27607, 26.30919, 26.34217, 26.37499, 26.40767, 26.4402, 
    26.47258, 26.5048, 26.53688, 26.56881, 26.60059, 26.63222, 26.66369, 
    26.69502, 26.72619, 26.75721, 26.78808, 26.8188, 26.84937, 26.87978, 
    26.91004, 26.94015, 26.9701, 26.9999, 27.02955, 27.05904, 27.08838, 
    27.11757, 27.1466, 27.17547, 27.2042, 27.23276, 27.26117, 27.28942, 
    27.31752, 27.34547, 27.37325, 27.40088, 27.42836, 27.45567, 27.48283, 
    27.50983, 27.53668, 27.56336, 27.58989, 27.61626, 27.64248, 27.66853, 
    27.69443, 27.72016, 27.74574, 27.77115, 27.79641, 27.82151, 27.84645, 
    27.87123, 27.89584, 27.9203, 27.9446, 27.96873, 27.99271, 28.01652, 
    28.04017, 28.06366, 28.08699, 28.11015, 28.13316, 28.156, 28.17867, 
    28.20119, 28.22354, 28.24573, 28.26776, 28.28962, 28.31132, 28.33285, 
    28.35422, 28.37543, 28.39647, 28.41735, 28.43806, 28.4586, 28.47899, 
    28.4992, 28.51925, 28.53914, 28.55886, 28.57841, 28.5978, 28.61702, 
    28.63608, 28.65497, 28.67369, 28.69224, 28.71063, 28.72885, 28.74691, 
    28.76479, 28.78251, 28.80006, 28.81744, 28.83466, 28.8517, 28.86858, 
    28.88529, 28.90183, 28.9182, 28.9344, 28.95044, 28.9663, 28.98199, 
    28.99752, 29.01287, 29.02806, 29.04308, 29.05792, 29.0726, 29.0871, 
    29.10144, 29.1156, 29.1296, 29.14342, 29.15707, 29.17055, 29.18386, 
    29.197, 29.20997, 29.22276, 29.23539, 29.24784, 29.26012, 29.27223, 
    29.28417, 29.29593, 29.30753, 29.31894, 29.33019, 29.34127, 29.35217, 
    29.3629, 29.37346, 29.38384, 29.39405, 29.40409, 29.41396, 29.42365, 
    29.43317, 29.44251, 29.45168, 29.46068, 29.46951, 29.47816, 29.48663, 
    29.49494, 29.50307, 29.51102, 29.5188, 29.52641, 29.53384, 29.5411, 
    29.54818, 29.55509, 29.56182, 29.56839, 29.57477, 29.58098, 29.58702, 
    29.59288, 29.59857, 29.60408, 29.60942, 29.61458, 29.61956, 29.62438, 
    29.62901, 29.63347, 29.63776, 29.64187, 29.64581, 29.64957, 29.65315, 
    29.65656, 29.6598, 29.66286, 29.66574, 29.66845, 29.67098, 29.67334, 
    29.67552, 29.67752, 29.67936, 29.68101, 29.68249, 29.68379, 29.68492, 
    29.68587, 29.68665, 29.68725, 29.68768, 29.68793, 29.688, 29.6879, 
    29.68762, 29.68717, 29.68654, 29.68573, 29.68475, 29.6836, 29.68227, 
    29.68076, 29.67908, 29.67722, 29.67519, 29.67298, 29.67059, 29.66803, 
    29.66529, 29.66238, 29.6593, 29.65603, 29.6526, 29.64898, 29.6452, 
    29.64123, 29.63709, 29.63278, 29.62829, 29.62363, 29.61879, 29.61377, 
    29.60858, 29.60322, 29.59768, 29.59196, 29.58607, 29.58001, 29.57377, 
    29.56736, 29.56077, 29.55401, 29.54707, 29.53996, 29.53268, 29.52522, 
    29.51758, 29.50977, 29.50179, 29.49364, 29.4853, 29.4768, 29.46812, 
    29.45927, 29.45024, 29.44105, 29.43167, 29.42213, 29.41241, 29.40252, 
    29.39245, 29.38221, 29.3718, 29.36122, 29.35046, 29.33953, 29.32843, 
    29.31715, 29.3057, 29.29408, 29.28229, 29.27033, 29.25819, 29.24588, 
    29.2334, 29.22075, 29.20793, 29.19493, 29.18177, 29.16843, 29.15492, 
    29.14124, 29.12739, 29.11337, 29.09918, 29.08482, 29.07029, 29.05559, 
    29.04071, 29.02567, 29.01046, 28.99508, 28.97952, 28.9638, 28.94791, 
    28.93185, 28.91562, 28.89922, 28.88266, 28.86592, 28.84902, 28.83194, 
    28.8147, 28.79729, 28.77972, 28.76197, 28.74406, 28.72598, 28.70774, 
    28.68932, 28.67074, 28.65199, 28.63308, 28.61399, 28.59475, 28.57533, 
    28.55575, 28.53601, 28.51609, 28.49602, 28.47577, 28.45537, 28.43479, 
    28.41405, 28.39315, 28.37208, 28.35085, 28.32945, 28.30789, 28.28617, 
    28.26428, 28.24223, 28.22002, 28.19764, 28.1751, 28.15239, 28.12953, 
    28.1065, 28.08331, 28.05995, 28.03644, 28.01276, 27.98892, 27.96493, 
    27.94076, 27.91644, 27.89196, 27.86732, 27.84251, 27.81755, 27.79243, 
    27.76715, 27.7417, 27.7161, 27.69034, 27.66442, 27.63834, 27.6121, 
    27.58571, 27.55915, 27.53244, 27.50557, 27.47855, 27.45136, 27.42402, 
    27.39652, 27.36887, 27.34106, 27.31309, 27.28497, 27.25669, 27.22825, 
    27.19966, 27.17092,
  23.95871, 24.00089, 24.04294, 24.08485, 24.12663, 24.16828, 24.20979, 
    24.25117, 24.29242, 24.33353, 24.37451, 24.41535, 24.45605, 24.49662, 
    24.53706, 24.57736, 24.61752, 24.65755, 24.69744, 24.73719, 24.77681, 
    24.81628, 24.85563, 24.89483, 24.93389, 24.97282, 25.0116, 25.05025, 
    25.08876, 25.12713, 25.16536, 25.20345, 25.2414, 25.2792, 25.31687, 
    25.3544, 25.39178, 25.42902, 25.46613, 25.50308, 25.5399, 25.57658, 
    25.61311, 25.6495, 25.68574, 25.72184, 25.7578, 25.79361, 25.82928, 
    25.86481, 25.90019, 25.93542, 25.97051, 26.00545, 26.04025, 26.0749, 
    26.10941, 26.14377, 26.17798, 26.21204, 26.24596, 26.27973, 26.31335, 
    26.34683, 26.38015, 26.41333, 26.44636, 26.47924, 26.51197, 26.54455, 
    26.57698, 26.60926, 26.6414, 26.67338, 26.70521, 26.73689, 26.76841, 
    26.79979, 26.83102, 26.86209, 26.89301, 26.92378, 26.9544, 26.98486, 
    27.01517, 27.04533, 27.07533, 27.10518, 27.13488, 27.16442, 27.19381, 
    27.22305, 27.25213, 27.28105, 27.30982, 27.33843, 27.36689, 27.3952, 
    27.42334, 27.45133, 27.47917, 27.50684, 27.53436, 27.56173, 27.58893, 
    27.61598, 27.64287, 27.6696, 27.69618, 27.72259, 27.74885, 27.77495, 
    27.80089, 27.82667, 27.85229, 27.87775, 27.90305, 27.92819, 27.95317, 
    27.97799, 28.00265, 28.02715, 28.05149, 28.07567, 28.09968, 28.12354, 
    28.14723, 28.17076, 28.19413, 28.21733, 28.24038, 28.26326, 28.28597, 
    28.30853, 28.33092, 28.35315, 28.37521, 28.39711, 28.41885, 28.44042, 
    28.46183, 28.48307, 28.50415, 28.52506, 28.54581, 28.56639, 28.58681, 
    28.60707, 28.62715, 28.64707, 28.66683, 28.68641, 28.70584, 28.72509, 
    28.74418, 28.7631, 28.78186, 28.80045, 28.81887, 28.83712, 28.85521, 
    28.87312, 28.89087, 28.90845, 28.92587, 28.94311, 28.96019, 28.9771, 
    28.99384, 29.0104, 29.02681, 29.04304, 29.0591, 29.07499, 29.09071, 
    29.10627, 29.12165, 29.13686, 29.15191, 29.16678, 29.18148, 29.19601, 
    29.21037, 29.22456, 29.23858, 29.25243, 29.26611, 29.27961, 29.29295, 
    29.30611, 29.3191, 29.33192, 29.34456, 29.35704, 29.36934, 29.38147, 
    29.39343, 29.40522, 29.41683, 29.42827, 29.43954, 29.45064, 29.46156, 
    29.47231, 29.48288, 29.49329, 29.50352, 29.51357, 29.52346, 29.53316, 
    29.5427, 29.55206, 29.56125, 29.57027, 29.57911, 29.58777, 29.59627, 
    29.60458, 29.61273, 29.6207, 29.62849, 29.63611, 29.64356, 29.65083, 
    29.65793, 29.66485, 29.67159, 29.67817, 29.68456, 29.69079, 29.69683, 
    29.70271, 29.7084, 29.71392, 29.71927, 29.72444, 29.72944, 29.73426, 
    29.7389, 29.74337, 29.74767, 29.75179, 29.75573, 29.7595, 29.76309, 
    29.7665, 29.76974, 29.77281, 29.7757, 29.77841, 29.78095, 29.78331, 
    29.7855, 29.78751, 29.78934, 29.791, 29.79248, 29.79379, 29.79491, 
    29.79587, 29.79665, 29.79725, 29.79768, 29.79793, 29.798, 29.7979, 
    29.79762, 29.79716, 29.79654, 29.79573, 29.79475, 29.79359, 29.79226, 
    29.79075, 29.78906, 29.7872, 29.78516, 29.78295, 29.78056, 29.77799, 
    29.77525, 29.77234, 29.76925, 29.76598, 29.76253, 29.75891, 29.75512, 
    29.75115, 29.747, 29.74268, 29.73818, 29.73351, 29.72866, 29.72364, 
    29.71844, 29.71306, 29.70751, 29.70179, 29.69589, 29.68981, 29.68356, 
    29.67714, 29.67054, 29.66376, 29.65681, 29.64969, 29.64239, 29.63492, 
    29.62727, 29.61945, 29.61145, 29.60328, 29.59493, 29.58641, 29.57772, 
    29.56885, 29.55981, 29.55059, 29.5412, 29.53164, 29.5219, 29.51199, 
    29.50191, 29.49165, 29.48122, 29.47062, 29.45984, 29.44889, 29.43777, 
    29.42647, 29.415, 29.40336, 29.39155, 29.37957, 29.36741, 29.35508, 
    29.34258, 29.3299, 29.31705, 29.30404, 29.29085, 29.27749, 29.26395, 
    29.25025, 29.23638, 29.22233, 29.20811, 29.19372, 29.17916, 29.16444, 
    29.14954, 29.13447, 29.11923, 29.10382, 29.08824, 29.07249, 29.05657, 
    29.04048, 29.02422, 29.0078, 28.9912, 28.97443, 28.9575, 28.9404, 
    28.92312, 28.90568, 28.88808, 28.8703, 28.85236, 28.83424, 28.81596, 
    28.79752, 28.7789, 28.76012, 28.74117, 28.72206, 28.70278, 28.68333, 
    28.66371, 28.64393, 28.62399, 28.60387, 28.58359, 28.56315, 28.54254, 
    28.52176, 28.50083, 28.47972, 28.45845, 28.43702, 28.41542, 28.39366, 
    28.37173, 28.34964, 28.32739, 28.30497, 28.28239, 28.25965, 28.23674, 
    28.21367, 28.19044, 28.16705, 28.14349, 28.11977, 28.09589, 28.07185, 
    28.04765, 28.02329, 27.99876, 27.97408, 27.94923, 27.92422, 27.89906, 
    27.87373, 27.84824, 27.8226, 27.79679, 27.77083, 27.74471, 27.71842, 
    27.69198, 27.66538, 27.63863, 27.61171, 27.58464, 27.55741, 27.53002, 
    27.50248, 27.47477, 27.44691, 27.4189, 27.39073, 27.3624, 27.33392, 
    27.30528, 27.27649,
  24.05898, 24.10122, 24.14333, 24.1853, 24.22715, 24.26886, 24.31043, 
    24.35188, 24.39319, 24.43436, 24.4754, 24.5163, 24.55707, 24.59771, 
    24.6382, 24.67856, 24.71879, 24.75888, 24.79883, 24.83864, 24.87832, 
    24.91786, 24.95726, 24.99653, 25.03565, 25.07464, 25.11349, 25.15219, 
    25.19076, 25.22919, 25.26748, 25.30563, 25.34364, 25.38151, 25.41923, 
    25.45682, 25.49426, 25.53156, 25.56872, 25.60574, 25.64262, 25.67935, 
    25.71594, 25.75239, 25.78869, 25.82485, 25.86086, 25.89673, 25.93246, 
    25.96804, 26.00348, 26.03877, 26.07392, 26.10892, 26.14377, 26.17848, 
    26.21304, 26.24745, 26.28172, 26.31584, 26.34981, 26.38364, 26.41732, 
    26.45085, 26.48423, 26.51746, 26.55054, 26.58347, 26.61626, 26.64889, 
    26.68138, 26.71371, 26.7459, 26.77793, 26.80981, 26.84155, 26.87313, 
    26.90455, 26.93583, 26.96696, 26.99793, 27.02875, 27.05942, 27.08993, 
    27.12029, 27.1505, 27.18056, 27.21046, 27.24021, 27.2698, 27.29924, 
    27.32852, 27.35765, 27.38662, 27.41544, 27.4441, 27.47261, 27.50096, 
    27.52915, 27.55719, 27.58507, 27.61279, 27.64036, 27.66777, 27.69502, 
    27.72212, 27.74905, 27.77583, 27.80245, 27.82891, 27.85521, 27.88136, 
    27.90734, 27.93316, 27.95883, 27.98433, 28.00968, 28.03486, 28.05989, 
    28.08475, 28.10945, 28.134, 28.15837, 28.18259, 28.20665, 28.23055, 
    28.25428, 28.27785, 28.30126, 28.3245, 28.34759, 28.37051, 28.39327, 
    28.41586, 28.43829, 28.46056, 28.48266, 28.5046, 28.52637, 28.54798, 
    28.56943, 28.59071, 28.61182, 28.63277, 28.65356, 28.67418, 28.69463, 
    28.71492, 28.73504, 28.755, 28.77479, 28.79441, 28.81387, 28.83316, 
    28.85228, 28.87124, 28.89002, 28.90865, 28.9271, 28.94538, 28.9635, 
    28.98145, 28.99923, 29.01685, 29.03429, 29.05157, 29.06867, 29.08561, 
    29.10238, 29.11898, 29.13541, 29.15167, 29.16776, 29.18368, 29.19943, 
    29.21501, 29.23042, 29.24566, 29.26073, 29.27563, 29.29036, 29.30492, 
    29.3193, 29.33352, 29.34756, 29.36144, 29.37514, 29.38867, 29.40203, 
    29.41521, 29.42823, 29.44107, 29.45374, 29.46624, 29.47856, 29.49071, 
    29.50269, 29.5145, 29.52614, 29.5376, 29.54889, 29.56, 29.57094, 
    29.58171, 29.59231, 29.60273, 29.61298, 29.62305, 29.63295, 29.64268, 
    29.65224, 29.66161, 29.67082, 29.67985, 29.68871, 29.69739, 29.7059, 
    29.71423, 29.72239, 29.73037, 29.73818, 29.74582, 29.75327, 29.76056, 
    29.76767, 29.7746, 29.78136, 29.78795, 29.79436, 29.80059, 29.80665, 
    29.81253, 29.81824, 29.82377, 29.82913, 29.83431, 29.83931, 29.84414, 
    29.84879, 29.85327, 29.85758, 29.8617, 29.86565, 29.86943, 29.87302, 
    29.87645, 29.87969, 29.88276, 29.88566, 29.88838, 29.89092, 29.89328, 
    29.89547, 29.89749, 29.89932, 29.90098, 29.90247, 29.90378, 29.90491, 
    29.90586, 29.90664, 29.90725, 29.90767, 29.90792, 29.908, 29.9079, 
    29.90762, 29.90716, 29.90653, 29.90573, 29.90474, 29.90358, 29.90225, 
    29.90073, 29.89904, 29.89718, 29.89514, 29.89292, 29.89053, 29.88796, 
    29.88521, 29.88229, 29.87919, 29.87592, 29.87247, 29.86884, 29.86504, 
    29.86106, 29.85691, 29.85258, 29.84807, 29.84339, 29.83853, 29.8335, 
    29.82829, 29.82291, 29.81735, 29.81161, 29.8057, 29.79962, 29.79335, 
    29.78692, 29.78031, 29.77352, 29.76656, 29.75942, 29.75211, 29.74462, 
    29.73696, 29.72912, 29.72111, 29.71292, 29.70456, 29.69603, 29.68732, 
    29.67843, 29.66937, 29.66014, 29.65074, 29.64116, 29.6314, 29.62147, 
    29.61137, 29.60109, 29.59064, 29.58002, 29.56923, 29.55825, 29.54711, 
    29.5358, 29.52431, 29.51265, 29.50081, 29.4888, 29.47662, 29.46427, 
    29.45175, 29.43905, 29.42618, 29.41314, 29.39992, 29.38654, 29.37298, 
    29.35925, 29.34535, 29.33128, 29.31704, 29.30263, 29.28804, 29.27328, 
    29.25836, 29.24326, 29.22799, 29.21256, 29.19695, 29.18117, 29.16522, 
    29.14911, 29.13282, 29.11636, 29.09974, 29.08294, 29.06598, 29.04884, 
    29.03154, 29.01407, 28.99643, 28.97862, 28.96065, 28.9425, 28.92419, 
    28.90571, 28.88706, 28.86825, 28.84927, 28.83012, 28.8108, 28.79132, 
    28.77167, 28.75185, 28.73187, 28.71172, 28.69141, 28.67093, 28.65028, 
    28.62947, 28.6085, 28.58735, 28.56605, 28.54457, 28.52294, 28.50114, 
    28.47917, 28.45705, 28.43475, 28.4123, 28.38968, 28.36689, 28.34395, 
    28.32084, 28.29757, 28.27413, 28.25054, 28.22678, 28.20286, 28.17877, 
    28.15453, 28.13012, 28.10556, 28.08083, 28.05594, 28.03089, 28.00568, 
    27.98031, 27.95478, 27.92909, 27.90324, 27.87723, 27.85106, 27.82474, 
    27.79825, 27.77161, 27.7448, 27.71784, 27.69072, 27.66345, 27.63601, 
    27.60842, 27.58067, 27.55276, 27.5247, 27.49648, 27.46811, 27.43958, 
    27.41089, 27.38205,
  24.15922, 24.20152, 24.2437, 24.28574, 24.32765, 24.36942, 24.41106, 
    24.45257, 24.49394, 24.53518, 24.57628, 24.61724, 24.65808, 24.69877, 
    24.73933, 24.77976, 24.82004, 24.86019, 24.90021, 24.94008, 24.97982, 
    25.01942, 25.05889, 25.09821, 25.1374, 25.17644, 25.21535, 25.25412, 
    25.29275, 25.33124, 25.36959, 25.4078, 25.44587, 25.48379, 25.52158, 
    25.55923, 25.59673, 25.63409, 25.67131, 25.70839, 25.74532, 25.78211, 
    25.81876, 25.85526, 25.89162, 25.92784, 25.96391, 25.99984, 26.03563, 
    26.07127, 26.10676, 26.14211, 26.17731, 26.21237, 26.24728, 26.28204, 
    26.31666, 26.35113, 26.38545, 26.41963, 26.45366, 26.48754, 26.52127, 
    26.55485, 26.58829, 26.62157, 26.65471, 26.6877, 26.72054, 26.75323, 
    26.78576, 26.81815, 26.85039, 26.88247, 26.91441, 26.9462, 26.97783, 
    27.00931, 27.04064, 27.07182, 27.10284, 27.13371, 27.16443, 27.195, 
    27.22541, 27.25567, 27.28577, 27.31572, 27.34552, 27.37516, 27.40465, 
    27.43398, 27.46316, 27.49218, 27.52105, 27.54976, 27.57831, 27.60671, 
    27.63495, 27.66304, 27.69097, 27.71874, 27.74635, 27.77381, 27.80111, 
    27.82825, 27.85523, 27.88205, 27.90872, 27.93522, 27.96157, 27.98776, 
    28.01379, 28.03966, 28.06536, 28.09091, 28.1163, 28.14153, 28.1666, 
    28.1915, 28.21625, 28.24083, 28.26525, 28.28952, 28.31361, 28.33755, 
    28.36133, 28.38494, 28.40839, 28.43167, 28.4548, 28.47776, 28.50056, 
    28.52319, 28.54566, 28.56796, 28.5901, 28.61208, 28.63389, 28.65554, 
    28.67702, 28.69834, 28.71949, 28.74048, 28.7613, 28.78196, 28.80245, 
    28.82277, 28.84293, 28.86292, 28.88275, 28.9024, 28.9219, 28.94122, 
    28.96038, 28.97936, 28.99819, 29.01684, 29.03533, 29.05364, 29.07179, 
    29.08978, 29.10759, 29.12523, 29.14271, 29.16001, 29.17715, 29.19412, 
    29.21092, 29.22755, 29.24401, 29.2603, 29.27641, 29.29236, 29.30814, 
    29.32375, 29.33919, 29.35446, 29.36956, 29.38448, 29.39924, 29.41382, 
    29.42823, 29.44247, 29.45654, 29.47044, 29.48417, 29.49772, 29.5111, 
    29.52431, 29.53735, 29.55022, 29.56291, 29.57543, 29.58778, 29.59995, 
    29.61195, 29.62378, 29.63544, 29.64692, 29.65823, 29.66937, 29.68033, 
    29.69112, 29.70173, 29.71217, 29.72244, 29.73253, 29.74245, 29.7522, 
    29.76177, 29.77116, 29.78038, 29.78943, 29.79831, 29.807, 29.81553, 
    29.82387, 29.83205, 29.84005, 29.84787, 29.85552, 29.86299, 29.87029, 
    29.87741, 29.88436, 29.89113, 29.89773, 29.90415, 29.91039, 29.91646, 
    29.92236, 29.92807, 29.93362, 29.93898, 29.94417, 29.94919, 29.95403, 
    29.95869, 29.96317, 29.96748, 29.97162, 29.97557, 29.97935, 29.98296, 
    29.98639, 29.98964, 29.99272, 29.99562, 29.99834, 30.00089, 30.00326, 
    30.00545, 30.00747, 30.00931, 30.01097, 30.01246, 30.01377, 30.0149, 
    30.01586, 30.01664, 30.01725, 30.01767, 30.01793, 30.018, 30.0179, 
    30.01762, 30.01716, 30.01653, 30.01572, 30.01474, 30.01357, 30.01224, 
    30.01072, 30.00903, 30.00716, 30.00512, 30.00289, 30.0005, 29.99792, 
    29.99517, 29.99224, 29.98914, 29.98586, 29.9824, 29.97877, 29.97496, 
    29.97097, 29.96681, 29.96247, 29.95796, 29.95327, 29.9484, 29.94336, 
    29.93814, 29.93275, 29.92718, 29.92144, 29.91551, 29.90942, 29.90314, 
    29.8967, 29.89007, 29.88327, 29.8763, 29.86915, 29.86182, 29.85432, 
    29.84664, 29.83879, 29.83077, 29.82257, 29.81419, 29.80564, 29.79691, 
    29.78801, 29.77894, 29.76969, 29.76027, 29.75067, 29.74089, 29.73095, 
    29.72083, 29.71053, 29.70006, 29.68942, 29.67861, 29.66762, 29.65645, 
    29.64512, 29.63361, 29.62192, 29.61007, 29.59804, 29.58584, 29.57346, 
    29.56091, 29.54819, 29.5353, 29.52224, 29.509, 29.49559, 29.48201, 
    29.46825, 29.45433, 29.44023, 29.42596, 29.41153, 29.39691, 29.38213, 
    29.36718, 29.35205, 29.33676, 29.32129, 29.30566, 29.28985, 29.27388, 
    29.25773, 29.24142, 29.22493, 29.20827, 29.19145, 29.17445, 29.15729, 
    29.13996, 29.12245, 29.10478, 29.08694, 29.06893, 29.05076, 29.03241, 
    29.0139, 28.99522, 28.97637, 28.95736, 28.93817, 28.91882, 28.89931, 
    28.87962, 28.85977, 28.83975, 28.81957, 28.79922, 28.7787, 28.75802, 
    28.73717, 28.71616, 28.69498, 28.67364, 28.65213, 28.63045, 28.60862, 
    28.58661, 28.56445, 28.54211, 28.51962, 28.49696, 28.47414, 28.45115, 
    28.428, 28.40469, 28.38121, 28.35758, 28.33378, 28.30981, 28.28569, 
    28.2614, 28.23695, 28.21235, 28.18757, 28.16264, 28.13755, 28.1123, 
    28.08688, 28.06131, 28.03557, 28.00968, 27.98363, 27.95741, 27.93104, 
    27.90451, 27.87782, 27.85097, 27.82397, 27.7968, 27.76948, 27.74199, 
    27.71436, 27.68656, 27.65861, 27.6305, 27.60223, 27.57381, 27.54523, 
    27.51649, 27.4876,
  24.25945, 24.30182, 24.34406, 24.38616, 24.42813, 24.46997, 24.51167, 
    24.55324, 24.59468, 24.63598, 24.67714, 24.71817, 24.75907, 24.79982, 
    24.84045, 24.88093, 24.92128, 24.96149, 25.00157, 25.04151, 25.08131, 
    25.12097, 25.16049, 25.19988, 25.23913, 25.27824, 25.31721, 25.35604, 
    25.39472, 25.43327, 25.47168, 25.50995, 25.54808, 25.58607, 25.62391, 
    25.66162, 25.69918, 25.7366, 25.77388, 25.81102, 25.84801, 25.88486, 
    25.92157, 25.95813, 25.99455, 26.03082, 26.06695, 26.10294, 26.13878, 
    26.17448, 26.21003, 26.24543, 26.28069, 26.31581, 26.35077, 26.38559, 
    26.42027, 26.45479, 26.48917, 26.5234, 26.55749, 26.59142, 26.62521, 
    26.65885, 26.69234, 26.72568, 26.75887, 26.79191, 26.8248, 26.85755, 
    26.89014, 26.92258, 26.95487, 26.98701, 27.019, 27.05083, 27.08252, 
    27.11405, 27.14543, 27.17666, 27.20774, 27.23866, 27.26943, 27.30005, 
    27.33051, 27.36082, 27.39098, 27.42098, 27.45083, 27.48052, 27.51006, 
    27.53944, 27.56866, 27.59773, 27.62665, 27.65541, 27.68401, 27.71246, 
    27.74075, 27.76888, 27.79686, 27.82467, 27.85233, 27.87984, 27.90718, 
    27.93437, 27.9614, 27.98827, 28.01498, 28.04153, 28.06792, 28.09415, 
    28.12023, 28.14614, 28.17189, 28.19748, 28.22292, 28.24819, 28.2733, 
    28.29825, 28.32304, 28.34766, 28.37213, 28.39643, 28.42057, 28.44455, 
    28.46836, 28.49202, 28.51551, 28.53884, 28.562, 28.585, 28.60784, 
    28.63051, 28.65302, 28.67536, 28.69754, 28.71956, 28.74141, 28.76309, 
    28.78461, 28.80597, 28.82716, 28.84818, 28.86904, 28.88974, 28.91026, 
    28.93062, 28.95082, 28.97084, 28.9907, 29.01039, 29.02992, 29.04928, 
    29.06847, 29.08749, 29.10634, 29.12503, 29.14355, 29.1619, 29.18008, 
    29.1981, 29.21594, 29.23362, 29.25112, 29.26846, 29.28563, 29.30263, 
    29.31945, 29.33611, 29.3526, 29.36892, 29.38507, 29.40105, 29.41685, 
    29.43249, 29.44796, 29.46325, 29.47838, 29.49333, 29.50811, 29.52272, 
    29.53716, 29.55143, 29.56552, 29.57944, 29.59319, 29.60677, 29.62018, 
    29.63341, 29.64647, 29.65936, 29.67208, 29.68462, 29.69699, 29.70919, 
    29.72121, 29.73306, 29.74474, 29.75624, 29.76757, 29.77873, 29.78971, 
    29.80052, 29.81115, 29.82161, 29.8319, 29.84201, 29.85195, 29.86171, 
    29.8713, 29.88071, 29.88995, 29.89901, 29.9079, 29.91662, 29.92516, 
    29.93352, 29.94171, 29.94972, 29.95756, 29.96522, 29.97271, 29.98002, 
    29.98715, 29.99411, 30.0009, 30.00751, 30.01394, 30.0202, 30.02628, 
    30.03218, 30.03791, 30.04346, 30.04884, 30.05404, 30.05906, 30.06391, 
    30.06858, 30.07307, 30.07739, 30.08153, 30.0855, 30.08928, 30.0929, 
    30.09633, 30.09959, 30.10267, 30.10558, 30.1083, 30.11086, 30.11323, 
    30.11543, 30.11745, 30.11929, 30.12096, 30.12245, 30.12376, 30.1249, 
    30.12586, 30.12664, 30.12724, 30.12767, 30.12793, 30.128, 30.1279, 
    30.12762, 30.12716, 30.12653, 30.12572, 30.12473, 30.12357, 30.12222, 
    30.12071, 30.11901, 30.11714, 30.11509, 30.11287, 30.11046, 30.10788, 
    30.10513, 30.1022, 30.09909, 30.0958, 30.09234, 30.0887, 30.08488, 
    30.08089, 30.07672, 30.07237, 30.06785, 30.06315, 30.05828, 30.05323, 
    30.048, 30.04259, 30.03701, 30.03126, 30.02533, 30.01922, 30.01293, 
    30.00647, 29.99984, 29.99302, 29.98604, 29.97887, 29.97153, 29.96402, 
    29.95633, 29.94846, 29.94042, 29.93221, 29.92382, 29.91525, 29.90651, 
    29.89759, 29.8885, 29.87923, 29.86979, 29.86018, 29.85039, 29.84042, 
    29.83028, 29.81997, 29.80948, 29.79882, 29.78798, 29.77698, 29.76579, 
    29.75443, 29.7429, 29.7312, 29.71932, 29.70727, 29.69505, 29.68265, 
    29.67008, 29.65734, 29.64442, 29.63133, 29.61807, 29.60464, 29.59103, 
    29.57725, 29.5633, 29.54918, 29.53489, 29.52042, 29.50578, 29.49098, 
    29.476, 29.46085, 29.44552, 29.43003, 29.41437, 29.39853, 29.38253, 
    29.36635, 29.35001, 29.33349, 29.3168, 29.29995, 29.28292, 29.26573, 
    29.24837, 29.23083, 29.21313, 29.19526, 29.17722, 29.15901, 29.14063, 
    29.12209, 29.10337, 29.08449, 29.06544, 29.04623, 29.02684, 29.00729, 
    28.98757, 28.96768, 28.94763, 28.92741, 28.90703, 28.88647, 28.86576, 
    28.84487, 28.82382, 28.8026, 28.78122, 28.75968, 28.73796, 28.71609, 
    28.69405, 28.67184, 28.64947, 28.62693, 28.60423, 28.58137, 28.55835, 
    28.53516, 28.5118, 28.48829, 28.46461, 28.44077, 28.41676, 28.3926, 
    28.36827, 28.34378, 28.31913, 28.29431, 28.26934, 28.2442, 28.21891, 
    28.19345, 28.16783, 28.14205, 28.11611, 28.09002, 28.06376, 28.03734, 
    28.01076, 27.98403, 27.95713, 27.93008, 27.90287, 27.8755, 27.84797, 
    27.82028, 27.79244, 27.76444, 27.73628, 27.70797, 27.6795, 27.65087, 
    27.62209, 27.59315,
  24.35966, 24.40209, 24.4444, 24.48656, 24.5286, 24.5705, 24.61227, 24.6539, 
    24.6954, 24.73676, 24.77799, 24.81908, 24.86004, 24.90086, 24.94154, 
    24.98209, 25.0225, 25.06278, 25.10292, 25.14292, 25.18278, 25.2225, 
    25.26209, 25.30154, 25.34084, 25.38001, 25.41904, 25.45793, 25.49669, 
    25.5353, 25.57376, 25.61209, 25.65028, 25.68833, 25.72623, 25.764, 
    25.80162, 25.8391, 25.87644, 25.91363, 25.95069, 25.98759, 26.02436, 
    26.06098, 26.09746, 26.13379, 26.16998, 26.20602, 26.24192, 26.27768, 
    26.31328, 26.34875, 26.38406, 26.41923, 26.45426, 26.48913, 26.52386, 
    26.55844, 26.59288, 26.62717, 26.6613, 26.6953, 26.72914, 26.76283, 
    26.79638, 26.82977, 26.86302, 26.89611, 26.92906, 26.96186, 26.9945, 
    27.027, 27.05934, 27.09153, 27.12357, 27.15546, 27.1872, 27.21879, 
    27.25022, 27.2815, 27.31263, 27.3436, 27.37443, 27.40509, 27.43561, 
    27.46597, 27.49617, 27.52623, 27.55612, 27.58587, 27.61545, 27.64488, 
    27.67416, 27.70328, 27.73224, 27.76105, 27.7897, 27.8182, 27.84653, 
    27.87471, 27.90274, 27.9306, 27.95831, 27.98586, 28.01325, 28.04048, 
    28.06756, 28.09447, 28.12123, 28.14783, 28.17426, 28.20054, 28.22666, 
    28.25262, 28.27841, 28.30405, 28.32953, 28.35484, 28.38, 28.40499, 
    28.42982, 28.45449, 28.47899, 28.50334, 28.52752, 28.55154, 28.5754, 
    28.59909, 28.62263, 28.64599, 28.6692, 28.69224, 28.71511, 28.73783, 
    28.76037, 28.78276, 28.80498, 28.82703, 28.84892, 28.87064, 28.8922, 
    28.9136, 28.93482, 28.95588, 28.97678, 28.99751, 29.01807, 29.03846, 
    29.05869, 29.07875, 29.09865, 29.11838, 29.13794, 29.15733, 29.17655, 
    29.19561, 29.2145, 29.23322, 29.25177, 29.27015, 29.28837, 29.30641, 
    29.32429, 29.342, 29.35954, 29.3769, 29.3941, 29.41113, 29.42799, 
    29.44468, 29.46119, 29.47754, 29.49372, 29.50973, 29.52556, 29.54123, 
    29.55672, 29.57204, 29.5872, 29.60218, 29.61698, 29.63162, 29.64608, 
    29.66038, 29.6745, 29.68845, 29.70222, 29.71582, 29.72925, 29.74251, 
    29.7556, 29.76851, 29.78125, 29.79381, 29.80621, 29.81842, 29.83047, 
    29.84234, 29.85404, 29.86556, 29.87691, 29.88809, 29.89909, 29.90992, 
    29.92057, 29.93105, 29.94136, 29.95149, 29.96144, 29.97122, 29.98083, 
    29.99026, 29.99951, 30.00859, 30.0175, 30.02623, 30.03478, 30.04316, 
    30.05136, 30.05939, 30.06725, 30.07492, 30.08242, 30.08975, 30.0969, 
    30.10387, 30.11066, 30.11728, 30.12373, 30.13, 30.13609, 30.142, 
    30.14774, 30.15331, 30.15869, 30.1639, 30.16893, 30.17379, 30.17847, 
    30.18297, 30.1873, 30.19145, 30.19542, 30.19921, 30.20283, 30.20627, 
    30.20954, 30.21262, 30.21553, 30.21827, 30.22082, 30.2232, 30.2254, 
    30.22743, 30.22927, 30.23095, 30.23244, 30.23375, 30.23489, 30.23585, 
    30.23664, 30.23724, 30.23767, 30.23792, 30.238, 30.2379, 30.23762, 
    30.23716, 30.23652, 30.23571, 30.23472, 30.23356, 30.23221, 30.23069, 
    30.22899, 30.22712, 30.22507, 30.22284, 30.22043, 30.21785, 30.21509, 
    30.21215, 30.20903, 30.20574, 30.20227, 30.19863, 30.1948, 30.1908, 
    30.18662, 30.18227, 30.17774, 30.17303, 30.16815, 30.16309, 30.15785, 
    30.15244, 30.14685, 30.14108, 30.13514, 30.12902, 30.12272, 30.11625, 
    30.1096, 30.10278, 30.09578, 30.0886, 30.08125, 30.07372, 30.06602, 
    30.05814, 30.05008, 30.04185, 30.03344, 30.02486, 30.0161, 30.00717, 
    29.99806, 29.98878, 29.97932, 29.96969, 29.95988, 29.9499, 29.93974, 
    29.92941, 29.9189, 29.90822, 29.89736, 29.88633, 29.87513, 29.86375, 
    29.8522, 29.84048, 29.82858, 29.8165, 29.80426, 29.79184, 29.77925, 
    29.76648, 29.75354, 29.74043, 29.72714, 29.71368, 29.70005, 29.68625, 
    29.67228, 29.65813, 29.64381, 29.62932, 29.61465, 29.59982, 29.58481, 
    29.56963, 29.55428, 29.53876, 29.52307, 29.50721, 29.49117, 29.47497, 
    29.45859, 29.44205, 29.42533, 29.40845, 29.39139, 29.37417, 29.35677, 
    29.33921, 29.32147, 29.30357, 29.2855, 29.26726, 29.24885, 29.23027, 
    29.21152, 29.19261, 29.17352, 29.15427, 29.13485, 29.11527, 29.09551, 
    29.07559, 29.0555, 29.03525, 29.01483, 28.99424, 28.97348, 28.95256, 
    28.93147, 28.91022, 28.8888, 28.86722, 28.84547, 28.82355, 28.80147, 
    28.77923, 28.75682, 28.73424, 28.71151, 28.6886, 28.66554, 28.64231, 
    28.61891, 28.59536, 28.57164, 28.54775, 28.52371, 28.4995, 28.47513, 
    28.4506, 28.4259, 28.40104, 28.37603, 28.35085, 28.32551, 28.30001, 
    28.27435, 28.24852, 28.22254, 28.1964, 28.17009, 28.14363, 28.11701, 
    28.09023, 28.06329, 28.03619, 28.00893, 27.98151, 27.95394, 27.9262, 
    27.89832, 27.87027, 27.84206, 27.8137, 27.78518, 27.7565, 27.72767, 
    27.69868,
  24.45985, 24.50235, 24.54472, 24.58695, 24.62905, 24.67101, 24.71284, 
    24.75454, 24.7961, 24.83753, 24.87882, 24.91998, 24.961, 25.00188, 
    25.04263, 25.08324, 25.12371, 25.16405, 25.20425, 25.24431, 25.28424, 
    25.32402, 25.36367, 25.40318, 25.44255, 25.48178, 25.52087, 25.55982, 
    25.59863, 25.6373, 25.67583, 25.71422, 25.75247, 25.79058, 25.82854, 
    25.86637, 25.90405, 25.94159, 25.97898, 26.01624, 26.05335, 26.09031, 
    26.12714, 26.16382, 26.20036, 26.23675, 26.27299, 26.30909, 26.34505, 
    26.38086, 26.41653, 26.45205, 26.48742, 26.52265, 26.55773, 26.59266, 
    26.62745, 26.66208, 26.69658, 26.73092, 26.76511, 26.79916, 26.83306, 
    26.8668, 26.9004, 26.93386, 26.96716, 27.00031, 27.03331, 27.06615, 
    27.09885, 27.1314, 27.1638, 27.19605, 27.22814, 27.26008, 27.29187, 
    27.32351, 27.355, 27.38633, 27.41751, 27.44854, 27.47941, 27.51013, 
    27.54069, 27.5711, 27.60136, 27.63146, 27.66141, 27.6912, 27.72084, 
    27.75032, 27.77964, 27.80881, 27.83783, 27.86668, 27.89538, 27.92393, 
    27.95231, 27.98054, 28.00861, 28.03652, 28.06428, 28.09187, 28.11931, 
    28.14659, 28.17371, 28.20067, 28.22747, 28.25412, 28.2806, 28.30692, 
    28.33309, 28.35909, 28.38493, 28.41061, 28.43613, 28.46149, 28.48668, 
    28.51172, 28.53659, 28.56131, 28.58586, 28.61024, 28.63447, 28.65853, 
    28.68243, 28.70616, 28.72973, 28.75314, 28.77639, 28.79947, 28.82238, 
    28.84514, 28.86772, 28.89015, 28.91241, 28.9345, 28.95642, 28.97819, 
    28.99978, 29.02121, 29.04248, 29.06358, 29.08451, 29.10527, 29.12587, 
    29.1463, 29.16657, 29.18666, 29.20659, 29.22636, 29.24595, 29.26538, 
    29.28464, 29.30373, 29.32265, 29.3414, 29.35999, 29.3784, 29.39665, 
    29.41473, 29.43264, 29.45037, 29.46794, 29.48534, 29.50257, 29.51963, 
    29.53652, 29.55324, 29.56979, 29.58616, 29.60237, 29.6184, 29.63427, 
    29.64996, 29.66548, 29.68083, 29.69601, 29.71102, 29.72585, 29.74052, 
    29.75501, 29.76933, 29.78347, 29.79744, 29.81124, 29.82487, 29.83833, 
    29.85161, 29.86472, 29.87765, 29.89042, 29.903, 29.91542, 29.92766, 
    29.93973, 29.95162, 29.96334, 29.97488, 29.98625, 29.99745, 30.00847, 
    30.01932, 30.02999, 30.04049, 30.05081, 30.06096, 30.07094, 30.08073, 
    30.09036, 30.0998, 30.10908, 30.11817, 30.12709, 30.13584, 30.14441, 
    30.15281, 30.16102, 30.16907, 30.17693, 30.18462, 30.19214, 30.19947, 
    30.20664, 30.21362, 30.22043, 30.22706, 30.23352, 30.2398, 30.2459, 
    30.25183, 30.25758, 30.26315, 30.26855, 30.27377, 30.27881, 30.28367, 
    30.28836, 30.29287, 30.2972, 30.30136, 30.30534, 30.30914, 30.31277, 
    30.31622, 30.31948, 30.32258, 30.32549, 30.32823, 30.33079, 30.33318, 
    30.33538, 30.33741, 30.33926, 30.34093, 30.34243, 30.34375, 30.34489, 
    30.34585, 30.34663, 30.34724, 30.34767, 30.34793, 30.348, 30.3479, 
    30.34762, 30.34716, 30.34652, 30.34571, 30.34472, 30.34355, 30.3422, 
    30.34068, 30.33898, 30.3371, 30.33504, 30.33281, 30.3304, 30.32781, 
    30.32504, 30.3221, 30.31898, 30.31568, 30.31221, 30.30855, 30.30472, 
    30.30071, 30.29653, 30.29217, 30.28763, 30.28291, 30.27802, 30.27295, 
    30.2677, 30.26228, 30.25668, 30.2509, 30.24495, 30.23882, 30.23251, 
    30.22603, 30.21937, 30.21253, 30.20551, 30.19833, 30.19096, 30.18342, 
    30.1757, 30.1678, 30.15973, 30.15149, 30.14307, 30.13447, 30.1257, 
    30.11675, 30.10762, 30.09832, 30.08885, 30.0792, 30.06937, 30.05937, 
    30.04919, 30.03884, 30.02832, 30.01762, 30.00674, 29.99569, 29.98447, 
    29.97307, 29.9615, 29.94975, 29.93783, 29.92573, 29.91347, 29.90102, 
    29.88841, 29.87562, 29.86266, 29.84952, 29.83621, 29.82273, 29.80907, 
    29.79525, 29.78124, 29.76707, 29.75273, 29.73821, 29.72352, 29.70866, 
    29.69362, 29.67842, 29.66304, 29.64749, 29.63177, 29.61588, 29.59982, 
    29.58358, 29.56718, 29.55061, 29.53386, 29.51694, 29.49986, 29.4826, 
    29.46518, 29.44758, 29.42981, 29.41188, 29.39377, 29.3755, 29.35706, 
    29.33845, 29.31967, 29.30072, 29.2816, 29.26232, 29.24286, 29.22324, 
    29.20345, 29.1835, 29.16337, 29.14308, 29.12262, 29.102, 29.08121, 
    29.06025, 29.03913, 29.01783, 28.99638, 28.97475, 28.95297, 28.93101, 
    28.9089, 28.88661, 28.86416, 28.84155, 28.81877, 28.79583, 28.77272, 
    28.74945, 28.72602, 28.70242, 28.67866, 28.65473, 28.63065, 28.6064, 
    28.58198, 28.55741, 28.53267, 28.50777, 28.48271, 28.45749, 28.4321, 
    28.40656, 28.38085, 28.35498, 28.32896, 28.30277, 28.27642, 28.24991, 
    28.22325, 28.19642, 28.16943, 28.14229, 28.11498, 28.08752, 28.0599, 
    28.03212, 28.00418, 27.97608, 27.94783, 27.91942, 27.89085, 27.86213, 
    27.83325, 27.80421,
  24.56003, 24.6026, 24.64503, 24.68732, 24.72949, 24.77151, 24.81341, 
    24.85517, 24.89679, 24.93828, 24.97964, 25.02086, 25.06194, 25.10289, 
    25.1437, 25.18437, 25.22491, 25.2653, 25.30557, 25.34569, 25.38568, 
    25.42552, 25.46523, 25.5048, 25.54423, 25.58352, 25.62268, 25.66169, 
    25.70056, 25.73929, 25.77788, 25.81633, 25.85464, 25.89281, 25.93084, 
    25.96872, 26.00646, 26.04406, 26.08152, 26.11883, 26.156, 26.19302, 
    26.22991, 26.26665, 26.30324, 26.33969, 26.37599, 26.41215, 26.44817, 
    26.48404, 26.51976, 26.55533, 26.59076, 26.62605, 26.66119, 26.69617, 
    26.73102, 26.76571, 26.80026, 26.83466, 26.86891, 26.90301, 26.93696, 
    26.97077, 27.00442, 27.03793, 27.07128, 27.10448, 27.13754, 27.17044, 
    27.2032, 27.2358, 27.26825, 27.30055, 27.3327, 27.36469, 27.39653, 
    27.42822, 27.45976, 27.49115, 27.52238, 27.55346, 27.58438, 27.61515, 
    27.64577, 27.67623, 27.70654, 27.73669, 27.76669, 27.79653, 27.82622, 
    27.85575, 27.88512, 27.91434, 27.9434, 27.97231, 28.00105, 28.02965, 
    28.05808, 28.08636, 28.11447, 28.14243, 28.17023, 28.19788, 28.22536, 
    28.25269, 28.27986, 28.30686, 28.33371, 28.3604, 28.38693, 28.4133, 
    28.4395, 28.46555, 28.49144, 28.51716, 28.54272, 28.56813, 28.59337, 
    28.61845, 28.64336, 28.66812, 28.69271, 28.71714, 28.74141, 28.76551, 
    28.78945, 28.81322, 28.83684, 28.86029, 28.88357, 28.90669, 28.92965, 
    28.95244, 28.97507, 28.99753, 29.01983, 29.04196, 29.06392, 29.08572, 
    29.10736, 29.12883, 29.15013, 29.17126, 29.19223, 29.21303, 29.23367, 
    29.25414, 29.27444, 29.29457, 29.31454, 29.33433, 29.35396, 29.37342, 
    29.39272, 29.41184, 29.4308, 29.44958, 29.4682, 29.48665, 29.50493, 
    29.52304, 29.54098, 29.55875, 29.57635, 29.59378, 29.61104, 29.62813, 
    29.64505, 29.66179, 29.67837, 29.69478, 29.71102, 29.72708, 29.74297, 
    29.75869, 29.77424, 29.78962, 29.80483, 29.81986, 29.83472, 29.84941, 
    29.86393, 29.87827, 29.89244, 29.90644, 29.92027, 29.93392, 29.9474, 
    29.9607, 29.97383, 29.98679, 29.99958, 30.01219, 30.02463, 30.03689, 
    30.04898, 30.06089, 30.07264, 30.0842, 30.09559, 30.10681, 30.11785, 
    30.12872, 30.13941, 30.14993, 30.16027, 30.17044, 30.18043, 30.19024, 
    30.19988, 30.20935, 30.21864, 30.22775, 30.23669, 30.24545, 30.25404, 
    30.26245, 30.27068, 30.27874, 30.28662, 30.29432, 30.30185, 30.3092, 
    30.31638, 30.32338, 30.3302, 30.33684, 30.34331, 30.3496, 30.35571, 
    30.36165, 30.36741, 30.37299, 30.3784, 30.38363, 30.38868, 30.39355, 
    30.39825, 30.40277, 30.40711, 30.41128, 30.41526, 30.41907, 30.4227, 
    30.42616, 30.42943, 30.43253, 30.43545, 30.43819, 30.44076, 30.44315, 
    30.44536, 30.44739, 30.44924, 30.45092, 30.45242, 30.45374, 30.45488, 
    30.45584, 30.45663, 30.45724, 30.45767, 30.45792, 30.458, 30.4579, 
    30.45761, 30.45716, 30.45652, 30.45571, 30.45471, 30.45354, 30.45219, 
    30.45067, 30.44896, 30.44708, 30.44502, 30.44278, 30.44037, 30.43777, 
    30.435, 30.43205, 30.42893, 30.42562, 30.42214, 30.41848, 30.41464, 
    30.41063, 30.40644, 30.40207, 30.39752, 30.39279, 30.38789, 30.38281, 
    30.37756, 30.37212, 30.36651, 30.36072, 30.35476, 30.34862, 30.3423, 
    30.3358, 30.32913, 30.32228, 30.31525, 30.30805, 30.30067, 30.29312, 
    30.28538, 30.27748, 30.26939, 30.26113, 30.25269, 30.24408, 30.23529, 
    30.22632, 30.21718, 30.20786, 30.19837, 30.1887, 30.17886, 30.16884, 
    30.15865, 30.14828, 30.13773, 30.12701, 30.11612, 30.10505, 30.0938, 
    30.08238, 30.07079, 30.05902, 30.04708, 30.03496, 30.02267, 30.01021, 
    29.99757, 29.98476, 29.97177, 29.95861, 29.94528, 29.93177, 29.91809, 
    29.90424, 29.89021, 29.87601, 29.86164, 29.8471, 29.83238, 29.81749, 
    29.80243, 29.7872, 29.7718, 29.75622, 29.74047, 29.72455, 29.70846, 
    29.6922, 29.67576, 29.65916, 29.64238, 29.62544, 29.60832, 29.59103, 
    29.57358, 29.55595, 29.53815, 29.52018, 29.50205, 29.48374, 29.46527, 
    29.44662, 29.42781, 29.40883, 29.38968, 29.37036, 29.35087, 29.33121, 
    29.31139, 29.2914, 29.27124, 29.25091, 29.23042, 29.20975, 29.18893, 
    29.16793, 29.14677, 29.12544, 29.10395, 29.08229, 29.06046, 29.03847, 
    29.01631, 28.99399, 28.9715, 28.94885, 28.92603, 28.90305, 28.8799, 
    28.85659, 28.83311, 28.80947, 28.78567, 28.76171, 28.73758, 28.71329, 
    28.68883, 28.66421, 28.63943, 28.61449, 28.58939, 28.56412, 28.53869, 
    28.5131, 28.48735, 28.46144, 28.43537, 28.40914, 28.38274, 28.35619, 
    28.32948, 28.3026, 28.27557, 28.24838, 28.22103, 28.19352, 28.16585, 
    28.13802, 28.11003, 28.08189, 28.05359, 28.02513, 27.99652, 27.96774, 
    27.93881, 27.90973,
  24.6602, 24.70282, 24.74532, 24.78768, 24.8299, 24.872, 24.91396, 24.95578, 
    24.99747, 25.03902, 25.08044, 25.12172, 25.16287, 25.20387, 25.24475, 
    25.28548, 25.32608, 25.36654, 25.40687, 25.44705, 25.4871, 25.52701, 
    25.56678, 25.60641, 25.64591, 25.68526, 25.72447, 25.76355, 25.80248, 
    25.84127, 25.87992, 25.91843, 25.9568, 25.99503, 26.03312, 26.07106, 
    26.10886, 26.14652, 26.18403, 26.22141, 26.25863, 26.29572, 26.33266, 
    26.36946, 26.40611, 26.44262, 26.47898, 26.5152, 26.55127, 26.5872, 
    26.62298, 26.65861, 26.6941, 26.72944, 26.76463, 26.79968, 26.83458, 
    26.86933, 26.90393, 26.93839, 26.97269, 27.00685, 27.04086, 27.07472, 
    27.10843, 27.14198, 27.1754, 27.20865, 27.24176, 27.27472, 27.30753, 
    27.34018, 27.37269, 27.40504, 27.43724, 27.46929, 27.50119, 27.53293, 
    27.56452, 27.59595, 27.62724, 27.65837, 27.68934, 27.72017, 27.75083, 
    27.78135, 27.8117, 27.84191, 27.87196, 27.90185, 27.93158, 27.96116, 
    27.99059, 28.01986, 28.04897, 28.07792, 28.10672, 28.13536, 28.16384, 
    28.19216, 28.22033, 28.24834, 28.27619, 28.30388, 28.33141, 28.35878, 
    28.38599, 28.41305, 28.43994, 28.46667, 28.49325, 28.51966, 28.54591, 
    28.57201, 28.59794, 28.6237, 28.64931, 28.67476, 28.70004, 28.72517, 
    28.75013, 28.77492, 28.79956, 28.82403, 28.84834, 28.87248, 28.89646, 
    28.92028, 28.94394, 28.96743, 28.99075, 29.01391, 29.03691, 29.05974, 
    29.08241, 29.10491, 29.12724, 29.14941, 29.17142, 29.19326, 29.21493, 
    29.23643, 29.25777, 29.27895, 29.29995, 29.32079, 29.34146, 29.36197, 
    29.3823, 29.40247, 29.42247, 29.4423, 29.46197, 29.48146, 29.50079, 
    29.51995, 29.53894, 29.55776, 29.57641, 29.59489, 29.6132, 29.63134, 
    29.64932, 29.66712, 29.68475, 29.70221, 29.7195, 29.73662, 29.75357, 
    29.77035, 29.78696, 29.80339, 29.81966, 29.83575, 29.85167, 29.86742, 
    29.883, 29.8984, 29.91364, 29.9287, 29.94359, 29.9583, 29.97285, 
    29.98722, 30.00141, 30.01543, 30.02929, 30.04296, 30.05647, 30.0698, 
    30.08295, 30.09593, 30.10874, 30.12138, 30.13384, 30.14612, 30.15823, 
    30.17017, 30.18193, 30.19352, 30.20493, 30.21617, 30.22723, 30.23812, 
    30.24883, 30.25937, 30.26973, 30.27991, 30.28992, 30.29975, 30.30941, 
    30.31889, 30.3282, 30.33733, 30.34628, 30.35506, 30.36366, 30.37209, 
    30.38034, 30.38841, 30.3963, 30.40402, 30.41156, 30.41893, 30.42612, 
    30.43313, 30.43996, 30.44662, 30.4531, 30.4594, 30.46553, 30.47147, 
    30.47725, 30.48284, 30.48825, 30.49349, 30.49855, 30.50344, 30.50814, 
    30.51267, 30.51702, 30.52119, 30.52518, 30.529, 30.53264, 30.5361, 
    30.53938, 30.54248, 30.54541, 30.54816, 30.55073, 30.55312, 30.55533, 
    30.55737, 30.55923, 30.56091, 30.56241, 30.56373, 30.56487, 30.56584, 
    30.56663, 30.56724, 30.56767, 30.56792, 30.568, 30.5679, 30.56762, 
    30.56716, 30.56652, 30.5657, 30.56471, 30.56353, 30.56218, 30.56065, 
    30.55894, 30.55706, 30.555, 30.55275, 30.55033, 30.54774, 30.54496, 
    30.54201, 30.53887, 30.53556, 30.53207, 30.52841, 30.52456, 30.52054, 
    30.51634, 30.51196, 30.50741, 30.50267, 30.49776, 30.49268, 30.48741, 
    30.48197, 30.47634, 30.47054, 30.46457, 30.45842, 30.45209, 30.44558, 
    30.43889, 30.43203, 30.42499, 30.41778, 30.41038, 30.40281, 30.39507, 
    30.38714, 30.37904, 30.37077, 30.36231, 30.35369, 30.34488, 30.3359, 
    30.32674, 30.31741, 30.3079, 30.29821, 30.28835, 30.27831, 30.2681, 
    30.25771, 30.24714, 30.23641, 30.22549, 30.2144, 30.20314, 30.1917, 
    30.18008, 30.16829, 30.15633, 30.14419, 30.13188, 30.11939, 30.10673, 
    30.09389, 30.08088, 30.0677, 30.05434, 30.04081, 30.02711, 30.01323, 
    29.99918, 29.98495, 29.97056, 29.95599, 29.94124, 29.92633, 29.91124, 
    29.89598, 29.88055, 29.86494, 29.84916, 29.83322, 29.8171, 29.8008, 
    29.78434, 29.76771, 29.7509, 29.73392, 29.71678, 29.69946, 29.68197, 
    29.66431, 29.64648, 29.62848, 29.61032, 29.59198, 29.57347, 29.55479, 
    29.53595, 29.51693, 29.49774, 29.47839, 29.45887, 29.43918, 29.41932, 
    29.39929, 29.3791, 29.35873, 29.3382, 29.31751, 29.29664, 29.27561, 
    29.25441, 29.23304, 29.21151, 29.18981, 29.16795, 29.14592, 29.12372, 
    29.10136, 29.07883, 29.05614, 29.03328, 29.01026, 28.98707, 28.96372, 
    28.9402, 28.91652, 28.89268, 28.86867, 28.8445, 28.82017, 28.79567, 
    28.77101, 28.74619, 28.7212, 28.69605, 28.67075, 28.64527, 28.61964, 
    28.59385, 28.56789, 28.54177, 28.51549, 28.48906, 28.46246, 28.4357, 
    28.40878, 28.3817, 28.35446, 28.32706, 28.29951, 28.27179, 28.24392, 
    28.21588, 28.18769, 28.15934, 28.13084, 28.10217, 28.07335, 28.04437, 
    28.01524,
  24.76034, 24.80304, 24.84559, 24.88802, 24.93031, 24.97247, 25.01449, 
    25.05637, 25.09813, 25.13974, 25.18122, 25.22257, 25.26378, 25.30485, 
    25.34579, 25.38658, 25.42725, 25.46777, 25.50816, 25.5484, 25.58851, 
    25.62848, 25.66832, 25.70801, 25.74756, 25.78698, 25.82625, 25.86539, 
    25.90438, 25.94324, 25.98195, 26.02052, 26.05895, 26.09723, 26.13538, 
    26.17338, 26.21124, 26.24896, 26.28654, 26.32397, 26.36126, 26.3984, 
    26.4354, 26.47226, 26.50897, 26.54553, 26.58195, 26.61823, 26.65436, 
    26.69034, 26.72618, 26.76187, 26.79742, 26.83282, 26.86807, 26.90317, 
    26.93813, 26.97293, 27.00759, 27.0421, 27.07646, 27.11068, 27.14474, 
    27.17866, 27.21242, 27.24603, 27.2795, 27.31281, 27.34598, 27.37899, 
    27.41185, 27.44456, 27.47712, 27.50952, 27.54178, 27.57388, 27.60583, 
    27.63762, 27.66926, 27.70075, 27.73209, 27.76327, 27.7943, 27.82517, 
    27.85589, 27.88645, 27.91686, 27.94712, 27.97721, 28.00716, 28.03694, 
    28.06657, 28.09605, 28.12536, 28.15452, 28.18353, 28.21237, 28.24106, 
    28.26959, 28.29796, 28.32618, 28.35423, 28.38213, 28.40987, 28.43744, 
    28.46486, 28.49212, 28.51922, 28.54616, 28.57294, 28.59956, 28.62602, 
    28.65232, 28.67845, 28.70443, 28.73024, 28.75589, 28.78139, 28.80671, 
    28.83188, 28.85688, 28.88172, 28.9064, 28.93091, 28.95526, 28.97945, 
    29.00347, 29.02733, 29.05103, 29.07456, 29.09793, 29.12113, 29.14416, 
    29.16703, 29.18974, 29.21228, 29.23466, 29.25686, 29.27891, 29.30079, 
    29.32249, 29.34404, 29.36542, 29.38663, 29.40767, 29.42854, 29.44925, 
    29.46979, 29.49016, 29.51037, 29.5304, 29.55027, 29.56997, 29.5895, 
    29.60886, 29.62805, 29.64708, 29.66593, 29.68461, 29.70313, 29.72147, 
    29.73965, 29.75765, 29.77548, 29.79315, 29.81064, 29.82796, 29.84511, 
    29.86209, 29.8789, 29.89554, 29.912, 29.9283, 29.94442, 29.96037, 
    29.97615, 29.99175, 30.00718, 30.02245, 30.03753, 30.05245, 30.06719, 
    30.08176, 30.09616, 30.11038, 30.12443, 30.1383, 30.152, 30.16553, 
    30.17889, 30.19207, 30.20507, 30.2179, 30.23056, 30.24304, 30.25535, 
    30.26748, 30.27944, 30.29122, 30.30283, 30.31427, 30.32552, 30.33661, 
    30.34751, 30.35824, 30.3688, 30.37918, 30.38938, 30.39941, 30.40926, 
    30.41894, 30.42844, 30.43776, 30.44691, 30.45588, 30.46467, 30.47329, 
    30.48173, 30.48999, 30.49808, 30.50599, 30.51372, 30.52128, 30.52866, 
    30.53586, 30.54288, 30.54973, 30.5564, 30.56289, 30.5692, 30.57534, 
    30.5813, 30.58708, 30.59268, 30.59811, 30.60336, 30.60843, 30.61332, 
    30.61803, 30.62257, 30.62692, 30.6311, 30.63511, 30.63893, 30.64257, 
    30.64604, 30.64933, 30.65244, 30.65537, 30.65812, 30.6607, 30.66309, 
    30.66531, 30.66735, 30.66921, 30.67089, 30.6724, 30.67372, 30.67487, 
    30.67584, 30.67663, 30.67724, 30.67767, 30.67793, 30.678, 30.6779, 
    30.67761, 30.67715, 30.67651, 30.6757, 30.6747, 30.67352, 30.67217, 
    30.67064, 30.66893, 30.66704, 30.66497, 30.66273, 30.6603, 30.6577, 
    30.65492, 30.65196, 30.64882, 30.6455, 30.64201, 30.63833, 30.63448, 
    30.63045, 30.62625, 30.62186, 30.6173, 30.61255, 30.60763, 30.60254, 
    30.59726, 30.59181, 30.58618, 30.58037, 30.57438, 30.56821, 30.56187, 
    30.55535, 30.54866, 30.54178, 30.53473, 30.5275, 30.52009, 30.51251, 
    30.50475, 30.49681, 30.4887, 30.48041, 30.47194, 30.46329, 30.45447, 
    30.44547, 30.4363, 30.42695, 30.41742, 30.40771, 30.39784, 30.38778, 
    30.37755, 30.36714, 30.35656, 30.3458, 30.33486, 30.32375, 30.31247, 
    30.30101, 30.28937, 30.27756, 30.26558, 30.25341, 30.24108, 30.22857, 
    30.21589, 30.20303, 30.18999, 30.17678, 30.1634, 30.14985, 30.13612, 
    30.12222, 30.10814, 30.09389, 30.07947, 30.06487, 30.0501, 30.03516, 
    30.02004, 30.00476, 29.9893, 29.97366, 29.95786, 29.94188, 29.92573, 
    29.90941, 29.89292, 29.87625, 29.85942, 29.84241, 29.82523, 29.80788, 
    29.79037, 29.77267, 29.75481, 29.73678, 29.71858, 29.70021, 29.68167, 
    29.66296, 29.64408, 29.62503, 29.60581, 29.58642, 29.56686, 29.54714, 
    29.52724, 29.50718, 29.48695, 29.46655, 29.44599, 29.42525, 29.40435, 
    29.38328, 29.36205, 29.34064, 29.31907, 29.29733, 29.27543, 29.25336, 
    29.23113, 29.20873, 29.18616, 29.16343, 29.14053, 29.11747, 29.09424, 
    29.07085, 29.04729, 29.02357, 28.99968, 28.97564, 28.95142, 28.92705, 
    28.90251, 28.8778, 28.85294, 28.82791, 28.80272, 28.77736, 28.75185, 
    28.72617, 28.70033, 28.67433, 28.64817, 28.62185, 28.59536, 28.56872, 
    28.54191, 28.51495, 28.48782, 28.46054, 28.43309, 28.40549, 28.37773, 
    28.3498, 28.32172, 28.29349, 28.26509, 28.23653, 28.20782, 28.17895, 
    28.14992, 28.12074,
  24.86047, 24.90323, 24.94585, 24.98834, 25.03069, 25.07292, 25.115, 
    25.15695, 25.19877, 25.24045, 25.28199, 25.3234, 25.36467, 25.40581, 
    25.44681, 25.48767, 25.52839, 25.56898, 25.60943, 25.64974, 25.68991, 
    25.72994, 25.76984, 25.80959, 25.84921, 25.88868, 25.92802, 25.96721, 
    26.00627, 26.04518, 26.08396, 26.12259, 26.16108, 26.19943, 26.23763, 
    26.2757, 26.31362, 26.35139, 26.38903, 26.42652, 26.46387, 26.50107, 
    26.53813, 26.57504, 26.61181, 26.64844, 26.68492, 26.72125, 26.75744, 
    26.79348, 26.82937, 26.86512, 26.90073, 26.93618, 26.97149, 27.00665, 
    27.04166, 27.07652, 27.11124, 27.14581, 27.18022, 27.21449, 27.24861, 
    27.28258, 27.3164, 27.35007, 27.38359, 27.41696, 27.45018, 27.48324, 
    27.51616, 27.54892, 27.58153, 27.61399, 27.6463, 27.67845, 27.71046, 
    27.7423, 27.774, 27.80554, 27.83693, 27.86816, 27.89924, 27.93017, 
    27.96094, 27.99155, 28.02201, 28.05231, 28.08246, 28.11246, 28.14229, 
    28.17197, 28.2015, 28.23086, 28.26007, 28.28912, 28.31802, 28.34675, 
    28.37533, 28.40375, 28.43201, 28.46012, 28.48806, 28.51585, 28.54347, 
    28.57094, 28.59825, 28.62539, 28.65238, 28.6792, 28.70587, 28.73237, 
    28.75871, 28.78489, 28.81091, 28.83677, 28.86247, 28.888, 28.91337, 
    28.93858, 28.96363, 28.98851, 29.01323, 29.03779, 29.06218, 29.08641, 
    29.11048, 29.13438, 29.15811, 29.18168, 29.20509, 29.22833, 29.25141, 
    29.27432, 29.29707, 29.31965, 29.34206, 29.36431, 29.38639, 29.40831, 
    29.43006, 29.45164, 29.47305, 29.4943, 29.51538, 29.53629, 29.55704, 
    29.57761, 29.59802, 29.61826, 29.63833, 29.65823, 29.67797, 29.69753, 
    29.71693, 29.73615, 29.75521, 29.7741, 29.79281, 29.81136, 29.82974, 
    29.84795, 29.86598, 29.88385, 29.90154, 29.91907, 29.93642, 29.9536, 
    29.97061, 29.98745, 30.00412, 30.02061, 30.03693, 30.05309, 30.06906, 
    30.08487, 30.1005, 30.11596, 30.13125, 30.14637, 30.16131, 30.17608, 
    30.19067, 30.20509, 30.21934, 30.23342, 30.24732, 30.26104, 30.2746, 
    30.28797, 30.30118, 30.31421, 30.32706, 30.33974, 30.35225, 30.36458, 
    30.37673, 30.38871, 30.40052, 30.41215, 30.4236, 30.43488, 30.44598, 
    30.45691, 30.46766, 30.47823, 30.48863, 30.49885, 30.5089, 30.51877, 
    30.52846, 30.53798, 30.54732, 30.55648, 30.56547, 30.57428, 30.58291, 
    30.59137, 30.59965, 30.60775, 30.61567, 30.62342, 30.63099, 30.63838, 
    30.6456, 30.65263, 30.65949, 30.66617, 30.67268, 30.679, 30.68515, 
    30.69112, 30.69691, 30.70252, 30.70796, 30.71322, 30.7183, 30.7232, 
    30.72792, 30.73246, 30.73683, 30.74102, 30.74503, 30.74886, 30.75251, 
    30.75598, 30.75927, 30.76239, 30.76533, 30.76809, 30.77066, 30.77307, 
    30.77529, 30.77733, 30.7792, 30.78088, 30.78239, 30.78371, 30.78486, 
    30.78583, 30.78662, 30.78724, 30.78767, 30.78792, 30.788, 30.7879, 
    30.78761, 30.78715, 30.78651, 30.78569, 30.78469, 30.78352, 30.78216, 
    30.78063, 30.77891, 30.77702, 30.77495, 30.7727, 30.77027, 30.76766, 
    30.76487, 30.76191, 30.75876, 30.75544, 30.75194, 30.74826, 30.7444, 
    30.74037, 30.73615, 30.73176, 30.72718, 30.72243, 30.7175, 30.7124, 
    30.70711, 30.70165, 30.69601, 30.69019, 30.68419, 30.67801, 30.67166, 
    30.66513, 30.65842, 30.65153, 30.64447, 30.63722, 30.6298, 30.62221, 
    30.61443, 30.60648, 30.59835, 30.59004, 30.58156, 30.5729, 30.56406, 
    30.55505, 30.54585, 30.53649, 30.52694, 30.51722, 30.50732, 30.49725, 
    30.487, 30.47657, 30.46597, 30.45519, 30.44423, 30.43311, 30.4218, 
    30.41032, 30.39866, 30.38683, 30.37482, 30.36264, 30.35028, 30.33775, 
    30.32504, 30.31216, 30.2991, 30.28587, 30.27246, 30.25888, 30.24513, 
    30.2312, 30.2171, 30.20282, 30.18838, 30.17375, 30.15896, 30.14399, 
    30.12885, 30.11353, 30.09804, 30.08238, 30.06655, 30.05054, 30.03436, 
    30.01801, 30.00149, 29.9848, 29.96793, 29.95089, 29.93369, 29.91631, 
    29.89875, 29.88103, 29.86314, 29.84508, 29.82684, 29.80844, 29.78987, 
    29.77112, 29.75221, 29.73312, 29.71387, 29.69445, 29.67486, 29.6551, 
    29.63517, 29.61507, 29.5948, 29.57437, 29.55376, 29.53299, 29.51205, 
    29.49095, 29.46968, 29.44823, 29.42663, 29.40485, 29.38291, 29.3608, 
    29.33853, 29.31609, 29.29348, 29.27071, 29.24777, 29.22467, 29.2014, 
    29.17797, 29.15437, 29.13061, 29.10668, 29.08259, 29.05833, 29.03392, 
    29.00933, 28.98459, 28.95968, 28.93461, 28.90937, 28.88397, 28.85842, 
    28.83269, 28.80681, 28.78076, 28.75456, 28.72819, 28.70166, 28.67497, 
    28.64812, 28.62111, 28.59394, 28.5666, 28.53911, 28.51146, 28.48365, 
    28.45568, 28.42756, 28.39927, 28.37082, 28.34222, 28.31346, 28.28454, 
    28.25546, 28.22623,
  24.96059, 25.00341, 25.04609, 25.08865, 25.13107, 25.17335, 25.2155, 
    25.25751, 25.29939, 25.34114, 25.38274, 25.42422, 25.46555, 25.50675, 
    25.54781, 25.58874, 25.62952, 25.67017, 25.71068, 25.75106, 25.79129, 
    25.83139, 25.87134, 25.91116, 25.95084, 25.99037, 26.02977, 26.06903, 
    26.10814, 26.14712, 26.18595, 26.22464, 26.2632, 26.3016, 26.33987, 
    26.37799, 26.41597, 26.45381, 26.4915, 26.52905, 26.56646, 26.60372, 
    26.64084, 26.67782, 26.71464, 26.75133, 26.78786, 26.82426, 26.8605, 
    26.8966, 26.93256, 26.96836, 27.00402, 27.03953, 27.0749, 27.11012, 
    27.14518, 27.1801, 27.21488, 27.2495, 27.28397, 27.3183, 27.35247, 
    27.3865, 27.42037, 27.4541, 27.48767, 27.52109, 27.55437, 27.58749, 
    27.62046, 27.65327, 27.68594, 27.71845, 27.75081, 27.78302, 27.81507, 
    27.84698, 27.87873, 27.91032, 27.94176, 27.97304, 28.00418, 28.03515, 
    28.06597, 28.09664, 28.12715, 28.15751, 28.1877, 28.21775, 28.24763, 
    28.27736, 28.30694, 28.33635, 28.36561, 28.39471, 28.42365, 28.45244, 
    28.48107, 28.50953, 28.53785, 28.566, 28.59399, 28.62182, 28.64949, 
    28.67701, 28.70436, 28.73155, 28.75858, 28.78545, 28.81216, 28.83871, 
    28.8651, 28.89133, 28.91739, 28.9433, 28.96904, 28.99461, 29.02003, 
    29.04528, 29.07037, 29.0953, 29.12006, 29.14466, 29.16909, 29.19337, 
    29.21747, 29.24142, 29.26519, 29.28881, 29.31225, 29.33554, 29.35865, 
    29.38161, 29.40439, 29.42701, 29.44946, 29.47175, 29.49387, 29.51583, 
    29.53761, 29.55923, 29.58068, 29.60197, 29.62308, 29.64403, 29.66481, 
    29.68543, 29.70587, 29.72615, 29.74625, 29.76619, 29.78596, 29.80556, 
    29.82499, 29.84425, 29.86334, 29.88226, 29.90101, 29.91959, 29.938, 
    29.95624, 29.97431, 29.99221, 30.00993, 30.02749, 30.04487, 30.06208, 
    30.07912, 30.09599, 30.11269, 30.12922, 30.14557, 30.16175, 30.17775, 
    30.19359, 30.20925, 30.22474, 30.24006, 30.2552, 30.27017, 30.28496, 
    30.29958, 30.31403, 30.3283, 30.3424, 30.35633, 30.37008, 30.38366, 
    30.39706, 30.41029, 30.42334, 30.43622, 30.44892, 30.46145, 30.4738, 
    30.48598, 30.49798, 30.50981, 30.52146, 30.53293, 30.54423, 30.55535, 
    30.5663, 30.57707, 30.58766, 30.59808, 30.60832, 30.61839, 30.62827, 
    30.63799, 30.64752, 30.65688, 30.66606, 30.67506, 30.68389, 30.69254, 
    30.70101, 30.7093, 30.71742, 30.72536, 30.73312, 30.7407, 30.74811, 
    30.75533, 30.76238, 30.76925, 30.77595, 30.78246, 30.7888, 30.79496, 
    30.80094, 30.80674, 30.81237, 30.81781, 30.82308, 30.82817, 30.83308, 
    30.83781, 30.84236, 30.84674, 30.85093, 30.85495, 30.85878, 30.86244, 
    30.86592, 30.86922, 30.87234, 30.87529, 30.87805, 30.88063, 30.88304, 
    30.88526, 30.88731, 30.88918, 30.89087, 30.89238, 30.89371, 30.89486, 
    30.89583, 30.89662, 30.89724, 30.89767, 30.89792, 30.898, 30.8979, 
    30.89761, 30.89715, 30.89651, 30.89569, 30.89469, 30.89351, 30.89215, 
    30.89061, 30.8889, 30.887, 30.88492, 30.88267, 30.88024, 30.87762, 
    30.87483, 30.87186, 30.86871, 30.86538, 30.86188, 30.85819, 30.85432, 
    30.85028, 30.84606, 30.84165, 30.83707, 30.83231, 30.82738, 30.82226, 
    30.81696, 30.81149, 30.80584, 30.80001, 30.794, 30.78781, 30.78144, 
    30.7749, 30.76818, 30.76128, 30.7542, 30.74695, 30.73951, 30.7319, 
    30.72411, 30.71614, 30.708, 30.69968, 30.69118, 30.6825, 30.67365, 
    30.66462, 30.65541, 30.64602, 30.63646, 30.62672, 30.61681, 30.60671, 
    30.59645, 30.586, 30.57538, 30.56458, 30.55361, 30.54246, 30.53113, 
    30.51963, 30.50795, 30.49609, 30.48406, 30.47186, 30.45948, 30.44692, 
    30.43419, 30.42129, 30.40821, 30.39495, 30.38152, 30.36792, 30.35414, 
    30.34019, 30.32606, 30.31176, 30.29728, 30.28263, 30.26781, 30.25281, 
    30.23764, 30.2223, 30.20679, 30.1911, 30.17523, 30.1592, 30.14299, 
    30.12661, 30.11006, 30.09334, 30.07644, 30.05937, 30.04213, 30.02472, 
    30.00714, 29.98939, 29.97146, 29.95337, 29.9351, 29.91666, 29.89806, 
    29.87928, 29.86033, 29.84122, 29.82193, 29.80247, 29.78284, 29.76305, 
    29.74308, 29.72295, 29.70265, 29.68218, 29.66154, 29.64073, 29.61975, 
    29.59861, 29.5773, 29.55582, 29.53418, 29.51236, 29.49038, 29.46824, 
    29.44592, 29.42344, 29.4008, 29.37799, 29.35501, 29.33187, 29.30856, 
    29.28508, 29.26144, 29.23764, 29.21367, 29.18954, 29.16524, 29.14078, 
    29.11615, 29.09137, 29.06641, 29.0413, 29.01602, 28.99058, 28.96498, 
    28.93921, 28.91328, 28.88719, 28.86094, 28.83453, 28.80795, 28.78121, 
    28.75432, 28.72726, 28.70004, 28.67266, 28.64513, 28.61743, 28.58957, 
    28.56155, 28.53338, 28.50504, 28.47655, 28.4479, 28.41909, 28.39012, 
    28.36099, 28.33171,
  25.06068, 25.10357, 25.14632, 25.18894, 25.23142, 25.27377, 25.31598, 
    25.35806, 25.4, 25.44181, 25.48348, 25.52502, 25.56642, 25.60768, 
    25.6488, 25.68979, 25.73064, 25.77135, 25.81192, 25.85236, 25.89266, 
    25.93281, 25.97283, 26.01271, 26.05245, 26.09205, 26.13151, 26.17082, 
    26.21, 26.24904, 26.28793, 26.32668, 26.3653, 26.40376, 26.44209, 
    26.48028, 26.51832, 26.55621, 26.59397, 26.63158, 26.66904, 26.70637, 
    26.74354, 26.78057, 26.81746, 26.8542, 26.8908, 26.92725, 26.96355, 
    26.99971, 27.03572, 27.07159, 27.1073, 27.14287, 27.1783, 27.21357, 
    27.24869, 27.28367, 27.3185, 27.35318, 27.38771, 27.42209, 27.45632, 
    27.4904, 27.52433, 27.55811, 27.59174, 27.62522, 27.65854, 27.69172, 
    27.72474, 27.75762, 27.79033, 27.8229, 27.85532, 27.88758, 27.91968, 
    27.95164, 27.98344, 28.01509, 28.04658, 28.07792, 28.1091, 28.14013, 
    28.171, 28.20172, 28.23228, 28.26268, 28.29293, 28.32303, 28.35296, 
    28.38274, 28.41237, 28.44183, 28.47114, 28.50029, 28.52928, 28.55812, 
    28.58679, 28.61531, 28.64367, 28.67187, 28.69991, 28.72779, 28.7555, 
    28.78306, 28.81046, 28.8377, 28.86478, 28.8917, 28.91846, 28.94505, 
    28.97148, 28.99776, 29.02386, 29.04981, 29.0756, 29.10122, 29.12668, 
    29.15197, 29.17711, 29.20208, 29.22688, 29.25152, 29.276, 29.30031, 
    29.32446, 29.34845, 29.37227, 29.39592, 29.41941, 29.44273, 29.46589, 
    29.48888, 29.51171, 29.53437, 29.55686, 29.57919, 29.60134, 29.62334, 
    29.64516, 29.66682, 29.68831, 29.70963, 29.73079, 29.75177, 29.77259, 
    29.79324, 29.81372, 29.83403, 29.85417, 29.87415, 29.89395, 29.91358, 
    29.93305, 29.95234, 29.97147, 29.99042, 30.0092, 30.02782, 30.04626, 
    30.06453, 30.08263, 30.10056, 30.11832, 30.13591, 30.15332, 30.17056, 
    30.18764, 30.20453, 30.22126, 30.23782, 30.2542, 30.27041, 30.28644, 
    30.30231, 30.318, 30.33351, 30.34886, 30.36403, 30.37902, 30.39384, 
    30.40849, 30.42296, 30.43726, 30.45139, 30.46534, 30.47912, 30.49272, 
    30.50615, 30.5194, 30.53247, 30.54537, 30.5581, 30.57065, 30.58302, 
    30.59522, 30.60725, 30.6191, 30.63077, 30.64226, 30.65358, 30.66472, 
    30.67569, 30.68648, 30.6971, 30.70753, 30.71779, 30.72787, 30.73778, 
    30.74751, 30.75706, 30.76644, 30.77563, 30.78465, 30.79349, 30.80216, 
    30.81064, 30.81895, 30.82709, 30.83504, 30.84281, 30.85041, 30.85783, 
    30.86507, 30.87213, 30.87902, 30.88572, 30.89225, 30.8986, 30.90477, 
    30.91076, 30.91657, 30.92221, 30.92767, 30.93294, 30.93804, 30.94296, 
    30.9477, 30.95226, 30.95664, 30.96084, 30.96487, 30.96871, 30.97238, 
    30.97586, 30.97917, 30.9823, 30.98524, 30.98801, 30.9906, 30.99301, 
    30.99524, 30.99729, 30.99916, 31.00085, 31.00237, 31.0037, 31.00485, 
    31.00583, 31.00662, 31.00723, 31.00767, 31.00792, 31.008, 31.0079, 
    31.00761, 31.00715, 31.00651, 31.00568, 31.00468, 31.0035, 31.00214, 
    31.0006, 30.99888, 30.99698, 30.9949, 30.99264, 30.9902, 30.98759, 
    30.98479, 30.98181, 30.97866, 30.97532, 30.97181, 30.96811, 30.96424, 
    30.96019, 30.95596, 30.95155, 30.94696, 30.94219, 30.93724, 30.93212, 
    30.92681, 30.92133, 30.91567, 30.90983, 30.90381, 30.89761, 30.89123, 
    30.88467, 30.87794, 30.87103, 30.86394, 30.85667, 30.84922, 30.8416, 
    30.83379, 30.82581, 30.81765, 30.80931, 30.8008, 30.79211, 30.78324, 
    30.77419, 30.76497, 30.75556, 30.74598, 30.73623, 30.72629, 30.71618, 
    30.70589, 30.69543, 30.68479, 30.67397, 30.66298, 30.6518, 30.64046, 
    30.62893, 30.61723, 30.60536, 30.59331, 30.58108, 30.56868, 30.5561, 
    30.54334, 30.53042, 30.51731, 30.50403, 30.49058, 30.47695, 30.46315, 
    30.44917, 30.43501, 30.42069, 30.40619, 30.39151, 30.37666, 30.36164, 
    30.34644, 30.33107, 30.31553, 30.29981, 30.28392, 30.26785, 30.25162, 
    30.23521, 30.21863, 30.20187, 30.18495, 30.16785, 30.15058, 30.13314, 
    30.11552, 30.09774, 30.07978, 30.06165, 30.04336, 30.02489, 30.00624, 
    29.98743, 29.96845, 29.9493, 29.92998, 29.91049, 29.89083, 29.871, 
    29.851, 29.83083, 29.81049, 29.78998, 29.76931, 29.74846, 29.72745, 
    29.70627, 29.68492, 29.6634, 29.64172, 29.61987, 29.59785, 29.57566, 
    29.55331, 29.53079, 29.50811, 29.48526, 29.46224, 29.43905, 29.4157, 
    29.39219, 29.36851, 29.34466, 29.32065, 29.29648, 29.27214, 29.24764, 
    29.22297, 29.19814, 29.17314, 29.14798, 29.12266, 29.09718, 29.07153, 
    29.04572, 29.01974, 28.99361, 28.96731, 28.94085, 28.91423, 28.88745, 
    28.86051, 28.8334, 28.80614, 28.77872, 28.75113, 28.72338, 28.69548, 
    28.66742, 28.63919, 28.61081, 28.58227, 28.55357, 28.52471, 28.49569, 
    28.46651, 28.43718,
  25.16076, 25.20371, 25.24653, 25.28921, 25.33176, 25.37417, 25.41645, 
    25.45859, 25.5006, 25.54247, 25.5842, 25.6258, 25.66726, 25.70859, 
    25.74977, 25.79082, 25.83174, 25.87251, 25.91315, 25.95365, 25.99401, 
    26.03423, 26.07431, 26.11425, 26.15405, 26.19371, 26.23323, 26.27261, 
    26.31185, 26.35094, 26.3899, 26.42871, 26.46738, 26.50591, 26.5443, 
    26.58254, 26.62065, 26.6586, 26.69642, 26.73409, 26.77161, 26.80899, 
    26.84623, 26.88332, 26.92027, 26.95707, 26.99372, 27.03023, 27.06659, 
    27.10281, 27.13888, 27.1748, 27.21057, 27.2462, 27.28168, 27.31701, 
    27.35219, 27.38723, 27.42211, 27.45685, 27.49143, 27.52587, 27.56016, 
    27.59429, 27.62828, 27.66211, 27.6958, 27.72933, 27.76271, 27.79594, 
    27.82902, 27.86195, 27.89472, 27.92734, 27.95981, 27.99212, 28.02428, 
    28.05629, 28.08814, 28.11984, 28.15139, 28.18278, 28.21401, 28.24509, 
    28.27602, 28.30679, 28.3374, 28.36786, 28.39816, 28.4283, 28.45829, 
    28.48812, 28.51779, 28.5473, 28.57666, 28.60586, 28.6349, 28.66379, 
    28.69251, 28.72108, 28.74948, 28.77773, 28.80581, 28.83374, 28.86151, 
    28.88911, 28.91656, 28.94385, 28.97097, 28.99793, 29.02474, 29.05138, 
    29.07786, 29.10417, 29.13033, 29.15632, 29.18215, 29.20782, 29.23332, 
    29.25866, 29.28383, 29.30885, 29.3337, 29.35838, 29.3829, 29.40726, 
    29.43145, 29.45547, 29.47933, 29.50303, 29.52656, 29.54992, 29.57312, 
    29.59615, 29.61902, 29.64172, 29.66425, 29.68661, 29.70881, 29.73084, 
    29.75271, 29.7744, 29.79593, 29.81729, 29.83848, 29.8595, 29.88036, 
    29.90104, 29.92156, 29.94191, 29.96209, 29.98209, 30.00193, 30.0216, 
    30.0411, 30.06043, 30.07959, 30.09858, 30.11739, 30.13604, 30.15452, 
    30.17282, 30.19095, 30.20892, 30.22671, 30.24432, 30.26177, 30.27904, 
    30.29614, 30.31307, 30.32983, 30.34641, 30.36283, 30.37906, 30.39513, 
    30.41102, 30.42674, 30.44228, 30.45765, 30.47285, 30.48787, 30.50272, 
    30.5174, 30.5319, 30.54622, 30.56037, 30.57435, 30.58815, 30.60178, 
    30.61523, 30.6285, 30.6416, 30.65453, 30.66728, 30.67985, 30.69225, 
    30.70447, 30.71651, 30.72838, 30.74008, 30.75159, 30.76293, 30.7741, 
    30.78508, 30.79589, 30.80652, 30.81698, 30.82726, 30.83736, 30.84728, 
    30.85703, 30.8666, 30.87599, 30.8852, 30.89424, 30.9031, 30.91178, 
    30.92028, 30.92861, 30.93675, 30.94472, 30.95251, 30.96012, 30.96755, 
    30.97481, 30.98188, 30.98878, 30.9955, 31.00204, 31.0084, 31.01458, 
    31.02058, 31.02641, 31.03205, 31.03752, 31.0428, 31.04791, 31.05284, 
    31.05759, 31.06216, 31.06655, 31.07076, 31.07479, 31.07864, 31.08231, 
    31.0858, 31.08912, 31.09225, 31.0952, 31.09797, 31.10057, 31.10298, 
    31.10522, 31.10727, 31.10915, 31.11084, 31.11236, 31.11369, 31.11485, 
    31.11582, 31.11662, 31.11723, 31.11767, 31.11792, 31.118, 31.1179, 
    31.11761, 31.11715, 31.1165, 31.11568, 31.11468, 31.11349, 31.11213, 
    31.11058, 31.10886, 31.10696, 31.10488, 31.10261, 31.10017, 31.09755, 
    31.09475, 31.09176, 31.0886, 31.08526, 31.08174, 31.07804, 31.07416, 
    31.0701, 31.06586, 31.06145, 31.05685, 31.05207, 31.04712, 31.04198, 
    31.03666, 31.03117, 31.0255, 31.01965, 31.01361, 31.0074, 31.00101, 
    30.99445, 30.9877, 30.98078, 30.97367, 30.96639, 30.95893, 30.95129, 
    30.94347, 30.93548, 30.9273, 30.91895, 30.91042, 30.90171, 30.89282, 
    30.88376, 30.87452, 30.8651, 30.8555, 30.84573, 30.83577, 30.82565, 
    30.81534, 30.80486, 30.79419, 30.78336, 30.77234, 30.76115, 30.74978, 
    30.73824, 30.72652, 30.71462, 30.70255, 30.6903, 30.67787, 30.66527, 
    30.65249, 30.63954, 30.62642, 30.61311, 30.59963, 30.58598, 30.57215, 
    30.55815, 30.54397, 30.52961, 30.51509, 30.50039, 30.48551, 30.47046, 
    30.45523, 30.43983, 30.42426, 30.40852, 30.3926, 30.37651, 30.36024, 
    30.3438, 30.32719, 30.31041, 30.29345, 30.27632, 30.25902, 30.24155, 
    30.2239, 30.20609, 30.1881, 30.16994, 30.15161, 30.1331, 30.11443, 
    30.09558, 30.07657, 30.05738, 30.03803, 30.0185, 29.99881, 29.97894, 
    29.9589, 29.9387, 29.91833, 29.89778, 29.87707, 29.85619, 29.83514, 
    29.81392, 29.79254, 29.77098, 29.74926, 29.72737, 29.70531, 29.68309, 
    29.6607, 29.63814, 29.61541, 29.59252, 29.56946, 29.54624, 29.52285, 
    29.49929, 29.47557, 29.45168, 29.42763, 29.40341, 29.37903, 29.35449, 
    29.32977, 29.3049, 29.27986, 29.25466, 29.22929, 29.20377, 29.17807, 
    29.15222, 29.1262, 29.10002, 29.07368, 29.04717, 29.02051, 28.99368, 
    28.96669, 28.93954, 28.91223, 28.88476, 28.85713, 28.82933, 28.80138, 
    28.77327, 28.745, 28.71657, 28.68798, 28.65923, 28.63032, 28.60125, 
    28.57203, 28.54265,
  25.26082, 25.30384, 25.34672, 25.38947, 25.43208, 25.47455, 25.5169, 
    25.5591, 25.60117, 25.64311, 25.68491, 25.72657, 25.76809, 25.80948, 
    25.85073, 25.89185, 25.93282, 25.97366, 26.01436, 26.05492, 26.09534, 
    26.13562, 26.17576, 26.21577, 26.25563, 26.29535, 26.33493, 26.37437, 
    26.41368, 26.45283, 26.49185, 26.53073, 26.56946, 26.60805, 26.64649, 
    26.6848, 26.72296, 26.76098, 26.79885, 26.83658, 26.87416, 26.91161, 
    26.9489, 26.98605, 27.02306, 27.05992, 27.09663, 27.1332, 27.16962, 
    27.20589, 27.24202, 27.278, 27.31383, 27.34951, 27.38505, 27.42044, 
    27.45568, 27.49077, 27.52571, 27.5605, 27.59514, 27.62964, 27.66398, 
    27.69817, 27.73221, 27.7661, 27.79984, 27.83343, 27.86687, 27.90015, 
    27.93328, 27.96626, 27.99909, 28.03177, 28.06429, 28.09665, 28.12887, 
    28.16093, 28.19284, 28.22459, 28.25619, 28.28763, 28.31891, 28.35005, 
    28.38102, 28.41184, 28.44251, 28.47301, 28.50337, 28.53356, 28.5636, 
    28.59348, 28.6232, 28.65277, 28.68217, 28.71142, 28.74051, 28.76944, 
    28.79822, 28.82683, 28.85529, 28.88358, 28.91171, 28.93969, 28.9675, 
    28.99516, 29.02265, 29.04998, 29.07715, 29.10416, 29.13101, 29.1577, 
    29.18422, 29.21058, 29.23678, 29.26282, 29.28869, 29.3144, 29.33995, 
    29.36534, 29.39055, 29.41561, 29.4405, 29.46523, 29.48979, 29.51419, 
    29.53842, 29.56249, 29.58639, 29.61013, 29.6337, 29.65711, 29.68034, 
    29.70342, 29.72632, 29.74906, 29.77163, 29.79404, 29.81627, 29.83834, 
    29.86024, 29.88198, 29.90355, 29.92494, 29.94617, 29.96723, 29.98812, 
    30.00884, 30.0294, 30.04978, 30.06999, 30.09004, 30.10991, 30.12962, 
    30.14915, 30.16851, 30.18771, 30.20673, 30.22558, 30.24426, 30.26277, 
    30.28111, 30.29927, 30.31726, 30.33508, 30.35274, 30.37021, 30.38752, 
    30.40465, 30.42161, 30.4384, 30.45501, 30.47145, 30.48772, 30.50381, 
    30.51973, 30.53548, 30.55105, 30.56645, 30.58167, 30.59672, 30.6116, 
    30.6263, 30.64083, 30.65518, 30.66935, 30.68336, 30.69718, 30.71083, 
    30.72431, 30.73761, 30.75073, 30.76368, 30.77645, 30.78905, 30.80147, 
    30.81371, 30.82578, 30.83767, 30.84938, 30.86092, 30.87228, 30.88346, 
    30.89447, 30.9053, 30.91595, 30.92643, 30.93673, 30.94684, 30.95679, 
    30.96655, 30.97614, 30.98555, 30.99478, 31.00383, 31.0127, 31.0214, 
    31.02992, 31.03826, 31.04642, 31.0544, 31.0622, 31.06983, 31.07728, 
    31.08455, 31.09163, 31.09854, 31.10527, 31.11182, 31.1182, 31.12439, 
    31.1304, 31.13624, 31.14189, 31.14737, 31.15266, 31.15778, 31.16272, 
    31.16747, 31.17205, 31.17645, 31.18067, 31.18471, 31.18857, 31.19225, 
    31.19574, 31.19906, 31.2022, 31.20516, 31.20794, 31.21054, 31.21296, 
    31.21519, 31.21725, 31.21913, 31.22083, 31.22235, 31.22368, 31.22484, 
    31.22582, 31.22661, 31.22723, 31.22767, 31.22792, 31.228, 31.2279, 
    31.22761, 31.22715, 31.2265, 31.22568, 31.22467, 31.22348, 31.22212, 
    31.22057, 31.21885, 31.21694, 31.21485, 31.21259, 31.21014, 31.20751, 
    31.2047, 31.20172, 31.19855, 31.1952, 31.19168, 31.18797, 31.18408, 
    31.18001, 31.17577, 31.17134, 31.16673, 31.16195, 31.15698, 31.15184, 
    31.14651, 31.14101, 31.13533, 31.12947, 31.12342, 31.1172, 31.1108, 
    31.10422, 31.09746, 31.09052, 31.08341, 31.07611, 31.06864, 31.06098, 
    31.05315, 31.04514, 31.03695, 31.02858, 31.02004, 31.01131, 31.00241, 
    30.99333, 30.98407, 30.97463, 30.96502, 30.95523, 30.94526, 30.93511, 
    30.92478, 30.91428, 30.9036, 30.89274, 30.88171, 30.8705, 30.85911, 
    30.84754, 30.8358, 30.82388, 30.81179, 30.79951, 30.78707, 30.77444, 
    30.76164, 30.74867, 30.73552, 30.72219, 30.70868, 30.69501, 30.68115, 
    30.66712, 30.65292, 30.63854, 30.62399, 30.60926, 30.59435, 30.57928, 
    30.56402, 30.5486, 30.533, 30.51722, 30.50128, 30.48516, 30.46886, 
    30.45239, 30.43575, 30.41894, 30.40195, 30.38479, 30.36746, 30.34995, 
    30.33228, 30.31443, 30.29641, 30.27822, 30.25985, 30.24132, 30.22261, 
    30.20373, 30.18468, 30.16546, 30.14607, 30.12651, 30.10678, 30.08688, 
    30.06681, 30.04657, 30.02616, 30.00558, 29.98483, 29.96391, 29.94282, 
    29.92157, 29.90014, 29.87855, 29.85679, 29.83486, 29.81277, 29.7905, 
    29.76807, 29.74548, 29.72271, 29.69978, 29.67668, 29.65342, 29.62998, 
    29.60639, 29.58262, 29.55869, 29.5346, 29.51034, 29.48592, 29.46133, 
    29.43658, 29.41166, 29.38658, 29.36133, 29.33592, 29.31035, 29.28461, 
    29.25871, 29.23265, 29.20642, 29.18004, 29.15349, 29.12678, 29.0999, 
    29.07287, 29.04567, 29.01831, 28.99079, 28.96311, 28.93527, 28.90727, 
    28.87911, 28.85079, 28.82232, 28.79368, 28.76488, 28.73592, 28.70681, 
    28.67753, 28.6481,
  25.36087, 25.40395, 25.44689, 25.4897, 25.53238, 25.57492, 25.61733, 
    25.6596, 25.70173, 25.74373, 25.78559, 25.82732, 25.86891, 25.91036, 
    25.95167, 25.99285, 26.03389, 26.07479, 26.11555, 26.15617, 26.19666, 
    26.237, 26.27721, 26.31727, 26.3572, 26.39698, 26.43662, 26.47613, 
    26.51549, 26.55471, 26.59379, 26.63272, 26.67152, 26.71017, 26.74867, 
    26.78704, 26.82526, 26.86334, 26.90127, 26.93906, 26.97671, 27.01421, 
    27.05156, 27.08877, 27.12583, 27.16275, 27.19952, 27.23615, 27.27263, 
    27.30896, 27.34515, 27.38118, 27.41707, 27.45282, 27.48841, 27.52386, 
    27.55915, 27.5943, 27.6293, 27.66414, 27.69884, 27.73339, 27.76779, 
    27.80204, 27.83614, 27.87008, 27.90388, 27.93752, 27.97101, 28.00435, 
    28.03754, 28.07057, 28.10345, 28.13618, 28.16876, 28.20118, 28.23345, 
    28.26556, 28.29752, 28.32932, 28.36097, 28.39247, 28.42381, 28.45499, 
    28.48602, 28.51689, 28.54761, 28.57817, 28.60857, 28.63881, 28.6689, 
    28.69883, 28.72861, 28.75822, 28.78768, 28.81697, 28.84611, 28.8751, 
    28.90392, 28.93258, 28.96108, 28.98942, 29.01761, 29.04563, 29.07349, 
    29.10119, 29.12873, 29.15611, 29.18333, 29.21038, 29.23728, 29.26401, 
    29.29058, 29.31699, 29.34323, 29.36931, 29.39523, 29.42099, 29.44658, 
    29.47201, 29.49727, 29.52237, 29.5473, 29.57207, 29.59668, 29.62112, 
    29.6454, 29.6695, 29.69345, 29.71723, 29.74084, 29.76428, 29.78756, 
    29.81067, 29.83362, 29.8564, 29.87901, 29.90145, 29.92373, 29.94584, 
    29.96778, 29.98955, 30.01115, 30.03259, 30.05386, 30.07495, 30.09588, 
    30.11664, 30.13723, 30.15765, 30.1779, 30.19798, 30.21789, 30.23763, 
    30.2572, 30.27659, 30.29582, 30.31488, 30.33376, 30.35247, 30.37102, 
    30.38939, 30.40758, 30.42561, 30.44346, 30.46114, 30.47865, 30.49599, 
    30.51315, 30.53014, 30.54696, 30.5636, 30.58007, 30.59637, 30.61249, 
    30.62844, 30.64421, 30.65981, 30.67524, 30.69049, 30.70557, 30.72047, 
    30.7352, 30.74975, 30.76413, 30.77833, 30.79236, 30.80621, 30.81989, 
    30.83339, 30.84671, 30.85986, 30.87283, 30.88562, 30.89824, 30.91069, 
    30.92295, 30.93504, 30.94695, 30.95869, 30.97025, 30.98163, 30.99283, 
    31.00386, 31.01471, 31.02538, 31.03587, 31.04619, 31.05633, 31.06629, 
    31.07607, 31.08567, 31.0951, 31.10435, 31.11342, 31.12231, 31.13102, 
    31.13955, 31.14791, 31.15608, 31.16408, 31.1719, 31.17954, 31.187, 
    31.19428, 31.20138, 31.2083, 31.21505, 31.22161, 31.22799, 31.2342, 
    31.24022, 31.24607, 31.25173, 31.25722, 31.26253, 31.26765, 31.2726, 
    31.27736, 31.28195, 31.28636, 31.29058, 31.29463, 31.29849, 31.30218, 
    31.30568, 31.30901, 31.31215, 31.31512, 31.3179, 31.32051, 31.32293, 
    31.32517, 31.32723, 31.32911, 31.33081, 31.33233, 31.33368, 31.33484, 
    31.33581, 31.33661, 31.33723, 31.33767, 31.33792, 31.338, 31.33789, 
    31.33761, 31.33714, 31.3365, 31.33567, 31.33466, 31.33348, 31.33211, 
    31.33056, 31.32883, 31.32692, 31.32483, 31.32256, 31.3201, 31.31747, 
    31.31466, 31.31167, 31.30849, 31.30514, 31.30161, 31.29789, 31.294, 
    31.28992, 31.28567, 31.28124, 31.27662, 31.27183, 31.26685, 31.2617, 
    31.25636, 31.25085, 31.24516, 31.23928, 31.23323, 31.227, 31.22058, 
    31.21399, 31.20722, 31.20027, 31.19314, 31.18583, 31.17834, 31.17068, 
    31.16283, 31.1548, 31.1466, 31.13822, 31.12965, 31.12091, 31.112, 
    31.1029, 31.09362, 31.08417, 31.07454, 31.06472, 31.05474, 31.04457, 
    31.03423, 31.0237, 31.013, 31.00213, 30.99107, 30.97984, 30.96843, 
    30.95684, 30.94508, 30.93314, 30.92102, 30.90873, 30.89626, 30.88361, 
    30.87079, 30.85779, 30.84461, 30.83126, 30.81773, 30.80403, 30.79015, 
    30.7761, 30.76187, 30.74746, 30.73288, 30.71813, 30.7032, 30.68809, 
    30.67281, 30.65736, 30.64173, 30.62593, 30.60995, 30.5938, 30.57748, 
    30.56098, 30.54431, 30.52746, 30.51045, 30.49326, 30.47589, 30.45836, 
    30.44065, 30.42277, 30.40471, 30.38649, 30.36809, 30.34953, 30.33078, 
    30.31187, 30.29279, 30.27354, 30.25411, 30.23452, 30.21475, 30.19481, 
    30.17471, 30.15443, 30.13398, 30.11337, 30.09258, 30.07163, 30.0505, 
    30.02921, 30.00775, 29.98612, 29.96432, 29.94235, 29.92022, 29.89791, 
    29.87544, 29.85281, 29.83, 29.80703, 29.78389, 29.76059, 29.73711, 
    29.71348, 29.68967, 29.6657, 29.64157, 29.61726, 29.5928, 29.56817, 
    29.54337, 29.51841, 29.49328, 29.46799, 29.44254, 29.41692, 29.39114, 
    29.3652, 29.33909, 29.31282, 29.28639, 29.25979, 29.23304, 29.20612, 
    29.17903, 29.15179, 29.12439, 29.09682, 29.06909, 29.04121, 29.01316, 
    28.98495, 28.95658, 28.92805, 28.89937, 28.87052, 28.84151, 28.81235, 
    28.78303, 28.75355,
  25.4609, 25.50404, 25.54705, 25.58993, 25.63267, 25.67527, 25.71774, 
    25.76008, 25.80228, 25.84434, 25.88626, 25.92805, 25.96971, 26.01122, 
    26.0526, 26.09384, 26.13494, 26.17591, 26.21673, 26.25741, 26.29796, 
    26.33837, 26.37864, 26.41876, 26.45875, 26.4986, 26.5383, 26.57787, 
    26.61729, 26.65657, 26.69571, 26.7347, 26.77356, 26.81227, 26.85084, 
    26.88927, 26.92755, 26.96568, 27.00368, 27.04153, 27.07923, 27.11679, 
    27.15421, 27.19147, 27.2286, 27.26558, 27.30241, 27.33909, 27.37563, 
    27.41202, 27.44826, 27.48436, 27.5203, 27.5561, 27.59175, 27.62726, 
    27.66261, 27.69781, 27.73287, 27.76778, 27.80253, 27.83714, 27.87159, 
    27.9059, 27.94005, 27.97405, 28.0079, 28.0416, 28.07514, 28.10854, 
    28.14178, 28.17487, 28.2078, 28.24059, 28.27321, 28.30569, 28.33801, 
    28.37018, 28.40219, 28.43405, 28.46575, 28.4973, 28.52869, 28.55993, 
    28.59101, 28.62193, 28.65269, 28.68331, 28.71376, 28.74405, 28.77419, 
    28.80417, 28.834, 28.86366, 28.89317, 28.92252, 28.95171, 28.98074, 
    29.00961, 29.03832, 29.06687, 29.09526, 29.12349, 29.15156, 29.17947, 
    29.20722, 29.2348, 29.26223, 29.2895, 29.3166, 29.34354, 29.37032, 
    29.39693, 29.42338, 29.44967, 29.4758, 29.50176, 29.52756, 29.5532, 
    29.57867, 29.60398, 29.62912, 29.6541, 29.67891, 29.70356, 29.72804, 
    29.75236, 29.77651, 29.8005, 29.82432, 29.84797, 29.87146, 29.89478, 
    29.91793, 29.94091, 29.96373, 29.98638, 30.00887, 30.03118, 30.05333, 
    30.07531, 30.09712, 30.11876, 30.14023, 30.16154, 30.18267, 30.20364, 
    30.22443, 30.24506, 30.26551, 30.2858, 30.30591, 30.32586, 30.34563, 
    30.36524, 30.38467, 30.40393, 30.42302, 30.44194, 30.46068, 30.47926, 
    30.49766, 30.51589, 30.53395, 30.55183, 30.56955, 30.58709, 30.60445, 
    30.62165, 30.63867, 30.65552, 30.67219, 30.68869, 30.70502, 30.72117, 
    30.73714, 30.75295, 30.76858, 30.78403, 30.79931, 30.81441, 30.82934, 
    30.8441, 30.85868, 30.87308, 30.88731, 30.90136, 30.91524, 30.92894, 
    30.94246, 30.95581, 30.96898, 30.98198, 30.99479, 31.00744, 31.0199, 
    31.03219, 31.0443, 31.05624, 31.06799, 31.07957, 31.09097, 31.1022, 
    31.11325, 31.12411, 31.13481, 31.14532, 31.15565, 31.16581, 31.17579, 
    31.18559, 31.19521, 31.20465, 31.21392, 31.223, 31.23191, 31.24064, 
    31.24919, 31.25756, 31.26575, 31.27376, 31.28159, 31.28925, 31.29672, 
    31.30401, 31.31113, 31.31807, 31.32482, 31.3314, 31.33779, 31.34401, 
    31.35004, 31.3559, 31.36158, 31.36707, 31.37239, 31.37752, 31.38248, 
    31.38725, 31.39185, 31.39626, 31.40049, 31.40455, 31.40842, 31.41211, 
    31.41562, 31.41895, 31.42211, 31.42508, 31.42786, 31.43047, 31.4329, 
    31.43515, 31.43721, 31.4391, 31.4408, 31.44233, 31.44367, 31.44483, 
    31.44581, 31.44661, 31.44723, 31.44767, 31.44792, 31.448, 31.4479, 
    31.44761, 31.44714, 31.4465, 31.44567, 31.44466, 31.44347, 31.4421, 
    31.44054, 31.43881, 31.4369, 31.4348, 31.43253, 31.43007, 31.42743, 
    31.42462, 31.42162, 31.41844, 31.41508, 31.41154, 31.40782, 31.40392, 
    31.39984, 31.39557, 31.39113, 31.38651, 31.38171, 31.37672, 31.37156, 
    31.36621, 31.36069, 31.35498, 31.3491, 31.34304, 31.33679, 31.33037, 
    31.32376, 31.31698, 31.31002, 31.30287, 31.29555, 31.28805, 31.28037, 
    31.27251, 31.26447, 31.25625, 31.24785, 31.23927, 31.23051, 31.22158, 
    31.21247, 31.20317, 31.1937, 31.18405, 31.17422, 31.16422, 31.15403, 
    31.14367, 31.13313, 31.12241, 31.11151, 31.10044, 31.08918, 31.07775, 
    31.06614, 31.05436, 31.0424, 31.03026, 31.01794, 31.00545, 30.99278, 
    30.97993, 30.96691, 30.95371, 30.94033, 30.92678, 30.91305, 30.89915, 
    30.88507, 30.87081, 30.85638, 30.84178, 30.82699, 30.81204, 30.7969, 
    30.7816, 30.76612, 30.75046, 30.73463, 30.71862, 30.70244, 30.68609, 
    30.66956, 30.65286, 30.63599, 30.61894, 30.60172, 30.58432, 30.56676, 
    30.54902, 30.53111, 30.51302, 30.49476, 30.47633, 30.45773, 30.43896, 
    30.42001, 30.40089, 30.38161, 30.36215, 30.34252, 30.32272, 30.30274, 
    30.2826, 30.26229, 30.24181, 30.22115, 30.20033, 30.17934, 30.15818, 
    30.13685, 30.11535, 30.09368, 30.07184, 30.04984, 30.02766, 30.00532, 
    29.98281, 29.96013, 29.93729, 29.91428, 29.8911, 29.86775, 29.84424, 
    29.82056, 29.79671, 29.7727, 29.74852, 29.72418, 29.69967, 29.675, 
    29.65016, 29.62515, 29.59999, 29.57465, 29.54915, 29.52349, 29.49767, 
    29.47168, 29.44553, 29.41921, 29.39273, 29.36609, 29.33929, 29.31232, 
    29.28519, 29.2579, 29.23045, 29.20284, 29.17506, 29.14713, 29.11903, 
    29.09078, 29.06236, 29.03379, 29.00505, 28.97615, 28.9471, 28.91788, 
    28.88851, 28.85898,
  25.56091, 25.60411, 25.64719, 25.69013, 25.73293, 25.7756, 25.81814, 
    25.86054, 25.9028, 25.94493, 25.98692, 26.02877, 26.07049, 26.11207, 
    26.15351, 26.19481, 26.23598, 26.277, 26.31789, 26.35864, 26.39925, 
    26.43972, 26.48005, 26.52024, 26.56029, 26.60019, 26.63996, 26.67959, 
    26.71907, 26.75841, 26.79762, 26.83667, 26.87559, 26.91436, 26.95299, 
    26.99148, 27.02982, 27.06802, 27.10607, 27.14398, 27.18174, 27.21936, 
    27.25684, 27.29416, 27.33135, 27.36838, 27.40527, 27.44202, 27.47861, 
    27.51506, 27.55136, 27.58752, 27.62352, 27.65938, 27.69509, 27.73065, 
    27.76606, 27.80132, 27.83643, 27.87139, 27.90621, 27.94087, 27.97538, 
    28.00974, 28.04395, 28.078, 28.11191, 28.14566, 28.17926, 28.21271, 
    28.24601, 28.27915, 28.31214, 28.34498, 28.37766, 28.41019, 28.44257, 
    28.47479, 28.50685, 28.53876, 28.57052, 28.60212, 28.63356, 28.66485, 
    28.69598, 28.72696, 28.75777, 28.78844, 28.81894, 28.84929, 28.87948, 
    28.90951, 28.93938, 28.9691, 28.99865, 29.02805, 29.05729, 29.08637, 
    29.11529, 29.14405, 29.17265, 29.20109, 29.22936, 29.25748, 29.28544, 
    29.31323, 29.34087, 29.36834, 29.39565, 29.4228, 29.44979, 29.47661, 
    29.50327, 29.52977, 29.55611, 29.58228, 29.60829, 29.63413, 29.65981, 
    29.68533, 29.71068, 29.73586, 29.76088, 29.78574, 29.81043, 29.83496, 
    29.85932, 29.88351, 29.90754, 29.9314, 29.95509, 29.97862, 30.00198, 
    30.02518, 30.0482, 30.07106, 30.09375, 30.11627, 30.13863, 30.16081, 
    30.18283, 30.20468, 30.22636, 30.24787, 30.26921, 30.29038, 30.31139, 
    30.33222, 30.35288, 30.37337, 30.39369, 30.41385, 30.43382, 30.45363, 
    30.47327, 30.49274, 30.51204, 30.53116, 30.55011, 30.56889, 30.5875, 
    30.60593, 30.6242, 30.64229, 30.6602, 30.67795, 30.69552, 30.71292, 
    30.73014, 30.74719, 30.76407, 30.78078, 30.7973, 30.81366, 30.82984, 
    30.84585, 30.86168, 30.87733, 30.89282, 30.90812, 30.92326, 30.93821, 
    30.95299, 30.9676, 30.98203, 30.99628, 31.01036, 31.02426, 31.03799, 
    31.05153, 31.06491, 31.0781, 31.09112, 31.10396, 31.11663, 31.12912, 
    31.14143, 31.15356, 31.16552, 31.1773, 31.1889, 31.20032, 31.21156, 
    31.22263, 31.23352, 31.24423, 31.25476, 31.26512, 31.27529, 31.28529, 
    31.29511, 31.30474, 31.31421, 31.32349, 31.33259, 31.34151, 31.35026, 
    31.35882, 31.36721, 31.37541, 31.38344, 31.39129, 31.39895, 31.40644, 
    31.41375, 31.42088, 31.42783, 31.43459, 31.44118, 31.44759, 31.45382, 
    31.45986, 31.46573, 31.47142, 31.47692, 31.48225, 31.48739, 31.49236, 
    31.49714, 31.50174, 31.50616, 31.51041, 31.51447, 31.51835, 31.52205, 
    31.52556, 31.5289, 31.53206, 31.53503, 31.53783, 31.54044, 31.54287, 
    31.54512, 31.54719, 31.54908, 31.55079, 31.55231, 31.55366, 31.55482, 
    31.55581, 31.55661, 31.55723, 31.55766, 31.55792, 31.558, 31.55789, 
    31.55761, 31.55714, 31.55649, 31.55566, 31.55465, 31.55346, 31.55208, 
    31.55053, 31.54879, 31.54688, 31.54478, 31.5425, 31.54004, 31.5374, 
    31.53457, 31.53157, 31.52839, 31.52502, 31.52147, 31.51775, 31.51384, 
    31.50975, 31.50548, 31.50103, 31.4964, 31.49158, 31.48659, 31.48142, 
    31.47606, 31.47053, 31.46481, 31.45892, 31.45284, 31.44659, 31.44015, 
    31.43353, 31.42674, 31.41976, 31.41261, 31.40527, 31.39775, 31.39006, 
    31.38218, 31.37413, 31.36589, 31.35748, 31.34889, 31.34011, 31.33116, 
    31.32203, 31.31272, 31.30323, 31.29357, 31.28372, 31.27369, 31.26349, 
    31.25311, 31.24255, 31.23181, 31.22089, 31.2098, 31.19852, 31.18707, 
    31.17544, 31.16364, 31.15165, 31.13949, 31.12715, 31.11464, 31.10194, 
    31.08908, 31.07603, 31.0628, 31.0494, 31.03583, 31.02207, 31.00814, 
    30.99404, 30.97976, 30.9653, 30.95067, 30.93586, 30.92087, 30.90571, 
    30.89038, 30.87487, 30.85919, 30.84333, 30.82729, 30.81108, 30.7947, 
    30.77814, 30.76141, 30.74451, 30.72743, 30.71018, 30.69275, 30.67515, 
    30.65738, 30.63944, 30.62132, 30.60303, 30.58457, 30.56593, 30.54712, 
    30.52814, 30.509, 30.48967, 30.47018, 30.45051, 30.43068, 30.41067, 
    30.39049, 30.37014, 30.34962, 30.32893, 30.30807, 30.28705, 30.26585, 
    30.24448, 30.22294, 30.20123, 30.17936, 30.15732, 30.1351, 30.11272, 
    30.09017, 30.06746, 30.04457, 30.02152, 29.9983, 29.97491, 29.95136, 
    29.92764, 29.90375, 29.87969, 29.85547, 29.83109, 29.80654, 29.78182, 
    29.75694, 29.73189, 29.70668, 29.6813, 29.65576, 29.63005, 29.60418, 
    29.57815, 29.55195, 29.52559, 29.49907, 29.47238, 29.44553, 29.41852, 
    29.39134, 29.36401, 29.33651, 29.30885, 29.28103, 29.25304, 29.2249, 
    29.1966, 29.16813, 29.13951, 29.11072, 29.08178, 29.05267, 29.02341, 
    28.99399, 28.96441,
  25.6609, 25.70417, 25.74731, 25.79032, 25.83319, 25.87592, 25.91852, 
    25.96099, 26.00331, 26.0455, 26.08756, 26.12947, 26.17125, 26.2129, 
    26.2544, 26.29577, 26.337, 26.37809, 26.41904, 26.45985, 26.50052, 
    26.54105, 26.58144, 26.62169, 26.66181, 26.70178, 26.74161, 26.78129, 
    26.82084, 26.86024, 26.89951, 26.93863, 26.9776, 27.01644, 27.05513, 
    27.09367, 27.13207, 27.17033, 27.20845, 27.24642, 27.28424, 27.32192, 
    27.35945, 27.39684, 27.43408, 27.47118, 27.50813, 27.54493, 27.58158, 
    27.61809, 27.65445, 27.69066, 27.72673, 27.76264, 27.79841, 27.83402, 
    27.86949, 27.90481, 27.93998, 27.975, 28.00987, 28.04459, 28.07915, 
    28.11357, 28.14783, 28.18195, 28.21591, 28.24972, 28.28337, 28.31688, 
    28.35023, 28.38343, 28.41647, 28.44936, 28.4821, 28.51468, 28.54711, 
    28.57938, 28.6115, 28.64347, 28.67527, 28.70692, 28.73842, 28.76976, 
    28.80095, 28.83197, 28.86284, 28.89356, 28.92411, 28.95451, 28.98475, 
    29.01483, 29.04476, 29.07452, 29.10413, 29.13357, 29.16286, 29.19199, 
    29.22096, 29.24977, 29.27842, 29.3069, 29.33523, 29.3634, 29.3914, 
    29.41924, 29.44693, 29.47445, 29.5018, 29.529, 29.55603, 29.5829, 
    29.60961, 29.63615, 29.66253, 29.68875, 29.7148, 29.74069, 29.76641, 
    29.79198, 29.81737, 29.8426, 29.86766, 29.89256, 29.9173, 29.94187, 
    29.96627, 29.9905, 30.01457, 30.03848, 30.06221, 30.08578, 30.10918, 
    30.13242, 30.15548, 30.17838, 30.20111, 30.22367, 30.24607, 30.26829, 
    30.29035, 30.31224, 30.33395, 30.3555, 30.37688, 30.39809, 30.41913, 
    30.44, 30.4607, 30.48123, 30.50159, 30.52177, 30.54179, 30.56163, 
    30.5813, 30.60081, 30.62014, 30.63929, 30.65828, 30.67709, 30.69573, 
    30.7142, 30.7325, 30.75062, 30.76857, 30.78635, 30.80395, 30.82138, 
    30.83863, 30.85572, 30.87262, 30.88936, 30.90592, 30.9223, 30.93851, 
    30.95455, 30.97041, 30.98609, 31.0016, 31.01694, 31.03209, 31.04708, 
    31.06189, 31.07652, 31.09097, 31.10525, 31.11936, 31.13328, 31.14703, 
    31.16061, 31.174, 31.18722, 31.20027, 31.21313, 31.22582, 31.23833, 
    31.25066, 31.26282, 31.2748, 31.2866, 31.29822, 31.30966, 31.32093, 
    31.33201, 31.34292, 31.35365, 31.3642, 31.37458, 31.38477, 31.39479, 
    31.40462, 31.41428, 31.42376, 31.43306, 31.44217, 31.45111, 31.45988, 
    31.46845, 31.47686, 31.48508, 31.49312, 31.50098, 31.50866, 31.51616, 
    31.52348, 31.53062, 31.53758, 31.54436, 31.55096, 31.55738, 31.56362, 
    31.56968, 31.57556, 31.58125, 31.58677, 31.59211, 31.59726, 31.60224, 
    31.60703, 31.61164, 31.61607, 31.62032, 31.62439, 31.62827, 31.63198, 
    31.6355, 31.63885, 31.64201, 31.64499, 31.64779, 31.65041, 31.65284, 
    31.6551, 31.65717, 31.65906, 31.66077, 31.6623, 31.66365, 31.66482, 
    31.6658, 31.6666, 31.66722, 31.66767, 31.66792, 31.668, 31.66789, 
    31.66761, 31.66714, 31.66649, 31.66566, 31.66464, 31.66345, 31.66207, 
    31.66052, 31.65878, 31.65686, 31.65475, 31.65247, 31.65001, 31.64736, 
    31.64453, 31.64152, 31.63833, 31.63496, 31.6314, 31.62767, 31.62375, 
    31.61966, 31.61538, 31.61092, 31.60628, 31.60146, 31.59646, 31.59127, 
    31.58591, 31.58037, 31.57464, 31.56874, 31.56265, 31.55638, 31.54993, 
    31.5433, 31.5365, 31.52951, 31.52234, 31.51499, 31.50746, 31.49975, 
    31.49186, 31.48379, 31.47554, 31.46711, 31.4585, 31.44971, 31.44074, 
    31.4316, 31.42227, 31.41276, 31.40308, 31.39321, 31.38317, 31.37295, 
    31.36255, 31.35197, 31.34121, 31.33027, 31.31916, 31.30786, 31.29639, 
    31.28474, 31.27291, 31.26091, 31.24872, 31.23636, 31.22382, 31.21111, 
    31.19821, 31.18514, 31.1719, 31.15847, 31.14487, 31.13109, 31.11714, 
    31.10301, 31.0887, 31.07421, 31.05956, 31.04472, 31.02971, 31.01452, 
    30.99916, 30.98362, 30.96791, 30.95202, 30.93596, 30.91972, 30.90331, 
    30.88672, 30.86996, 30.85303, 30.83592, 30.81863, 30.80118, 30.78355, 
    30.76574, 30.74776, 30.72962, 30.71129, 30.6928, 30.67413, 30.65529, 
    30.63627, 30.61709, 30.59773, 30.57821, 30.5585, 30.53863, 30.51859, 
    30.49837, 30.47799, 30.45744, 30.43671, 30.41581, 30.39475, 30.37351, 
    30.35211, 30.33053, 30.30878, 30.28687, 30.26479, 30.24254, 30.22012, 
    30.19753, 30.17477, 30.15184, 30.12875, 30.10549, 30.08206, 30.05847, 
    30.03471, 30.01078, 29.98668, 29.96242, 29.93799, 29.9134, 29.88864, 
    29.86371, 29.83862, 29.81336, 29.78794, 29.76236, 29.73661, 29.71069, 
    29.68461, 29.65837, 29.63196, 29.60539, 29.57866, 29.55177, 29.52471, 
    29.49749, 29.4701, 29.44256, 29.41485, 29.38698, 29.35895, 29.33076, 
    29.30241, 29.2739, 29.24522, 29.21639, 29.18739, 29.15824, 29.12893, 
    29.09945, 29.06982,
  25.76087, 25.80421, 25.84742, 25.89049, 25.93342, 25.97622, 26.01888, 
    26.06141, 26.1038, 26.14606, 26.18818, 26.23016, 26.272, 26.31371, 
    26.35528, 26.39671, 26.438, 26.47915, 26.52016, 26.56104, 26.60177, 
    26.64237, 26.68282, 26.72314, 26.76331, 26.80334, 26.84324, 26.88298, 
    26.92259, 26.96206, 27.00138, 27.04056, 27.0796, 27.11849, 27.15725, 
    27.19585, 27.23432, 27.27263, 27.31081, 27.34884, 27.38672, 27.42446, 
    27.46206, 27.4995, 27.5368, 27.57396, 27.61097, 27.64783, 27.68454, 
    27.72111, 27.75753, 27.79379, 27.82992, 27.86589, 27.90171, 27.93739, 
    27.97292, 28.00829, 28.04352, 28.07859, 28.11352, 28.14829, 28.18291, 
    28.21739, 28.25171, 28.28588, 28.31989, 28.35376, 28.38747, 28.42103, 
    28.45444, 28.48769, 28.52079, 28.55373, 28.58652, 28.61916, 28.65164, 
    28.68397, 28.71614, 28.74816, 28.78002, 28.81172, 28.84327, 28.87466, 
    28.9059, 28.93698, 28.9679, 28.99867, 29.02927, 29.05972, 29.09001, 
    29.12015, 29.15012, 29.17994, 29.20959, 29.23909, 29.26843, 29.2976, 
    29.32662, 29.35548, 29.38418, 29.41271, 29.44109, 29.4693, 29.49735, 
    29.52524, 29.55297, 29.58054, 29.60794, 29.63519, 29.66227, 29.68918, 
    29.71593, 29.74253, 29.76895, 29.79521, 29.82131, 29.84724, 29.87301, 
    29.89862, 29.92406, 29.94933, 29.97444, 29.99938, 30.02416, 30.04877, 
    30.07321, 30.09749, 30.1216, 30.14555, 30.16932, 30.19293, 30.21638, 
    30.23965, 30.26276, 30.2857, 30.30847, 30.33107, 30.3535, 30.37576, 
    30.39786, 30.41979, 30.44154, 30.46313, 30.48455, 30.50579, 30.52687, 
    30.54778, 30.56851, 30.58908, 30.60947, 30.62969, 30.64974, 30.66962, 
    30.68933, 30.70887, 30.72823, 30.74743, 30.76644, 30.78529, 30.80396, 
    30.82247, 30.8408, 30.85895, 30.87693, 30.89474, 30.91237, 30.92984, 
    30.94712, 30.96424, 30.98117, 30.99794, 31.01452, 31.03094, 31.04718, 
    31.06324, 31.07913, 31.09484, 31.11038, 31.12575, 31.14093, 31.15594, 
    31.17078, 31.18543, 31.19992, 31.21422, 31.22835, 31.2423, 31.25608, 
    31.26968, 31.2831, 31.29634, 31.30941, 31.3223, 31.33501, 31.34754, 
    31.3599, 31.37207, 31.38407, 31.3959, 31.40754, 31.419, 31.43029, 
    31.44139, 31.45232, 31.46307, 31.47364, 31.48404, 31.49425, 31.50428, 
    31.51414, 31.52381, 31.53331, 31.54262, 31.55176, 31.56071, 31.56949, 
    31.57809, 31.5865, 31.59474, 31.6028, 31.61067, 31.61837, 31.62588, 
    31.63322, 31.64037, 31.64734, 31.65414, 31.66075, 31.66718, 31.67343, 
    31.6795, 31.68539, 31.6911, 31.69662, 31.70197, 31.70713, 31.71211, 
    31.71692, 31.72153, 31.72597, 31.73023, 31.73431, 31.7382, 31.74191, 
    31.74544, 31.74879, 31.75196, 31.75495, 31.75775, 31.76037, 31.76282, 
    31.76508, 31.76715, 31.76905, 31.77076, 31.77229, 31.77364, 31.77481, 
    31.7758, 31.7766, 31.77722, 31.77766, 31.77792, 31.778, 31.77789, 
    31.77761, 31.77714, 31.77649, 31.77565, 31.77464, 31.77344, 31.77206, 
    31.7705, 31.76876, 31.76684, 31.76473, 31.76244, 31.75997, 31.75732, 
    31.75449, 31.75147, 31.74828, 31.7449, 31.74134, 31.7376, 31.73367, 
    31.72957, 31.72528, 31.72082, 31.71617, 31.71134, 31.70633, 31.70113, 
    31.69576, 31.6902, 31.68447, 31.67855, 31.67245, 31.66617, 31.65972, 
    31.65307, 31.64625, 31.63925, 31.63207, 31.62471, 31.61716, 31.60944, 
    31.60153, 31.59345, 31.58518, 31.57674, 31.56812, 31.55931, 31.55033, 
    31.54116, 31.53182, 31.52229, 31.51259, 31.50271, 31.49265, 31.4824, 
    31.47198, 31.46139, 31.45061, 31.43965, 31.42851, 31.4172, 31.40571, 
    31.39404, 31.38219, 31.37016, 31.35795, 31.34557, 31.33301, 31.32027, 
    31.30735, 31.29426, 31.28099, 31.26754, 31.25391, 31.24011, 31.22613, 
    31.21197, 31.19764, 31.18313, 31.16844, 31.15358, 31.13854, 31.12333, 
    31.10794, 31.09237, 31.07663, 31.06071, 31.04462, 31.02835, 31.01191, 
    30.9953, 30.9785, 30.96154, 30.9444, 30.92709, 30.9096, 30.89194, 
    30.8741, 30.85609, 30.83791, 30.81955, 30.80102, 30.78232, 30.76345, 
    30.7444, 30.72518, 30.70579, 30.68623, 30.66649, 30.64658, 30.6265, 
    30.60626, 30.58583, 30.56524, 30.54448, 30.52355, 30.50244, 30.48117, 
    30.45973, 30.43811, 30.41633, 30.39438, 30.37226, 30.34996, 30.32751, 
    30.30488, 30.28208, 30.25911, 30.23598, 30.21268, 30.18921, 30.16557, 
    30.14177, 30.1178, 30.09366, 30.06936, 30.04489, 30.02025, 29.99545, 
    29.97048, 29.94534, 29.92004, 29.89458, 29.86895, 29.84315, 29.81719, 
    29.79107, 29.76478, 29.73833, 29.71171, 29.68493, 29.65799, 29.63089, 
    29.60362, 29.57619, 29.5486, 29.52084, 29.49293, 29.46485, 29.43661, 
    29.40821, 29.37965, 29.35093, 29.32204, 29.293, 29.2638, 29.23443, 
    29.20491, 29.17523,
  25.86083, 25.90423, 25.9475, 25.99064, 26.03364, 26.0765, 26.11923, 
    26.16182, 26.20428, 26.2466, 26.28878, 26.33083, 26.37273, 26.41451, 
    26.45614, 26.49763, 26.53898, 26.5802, 26.62128, 26.66222, 26.70301, 
    26.74367, 26.78419, 26.82456, 26.8648, 26.9049, 26.94485, 26.98466, 
    27.02433, 27.06386, 27.10324, 27.14248, 27.18158, 27.22054, 27.25935, 
    27.29802, 27.33654, 27.37492, 27.41316, 27.45125, 27.48919, 27.52699, 
    27.56464, 27.60215, 27.63951, 27.67673, 27.71379, 27.75071, 27.78749, 
    27.82411, 27.86059, 27.89692, 27.93309, 27.96913, 28.00501, 28.04074, 
    28.07632, 28.11176, 28.14704, 28.18217, 28.21716, 28.25199, 28.28666, 
    28.32119, 28.35557, 28.3898, 28.42387, 28.45779, 28.49156, 28.52517, 
    28.55863, 28.59194, 28.62509, 28.65809, 28.69094, 28.72363, 28.75616, 
    28.78854, 28.82077, 28.85284, 28.88475, 28.91651, 28.94811, 28.97956, 
    29.01085, 29.04198, 29.07295, 29.10377, 29.13442, 29.16492, 29.19527, 
    29.22545, 29.25548, 29.28534, 29.31505, 29.34459, 29.37398, 29.40321, 
    29.43228, 29.46118, 29.48993, 29.51851, 29.54694, 29.5752, 29.6033, 
    29.63124, 29.65901, 29.68663, 29.71408, 29.74137, 29.76849, 29.79546, 
    29.82225, 29.84889, 29.87536, 29.90167, 29.92781, 29.95379, 29.9796, 
    30.00525, 30.03073, 30.05605, 30.0812, 30.10619, 30.13101, 30.15566, 
    30.18015, 30.20447, 30.22862, 30.25261, 30.27643, 30.30008, 30.32356, 
    30.34688, 30.37003, 30.39301, 30.41582, 30.43846, 30.46093, 30.48323, 
    30.50537, 30.52733, 30.54913, 30.57075, 30.59221, 30.61349, 30.63461, 
    30.65555, 30.67632, 30.69692, 30.71735, 30.73761, 30.7577, 30.77761, 
    30.79736, 30.81693, 30.83632, 30.85555, 30.87461, 30.89349, 30.91219, 
    30.93073, 30.94909, 30.96728, 30.98529, 31.00313, 31.0208, 31.03829, 
    31.05561, 31.07275, 31.08972, 31.10651, 31.12313, 31.13957, 31.15584, 
    31.17194, 31.18785, 31.2036, 31.21916, 31.23455, 31.24977, 31.2648, 
    31.27966, 31.29435, 31.30886, 31.32319, 31.33734, 31.35132, 31.36512, 
    31.37874, 31.39219, 31.40546, 31.41855, 31.43146, 31.44419, 31.45675, 
    31.46913, 31.48133, 31.49335, 31.50519, 31.51686, 31.52834, 31.53965, 
    31.55078, 31.56172, 31.57249, 31.58308, 31.59349, 31.60373, 31.61378, 
    31.62365, 31.63334, 31.64286, 31.65219, 31.66134, 31.67031, 31.67911, 
    31.68772, 31.69615, 31.7044, 31.71247, 31.72036, 31.72807, 31.7356, 
    31.74295, 31.75012, 31.7571, 31.76391, 31.77053, 31.77698, 31.78324, 
    31.78932, 31.79522, 31.80094, 31.80647, 31.81183, 31.817, 31.82199, 
    31.8268, 31.83143, 31.83588, 31.84014, 31.84422, 31.84813, 31.85185, 
    31.85538, 31.85874, 31.86191, 31.8649, 31.86771, 31.87034, 31.87279, 
    31.87505, 31.87713, 31.87903, 31.88075, 31.88228, 31.88363, 31.88481, 
    31.88579, 31.8866, 31.88722, 31.88766, 31.88792, 31.888, 31.88789, 
    31.88761, 31.88714, 31.88648, 31.88565, 31.88463, 31.88343, 31.88205, 
    31.88049, 31.87874, 31.87682, 31.8747, 31.87241, 31.86994, 31.86728, 
    31.86444, 31.86142, 31.85822, 31.85484, 31.85127, 31.84752, 31.84359, 
    31.83948, 31.83519, 31.83071, 31.82605, 31.82121, 31.81619, 31.81099, 
    31.80561, 31.80004, 31.7943, 31.78837, 31.78226, 31.77597, 31.7695, 
    31.76284, 31.75601, 31.74899, 31.7418, 31.73442, 31.72687, 31.71913, 
    31.71121, 31.70311, 31.69483, 31.68637, 31.67773, 31.66891, 31.65991, 
    31.65072, 31.64136, 31.63182, 31.6221, 31.6122, 31.60212, 31.59186, 
    31.58142, 31.5708, 31.56001, 31.54903, 31.53787, 31.52654, 31.51502, 
    31.50333, 31.49146, 31.47941, 31.46718, 31.45477, 31.44219, 31.42943, 
    31.41649, 31.40337, 31.39007, 31.3766, 31.36295, 31.34912, 31.33512, 
    31.32093, 31.30657, 31.29204, 31.27732, 31.26244, 31.24737, 31.23213, 
    31.21671, 31.20112, 31.18535, 31.1694, 31.15328, 31.13699, 31.12051, 
    31.10387, 31.08705, 31.07005, 31.05288, 31.03553, 31.01801, 31.00032, 
    30.98245, 30.96441, 30.9462, 30.92781, 30.90924, 30.89051, 30.8716, 
    30.85252, 30.83327, 30.81384, 30.79424, 30.77447, 30.75453, 30.73442, 
    30.71413, 30.69367, 30.67305, 30.65225, 30.63128, 30.61014, 30.58882, 
    30.56734, 30.54569, 30.52387, 30.50188, 30.47972, 30.45739, 30.43489, 
    30.41222, 30.38938, 30.36638, 30.3432, 30.31986, 30.29635, 30.27267, 
    30.24883, 30.22481, 30.20063, 30.17629, 30.15177, 30.12709, 30.10225, 
    30.07724, 30.05206, 30.02671, 30.0012, 29.97553, 29.94969, 29.92369, 
    29.89752, 29.87118, 29.84469, 29.81803, 29.7912, 29.76421, 29.73706, 
    29.70975, 29.68227, 29.65463, 29.62683, 29.59886, 29.57074, 29.54245, 
    29.514, 29.48539, 29.45662, 29.42769, 29.3986, 29.36934, 29.33993, 
    29.31036, 29.28063,
  25.96077, 26.00424, 26.04757, 26.09077, 26.13384, 26.17677, 26.21956, 
    26.26222, 26.30474, 26.34712, 26.38937, 26.43148, 26.47345, 26.51528, 
    26.55698, 26.59854, 26.63996, 26.68123, 26.72237, 26.76337, 26.80424, 
    26.84496, 26.88554, 26.92598, 26.96627, 27.00643, 27.04645, 27.08632, 
    27.12605, 27.16564, 27.20509, 27.24439, 27.28355, 27.32257, 27.36144, 
    27.40017, 27.43876, 27.4772, 27.51549, 27.55364, 27.59165, 27.62951, 
    27.66722, 27.70478, 27.7422, 27.77948, 27.8166, 27.85358, 27.89042, 
    27.9271, 27.96363, 28.00002, 28.03626, 28.07235, 28.10829, 28.14408, 
    28.17972, 28.21521, 28.25055, 28.28574, 28.32078, 28.35567, 28.3904, 
    28.42499, 28.45942, 28.4937, 28.52783, 28.56181, 28.59563, 28.6293, 
    28.66281, 28.69618, 28.72938, 28.76244, 28.79534, 28.82808, 28.86067, 
    28.89311, 28.92539, 28.95751, 28.98948, 29.02129, 29.05294, 29.08444, 
    29.11578, 29.14696, 29.17799, 29.20886, 29.23957, 29.27012, 29.30051, 
    29.33075, 29.36082, 29.39074, 29.42049, 29.45009, 29.47953, 29.5088, 
    29.53792, 29.56688, 29.59567, 29.6243, 29.65277, 29.68109, 29.70923, 
    29.73722, 29.76504, 29.79271, 29.8202, 29.84754, 29.87471, 29.90172, 
    29.92857, 29.95525, 29.98176, 30.00812, 30.0343, 30.06033, 30.08619, 
    30.11188, 30.13741, 30.16277, 30.18796, 30.21299, 30.23785, 30.26255, 
    30.28708, 30.31144, 30.33564, 30.35967, 30.38353, 30.40722, 30.43074, 
    30.4541, 30.47729, 30.50031, 30.52316, 30.54584, 30.56835, 30.5907, 
    30.61287, 30.63487, 30.65671, 30.67837, 30.69986, 30.72118, 30.74233, 
    30.76332, 30.78412, 30.80476, 30.82523, 30.84552, 30.86564, 30.8856, 
    30.90537, 30.92498, 30.94441, 30.96367, 30.98276, 31.00167, 31.02042, 
    31.03898, 31.05738, 31.0756, 31.09365, 31.11152, 31.12922, 31.14674, 
    31.16409, 31.18126, 31.19826, 31.21508, 31.23173, 31.24821, 31.2645, 
    31.28063, 31.29657, 31.31234, 31.32794, 31.34336, 31.3586, 31.37366, 
    31.38855, 31.40326, 31.4178, 31.43215, 31.44633, 31.46034, 31.47416, 
    31.48781, 31.50128, 31.51457, 31.52769, 31.54062, 31.55338, 31.56596, 
    31.57836, 31.59058, 31.60262, 31.61449, 31.62617, 31.63768, 31.64901, 
    31.66015, 31.67112, 31.68191, 31.69252, 31.70295, 31.7132, 31.72327, 
    31.73316, 31.74287, 31.7524, 31.76175, 31.77092, 31.77991, 31.78872, 
    31.79735, 31.8058, 31.81406, 31.82215, 31.83005, 31.83778, 31.84532, 
    31.85268, 31.85986, 31.86686, 31.87368, 31.88032, 31.88677, 31.89304, 
    31.89914, 31.90504, 31.91077, 31.91632, 31.92169, 31.92687, 31.93187, 
    31.93669, 31.94133, 31.94578, 31.95005, 31.95414, 31.95805, 31.96178, 
    31.96532, 31.96869, 31.97186, 31.97486, 31.97768, 31.98031, 31.98276, 
    31.98503, 31.98711, 31.98901, 31.99073, 31.99227, 31.99363, 31.9948, 
    31.99579, 31.9966, 31.99722, 31.99766, 31.99792, 31.998, 31.99789, 
    31.99761, 31.99714, 31.99648, 31.99565, 31.99463, 31.99343, 31.99204, 
    31.99047, 31.98873, 31.98679, 31.98468, 31.98238, 31.97991, 31.97724, 
    31.9744, 31.97137, 31.96817, 31.96478, 31.9612, 31.95745, 31.95351, 
    31.94939, 31.94509, 31.9406, 31.93594, 31.93109, 31.92606, 31.92085, 
    31.91545, 31.90988, 31.90412, 31.89818, 31.89206, 31.88576, 31.87928, 
    31.87261, 31.86577, 31.85874, 31.85153, 31.84414, 31.83657, 31.82882, 
    31.82088, 31.81277, 31.80447, 31.796, 31.78734, 31.7785, 31.76949, 
    31.76029, 31.75091, 31.74135, 31.73161, 31.72169, 31.71159, 31.70131, 
    31.69086, 31.68022, 31.6694, 31.6584, 31.64723, 31.63587, 31.62434, 
    31.61262, 31.60073, 31.58866, 31.57641, 31.56398, 31.55137, 31.53859, 
    31.52562, 31.51248, 31.49916, 31.48566, 31.47199, 31.45813, 31.4441, 
    31.42989, 31.41551, 31.40095, 31.38621, 31.37129, 31.3562, 31.34093, 
    31.32548, 31.30986, 31.29406, 31.27809, 31.26194, 31.24561, 31.22911, 
    31.21243, 31.19558, 31.17856, 31.16135, 31.14398, 31.12643, 31.1087, 
    31.0908, 31.07273, 31.05448, 31.03606, 31.01746, 30.9987, 30.97975, 
    30.96064, 30.94135, 30.92189, 30.90226, 30.88245, 30.86247, 30.84232, 
    30.822, 30.80151, 30.78084, 30.76001, 30.739, 30.71782, 30.69647, 
    30.67495, 30.65326, 30.6314, 30.60937, 30.58717, 30.5648, 30.54226, 
    30.51956, 30.49668, 30.47363, 30.45042, 30.42703, 30.40348, 30.37976, 
    30.35588, 30.33182, 30.3076, 30.28321, 30.25866, 30.23393, 30.20904, 
    30.18399, 30.15877, 30.13338, 30.10782, 30.08211, 30.05622, 30.03017, 
    30.00396, 29.97758, 29.95104, 29.92433, 29.89746, 29.87042, 29.84323, 
    29.81586, 29.78834, 29.76065, 29.7328, 29.70479, 29.67662, 29.64828, 
    29.61978, 29.59113, 29.56231, 29.53333, 29.50418, 29.47488, 29.44542, 
    29.4158, 29.38601,
  26.06069, 26.10423, 26.14762, 26.19089, 26.23402, 26.27701, 26.31987, 
    26.36259, 26.40518, 26.44763, 26.48994, 26.53211, 26.57415, 26.61604, 
    26.6578, 26.69942, 26.74091, 26.78225, 26.82345, 26.86452, 26.90544, 
    26.94623, 26.98687, 27.02737, 27.06773, 27.10795, 27.14803, 27.18797, 
    27.22776, 27.26741, 27.30692, 27.34628, 27.38551, 27.42458, 27.46352, 
    27.50231, 27.54095, 27.57945, 27.61781, 27.65602, 27.69409, 27.732, 
    27.76978, 27.8074, 27.84488, 27.88222, 27.9194, 27.95644, 27.99333, 
    28.03007, 28.06667, 28.10311, 28.13941, 28.17556, 28.21156, 28.2474, 
    28.2831, 28.31865, 28.35405, 28.38929, 28.42439, 28.45934, 28.49413, 
    28.52877, 28.56326, 28.5976, 28.63178, 28.66581, 28.69969, 28.73341, 
    28.76698, 28.8004, 28.83367, 28.86677, 28.89973, 28.93253, 28.96517, 
    28.99766, 29.02999, 29.06217, 29.09419, 29.12605, 29.15776, 29.18931, 
    29.2207, 29.25194, 29.28302, 29.31394, 29.3447, 29.3753, 29.40574, 
    29.43603, 29.46616, 29.49612, 29.52593, 29.55558, 29.58506, 29.61439, 
    29.64355, 29.67256, 29.7014, 29.73009, 29.75861, 29.78696, 29.81516, 
    29.84319, 29.87107, 29.89878, 29.92632, 29.9537, 29.98092, 30.00798, 
    30.03487, 30.0616, 30.08816, 30.11456, 30.14079, 30.16686, 30.19276, 
    30.2185, 30.24407, 30.26947, 30.29471, 30.31979, 30.34469, 30.36943, 
    30.394, 30.41841, 30.44265, 30.46672, 30.49062, 30.51435, 30.53792, 
    30.56132, 30.58455, 30.60761, 30.6305, 30.65322, 30.67577, 30.69815, 
    30.72036, 30.74241, 30.76428, 30.78598, 30.80751, 30.82887, 30.85006, 
    30.87108, 30.89192, 30.9126, 30.9331, 30.95343, 30.97359, 30.99357, 
    31.01339, 31.03303, 31.0525, 31.07179, 31.09091, 31.10986, 31.12864, 
    31.14724, 31.16566, 31.18392, 31.202, 31.2199, 31.23763, 31.25518, 
    31.27256, 31.28977, 31.3068, 31.32365, 31.34033, 31.35683, 31.37316, 
    31.38931, 31.40529, 31.42109, 31.43671, 31.45216, 31.46742, 31.48252, 
    31.49743, 31.51217, 31.52673, 31.54111, 31.55532, 31.56935, 31.5832, 
    31.59687, 31.61036, 31.62368, 31.63682, 31.64978, 31.66256, 31.67516, 
    31.68759, 31.69983, 31.71189, 31.72378, 31.73549, 31.74702, 31.75836, 
    31.76953, 31.78052, 31.79133, 31.80196, 31.81241, 31.82268, 31.83277, 
    31.84267, 31.8524, 31.86195, 31.87132, 31.8805, 31.88951, 31.89833, 
    31.90698, 31.91544, 31.92372, 31.93182, 31.93974, 31.94748, 31.95504, 
    31.96241, 31.96961, 31.97662, 31.98345, 31.9901, 31.99656, 32.00285, 
    32.00895, 32.01487, 32.02061, 32.02617, 32.03154, 32.03674, 32.04175, 
    32.04657, 32.05122, 32.05568, 32.05996, 32.06406, 32.06798, 32.07171, 
    32.07526, 32.07863, 32.08182, 32.08482, 32.08764, 32.09027, 32.09273, 
    32.095, 32.09709, 32.099, 32.10072, 32.10226, 32.10362, 32.10479, 
    32.10579, 32.10659, 32.10722, 32.10766, 32.10792, 32.108, 32.10789, 
    32.1076, 32.10713, 32.10648, 32.10564, 32.10462, 32.10342, 32.10203, 
    32.10046, 32.09871, 32.09678, 32.09465, 32.09235, 32.08987, 32.0872, 
    32.08436, 32.08133, 32.07811, 32.07471, 32.07113, 32.06737, 32.06343, 
    32.0593, 32.05499, 32.0505, 32.04582, 32.04097, 32.03593, 32.0307, 
    32.0253, 32.01972, 32.01395, 32.008, 32.00187, 31.99555, 31.98906, 
    31.98238, 31.97552, 31.96848, 31.96126, 31.95385, 31.94627, 31.9385, 
    31.93055, 31.92242, 31.91411, 31.90562, 31.89695, 31.8881, 31.87906, 
    31.86985, 31.86045, 31.85088, 31.84112, 31.83118, 31.82107, 31.81077, 
    31.80029, 31.78963, 31.7788, 31.76778, 31.75658, 31.7452, 31.73365, 
    31.72191, 31.71, 31.6979, 31.68563, 31.67318, 31.66055, 31.64774, 
    31.63475, 31.62159, 31.60824, 31.59472, 31.58102, 31.56714, 31.55309, 
    31.53885, 31.52444, 31.50985, 31.49508, 31.48014, 31.46502, 31.44972, 
    31.43425, 31.4186, 31.40277, 31.38677, 31.37059, 31.35424, 31.33771, 
    31.321, 31.30412, 31.28706, 31.26983, 31.25242, 31.23484, 31.21708, 
    31.19915, 31.18104, 31.16276, 31.14431, 31.12568, 31.10688, 31.0879, 
    31.06875, 31.04943, 31.02993, 31.01027, 30.99043, 30.97041, 30.95023, 
    30.92987, 30.90934, 30.88864, 30.86776, 30.84672, 30.8255, 30.80412, 
    30.78256, 30.76083, 30.73893, 30.71686, 30.69462, 30.67221, 30.64964, 
    30.62689, 30.60397, 30.58088, 30.55763, 30.5342, 30.51061, 30.48685, 
    30.46292, 30.43883, 30.41456, 30.39013, 30.36553, 30.34076, 30.31583, 
    30.29073, 30.26547, 30.24003, 30.21444, 30.18867, 30.16274, 30.13665, 
    30.11039, 30.08397, 30.05738, 30.03062, 30.00371, 29.97663, 29.94938, 
    29.92197, 29.8944, 29.86667, 29.83877, 29.81071, 29.78249, 29.7541, 
    29.72556, 29.69685, 29.66798, 29.63895, 29.60976, 29.58041, 29.5509, 
    29.52122, 29.49139,
  26.16059, 26.20419, 26.24766, 26.29099, 26.33418, 26.37724, 26.42017, 
    26.46295, 26.5056, 26.54811, 26.59049, 26.63273, 26.67483, 26.71679, 
    26.75861, 26.8003, 26.84184, 26.88325, 26.92452, 26.96564, 27.00663, 
    27.04748, 27.08818, 27.12875, 27.16917, 27.20945, 27.2496, 27.28959, 
    27.32945, 27.36916, 27.40873, 27.44816, 27.48744, 27.52658, 27.56558, 
    27.60443, 27.64314, 27.6817, 27.72011, 27.75838, 27.79651, 27.83449, 
    27.87232, 27.91001, 27.94755, 27.98494, 28.02219, 28.05928, 28.09623, 
    28.13304, 28.16969, 28.20619, 28.24255, 28.27875, 28.31481, 28.35072, 
    28.38647, 28.42208, 28.45753, 28.49284, 28.52799, 28.56299, 28.59784, 
    28.63254, 28.66708, 28.70148, 28.73572, 28.7698, 28.80374, 28.83752, 
    28.87115, 28.90462, 28.93793, 28.9711, 29.00411, 29.03696, 29.06966, 
    29.1022, 29.13459, 29.16682, 29.19889, 29.23081, 29.26257, 29.29417, 
    29.32562, 29.3569, 29.38803, 29.419, 29.44982, 29.48047, 29.51097, 
    29.5413, 29.57148, 29.6015, 29.63136, 29.66105, 29.69059, 29.71996, 
    29.74918, 29.77823, 29.80713, 29.83586, 29.86443, 29.89283, 29.92108, 
    29.94916, 29.97708, 30.00484, 30.03243, 30.05986, 30.08712, 30.11423, 
    30.14116, 30.16794, 30.19454, 30.22099, 30.24727, 30.27338, 30.29933, 
    30.32511, 30.35073, 30.37617, 30.40146, 30.42657, 30.45152, 30.47631, 
    30.50092, 30.52537, 30.54965, 30.57376, 30.59771, 30.62148, 30.64509, 
    30.66853, 30.6918, 30.7149, 30.73783, 30.76059, 30.78318, 30.8056, 
    30.82785, 30.84994, 30.87185, 30.89359, 30.91515, 30.93655, 30.95778, 
    30.97883, 30.99972, 31.02043, 31.04097, 31.06133, 31.08153, 31.10155, 
    31.1214, 31.14107, 31.16058, 31.1799, 31.19906, 31.21804, 31.23685, 
    31.25549, 31.27395, 31.29223, 31.31034, 31.32828, 31.34604, 31.36363, 
    31.38104, 31.39827, 31.41533, 31.43222, 31.44893, 31.46546, 31.48182, 
    31.498, 31.514, 31.52983, 31.54548, 31.56095, 31.57625, 31.59137, 
    31.60631, 31.62108, 31.63566, 31.65007, 31.66431, 31.67836, 31.69224, 
    31.70593, 31.71945, 31.73279, 31.74595, 31.75894, 31.77174, 31.78437, 
    31.79681, 31.80908, 31.82117, 31.83307, 31.8448, 31.85635, 31.86772, 
    31.87891, 31.88992, 31.90075, 31.91139, 31.92186, 31.93215, 31.94226, 
    31.95218, 31.96193, 31.9715, 31.98088, 31.99008, 31.99911, 32.00795, 
    32.01661, 32.02509, 32.03338, 32.0415, 32.04943, 32.05718, 32.06475, 
    32.07214, 32.07935, 32.08638, 32.09322, 32.09988, 32.10636, 32.11266, 
    32.11877, 32.1247, 32.13045, 32.13602, 32.1414, 32.14661, 32.15162, 
    32.15646, 32.16111, 32.16559, 32.16988, 32.17398, 32.17791, 32.18164, 
    32.1852, 32.18858, 32.19177, 32.19477, 32.1976, 32.20024, 32.2027, 
    32.20498, 32.20707, 32.20898, 32.21071, 32.21225, 32.21361, 32.21479, 
    32.21578, 32.21659, 32.21722, 32.21766, 32.21792, 32.218, 32.21789, 
    32.21761, 32.21713, 32.21648, 32.21564, 32.21461, 32.21341, 32.21202, 
    32.21045, 32.20869, 32.20675, 32.20463, 32.20233, 32.19984, 32.19717, 
    32.19431, 32.19128, 32.18806, 32.18465, 32.18106, 32.1773, 32.17334, 
    32.16921, 32.16489, 32.16039, 32.15571, 32.15084, 32.14579, 32.14056, 
    32.13515, 32.12955, 32.12378, 32.11781, 32.11167, 32.10535, 32.09884, 
    32.09215, 32.08528, 32.07822, 32.07099, 32.06357, 32.05597, 32.04819, 
    32.04023, 32.03208, 32.02376, 32.01525, 32.00656, 31.99769, 31.98864, 
    31.97941, 31.97, 31.9604, 31.95063, 31.94067, 31.93054, 31.92022, 
    31.90972, 31.89905, 31.88819, 31.87715, 31.86593, 31.85454, 31.84296, 
    31.8312, 31.81927, 31.80715, 31.79486, 31.78238, 31.76973, 31.7569, 
    31.74388, 31.73069, 31.71733, 31.70378, 31.69005, 31.67615, 31.66207, 
    31.64781, 31.63337, 31.61875, 31.60396, 31.58899, 31.57384, 31.55852, 
    31.54302, 31.52734, 31.51148, 31.49545, 31.47924, 31.46286, 31.4463, 
    31.42956, 31.41265, 31.39556, 31.3783, 31.36086, 31.34324, 31.32545, 
    31.30749, 31.28935, 31.27104, 31.25255, 31.23389, 31.21505, 31.19604, 
    31.17686, 31.1575, 31.13797, 31.11827, 31.09839, 31.07834, 31.05812, 
    31.03773, 31.01716, 30.99642, 30.97551, 30.95443, 30.93318, 30.91175, 
    30.89016, 30.86839, 30.84645, 30.82434, 30.80207, 30.77962, 30.757, 
    30.73421, 30.71125, 30.68813, 30.66483, 30.64137, 30.61773, 30.59393, 
    30.56996, 30.54582, 30.52151, 30.49704, 30.4724, 30.44759, 30.42261, 
    30.39747, 30.37216, 30.34668, 30.32104, 30.29523, 30.26926, 30.24312, 
    30.21682, 30.19035, 30.16371, 30.13691, 30.10995, 30.08282, 30.05553, 
    30.02807, 30.00046, 29.97267, 29.94473, 29.91662, 29.88835, 29.85992, 
    29.83132, 29.80257, 29.77365, 29.74457, 29.71533, 29.68593, 29.65637, 
    29.62664, 29.59676,
  26.26048, 26.30414, 26.34768, 26.39107, 26.43433, 26.47745, 26.52044, 
    26.56329, 26.60601, 26.64858, 26.69102, 26.73333, 26.77549, 26.81752, 
    26.85941, 26.90115, 26.94276, 26.98423, 27.02556, 27.06675, 27.10781, 
    27.14871, 27.18948, 27.23011, 27.2706, 27.31094, 27.35114, 27.3912, 
    27.43112, 27.4709, 27.51053, 27.55002, 27.58937, 27.62856, 27.66762, 
    27.70654, 27.7453, 27.78393, 27.8224, 27.86073, 27.89892, 27.93696, 
    27.97485, 28.0126, 28.0502, 28.08765, 28.12496, 28.16211, 28.19912, 
    28.23598, 28.27269, 28.30926, 28.34567, 28.38193, 28.41805, 28.45401, 
    28.48983, 28.52549, 28.561, 28.59636, 28.63157, 28.66663, 28.70154, 
    28.73629, 28.7709, 28.80535, 28.83964, 28.87379, 28.90777, 28.94161, 
    28.97529, 29.00882, 29.04219, 29.07541, 29.10847, 29.14138, 29.17413, 
    29.20673, 29.23917, 29.27145, 29.30358, 29.33555, 29.36736, 29.39902, 
    29.43052, 29.46186, 29.49304, 29.52406, 29.55493, 29.58563, 29.61618, 
    29.64657, 29.6768, 29.70687, 29.73677, 29.76652, 29.79611, 29.82553, 
    29.8548, 29.8839, 29.91284, 29.94162, 29.97024, 29.9987, 30.02699, 
    30.05512, 30.08308, 30.11089, 30.13853, 30.166, 30.19332, 30.22047, 
    30.24745, 30.27427, 30.30092, 30.32741, 30.35374, 30.37989, 30.40589, 
    30.43171, 30.45737, 30.48287, 30.5082, 30.53336, 30.55835, 30.58317, 
    30.60783, 30.63232, 30.65664, 30.6808, 30.70479, 30.7286, 30.75225, 
    30.77573, 30.79904, 30.82218, 30.84515, 30.86795, 30.89059, 30.91305, 
    30.93534, 30.95746, 30.97941, 31.00118, 31.02279, 31.04423, 31.06549, 
    31.08658, 31.1075, 31.12825, 31.14883, 31.16923, 31.18946, 31.20952, 
    31.2294, 31.24911, 31.26865, 31.28802, 31.30721, 31.32622, 31.34506, 
    31.36373, 31.38222, 31.40054, 31.41869, 31.43666, 31.45445, 31.47206, 
    31.48951, 31.50677, 31.52387, 31.54078, 31.55752, 31.57408, 31.59047, 
    31.60668, 31.62271, 31.63857, 31.65425, 31.66975, 31.68507, 31.70022, 
    31.71519, 31.72998, 31.74459, 31.75903, 31.77329, 31.78737, 31.80127, 
    31.81499, 31.82854, 31.8419, 31.85509, 31.86809, 31.88092, 31.89357, 
    31.90604, 31.91833, 31.93044, 31.94236, 31.95411, 31.96568, 31.97707, 
    31.98828, 31.99931, 32.01016, 32.02083, 32.03131, 32.04162, 32.05175, 
    32.0617, 32.07146, 32.08104, 32.09044, 32.09966, 32.1087, 32.11756, 
    32.12624, 32.13473, 32.14304, 32.15117, 32.15912, 32.16689, 32.17447, 
    32.18187, 32.18909, 32.19613, 32.20299, 32.20966, 32.21615, 32.22246, 
    32.22858, 32.23453, 32.24029, 32.24586, 32.25126, 32.25647, 32.2615, 
    32.26635, 32.27101, 32.27549, 32.27979, 32.2839, 32.28783, 32.29158, 
    32.29514, 32.29852, 32.30172, 32.30473, 32.30756, 32.31021, 32.31268, 
    32.31495, 32.31705, 32.31897, 32.32069, 32.32224, 32.3236, 32.32478, 
    32.32578, 32.32659, 32.32722, 32.32766, 32.32792, 32.328, 32.32789, 
    32.3276, 32.32713, 32.32647, 32.32563, 32.32461, 32.3234, 32.32201, 
    32.32043, 32.31867, 32.31673, 32.31461, 32.3123, 32.3098, 32.30713, 
    32.30427, 32.30123, 32.298, 32.29459, 32.291, 32.28722, 32.28326, 
    32.27912, 32.27479, 32.27028, 32.26559, 32.26072, 32.25566, 32.25042, 
    32.245, 32.23939, 32.2336, 32.22763, 32.22147, 32.21514, 32.20862, 
    32.20192, 32.19503, 32.18797, 32.18071, 32.17328, 32.16567, 32.15788, 
    32.1499, 32.14174, 32.1334, 32.12487, 32.11617, 32.10728, 32.09822, 
    32.08897, 32.07954, 32.06993, 32.06013, 32.05016, 32.04, 32.02967, 
    32.01915, 32.00846, 31.99758, 31.98652, 31.97528, 31.96387, 31.95227, 
    31.94049, 31.92853, 31.91639, 31.90408, 31.89158, 31.8789, 31.86605, 
    31.85301, 31.8398, 31.8264, 31.81283, 31.79908, 31.78515, 31.77105, 
    31.75676, 31.7423, 31.72765, 31.71283, 31.69784, 31.68266, 31.66731, 
    31.65178, 31.63607, 31.62019, 31.60413, 31.58789, 31.57148, 31.55488, 
    31.53812, 31.52118, 31.50406, 31.48676, 31.46929, 31.45164, 31.43382, 
    31.41583, 31.39766, 31.37931, 31.36079, 31.34209, 31.32323, 31.30418, 
    31.28496, 31.26557, 31.24601, 31.22627, 31.20636, 31.18627, 31.16601, 
    31.14558, 31.12498, 31.10421, 31.08326, 31.06214, 31.04085, 31.01939, 
    30.99775, 30.97595, 30.95397, 30.93182, 30.90951, 30.88702, 30.86436, 
    30.84153, 30.81853, 30.79537, 30.77203, 30.74852, 30.72485, 30.701, 
    30.67699, 30.65281, 30.62846, 30.60394, 30.57926, 30.55441, 30.52939, 
    30.5042, 30.47885, 30.45333, 30.42764, 30.40179, 30.37577, 30.34958, 
    30.32323, 30.29672, 30.27004, 30.24319, 30.21618, 30.18901, 30.16167, 
    30.13417, 30.1065, 30.07867, 30.05068, 30.02252, 29.9942, 29.96572, 
    29.93708, 29.90827, 29.87931, 29.85018, 29.82089, 29.79144, 29.76183, 
    29.73205, 29.70212,
  26.36034, 26.40408, 26.44767, 26.49113, 26.53446, 26.57765, 26.6207, 
    26.66362, 26.7064, 26.74904, 26.79154, 26.83391, 26.87614, 26.91823, 
    26.96018, 27.00199, 27.04366, 27.0852, 27.12659, 27.16785, 27.20896, 
    27.24993, 27.29077, 27.33146, 27.37201, 27.41241, 27.45268, 27.4928, 
    27.53278, 27.57262, 27.61231, 27.65187, 27.69127, 27.73053, 27.76965, 
    27.80863, 27.84745, 27.88614, 27.92468, 27.96307, 28.00132, 28.03942, 
    28.07737, 28.11518, 28.15283, 28.19035, 28.22771, 28.26493, 28.302, 
    28.33891, 28.37568, 28.41231, 28.44878, 28.4851, 28.52127, 28.5573, 
    28.59317, 28.62889, 28.66446, 28.69988, 28.73515, 28.77026, 28.80523, 
    28.84004, 28.8747, 28.9092, 28.94355, 28.97775, 29.0118, 29.04569, 
    29.07943, 29.11301, 29.14644, 29.17971, 29.21283, 29.24579, 29.2786, 
    29.31125, 29.34374, 29.37608, 29.40826, 29.44028, 29.47215, 29.50386, 
    29.53541, 29.5668, 29.59804, 29.62911, 29.66003, 29.69079, 29.72138, 
    29.75182, 29.7821, 29.81222, 29.84218, 29.87198, 29.90161, 29.93109, 
    29.9604, 29.98956, 30.01855, 30.04738, 30.07604, 30.10455, 30.13289, 
    30.16107, 30.18908, 30.21693, 30.24462, 30.27214, 30.2995, 30.3267, 
    30.35373, 30.38059, 30.40729, 30.43383, 30.4602, 30.4864, 30.51244, 
    30.53831, 30.56402, 30.58955, 30.61493, 30.64013, 30.66516, 30.69003, 
    30.71474, 30.73927, 30.76363, 30.78783, 30.81186, 30.83572, 30.85941, 
    30.88293, 30.90628, 30.92946, 30.95247, 30.97532, 30.99799, 31.02049, 
    31.04282, 31.06498, 31.08696, 31.10878, 31.13042, 31.1519, 31.1732, 
    31.19433, 31.21529, 31.23607, 31.25668, 31.27712, 31.29739, 31.31748, 
    31.3374, 31.35715, 31.37672, 31.39612, 31.41534, 31.43439, 31.45327, 
    31.47197, 31.4905, 31.50885, 31.52703, 31.54502, 31.56285, 31.5805, 
    31.59797, 31.61527, 31.63239, 31.64934, 31.66611, 31.6827, 31.69912, 
    31.71536, 31.73142, 31.7473, 31.76301, 31.77854, 31.79389, 31.80907, 
    31.82406, 31.83888, 31.85352, 31.86798, 31.88227, 31.89637, 31.9103, 
    31.92405, 31.93761, 31.951, 31.96421, 31.97725, 31.9901, 32.00277, 
    32.01526, 32.02757, 32.0397, 32.05165, 32.06342, 32.07502, 32.08643, 
    32.09766, 32.10871, 32.11958, 32.13026, 32.14077, 32.15109, 32.16124, 
    32.1712, 32.18098, 32.19059, 32.2, 32.20924, 32.2183, 32.22717, 32.23586, 
    32.24437, 32.2527, 32.26085, 32.26881, 32.27659, 32.28419, 32.2916, 
    32.29884, 32.30589, 32.31276, 32.31944, 32.32594, 32.33226, 32.3384, 
    32.34436, 32.35012, 32.35571, 32.36112, 32.36634, 32.37138, 32.37623, 
    32.38091, 32.38539, 32.3897, 32.39382, 32.39775, 32.40151, 32.40508, 
    32.40847, 32.41167, 32.41469, 32.41753, 32.42018, 32.42265, 32.42493, 
    32.42703, 32.42895, 32.43068, 32.43223, 32.43359, 32.43478, 32.43577, 
    32.43658, 32.43721, 32.43766, 32.43792, 32.438, 32.43789, 32.4376, 
    32.43713, 32.43647, 32.43563, 32.4346, 32.43339, 32.432, 32.43042, 
    32.42866, 32.42671, 32.42458, 32.42227, 32.41977, 32.41709, 32.41423, 
    32.41117, 32.40794, 32.40453, 32.40093, 32.39714, 32.39318, 32.38903, 
    32.38469, 32.38018, 32.37548, 32.37059, 32.36552, 32.36028, 32.35484, 
    32.34922, 32.34343, 32.33744, 32.33128, 32.32493, 32.3184, 32.31168, 
    32.30478, 32.2977, 32.29044, 32.283, 32.27537, 32.26756, 32.25957, 
    32.25139, 32.24304, 32.2345, 32.22578, 32.21688, 32.20779, 32.19852, 
    32.18908, 32.17945, 32.16964, 32.15965, 32.14947, 32.13912, 32.12858, 
    32.11787, 32.10697, 32.09589, 32.08463, 32.07319, 32.06157, 32.04977, 
    32.0378, 32.02563, 32.01329, 32.00077, 31.98808, 31.97519, 31.96214, 
    31.9489, 31.93548, 31.92188, 31.90811, 31.89416, 31.88002, 31.86571, 
    31.85122, 31.83655, 31.8217, 31.80668, 31.79148, 31.7761, 31.76054, 
    31.7448, 31.72889, 31.7128, 31.69653, 31.68009, 31.66347, 31.64667, 
    31.6297, 31.61255, 31.59522, 31.57772, 31.56004, 31.54219, 31.52416, 
    31.50596, 31.48758, 31.46902, 31.4503, 31.43139, 31.41232, 31.39306, 
    31.37364, 31.35404, 31.33426, 31.31432, 31.2942, 31.2739, 31.25344, 
    31.2328, 31.21198, 31.191, 31.16984, 31.14851, 31.12701, 31.10534, 
    31.0835, 31.06148, 31.0393, 31.01694, 30.99441, 30.97171, 30.94884, 
    30.92581, 30.9026, 30.87922, 30.85567, 30.83195, 30.80807, 30.78401, 
    30.75979, 30.7354, 30.71084, 30.68611, 30.66122, 30.63615, 30.61092, 
    30.58553, 30.55996, 30.53423, 30.50833, 30.48227, 30.45604, 30.42964, 
    30.40308, 30.37636, 30.34946, 30.32241, 30.29519, 30.2678, 30.24025, 
    30.21254, 30.18466, 30.15662, 30.12842, 30.10005, 30.07152, 30.04283, 
    30.01397, 29.98495, 29.95578, 29.92644, 29.89694, 29.86727, 29.83745, 
    29.80747,
  26.46019, 26.50399, 26.54765, 26.59118, 26.63457, 26.67782, 26.72094, 
    26.76392, 26.80677, 26.84947, 26.89204, 26.93447, 26.97677, 27.01892, 
    27.06094, 27.10281, 27.14455, 27.18615, 27.22761, 27.26892, 27.3101, 
    27.35114, 27.39203, 27.43279, 27.4734, 27.51387, 27.5542, 27.59438, 
    27.63442, 27.67432, 27.71408, 27.75369, 27.79316, 27.83249, 27.87167, 
    27.9107, 27.94959, 27.98834, 28.02694, 28.06539, 28.10369, 28.14186, 
    28.17987, 28.21774, 28.25546, 28.29303, 28.33045, 28.36773, 28.40486, 
    28.44183, 28.47866, 28.51534, 28.55187, 28.58826, 28.62449, 28.66057, 
    28.6965, 28.73228, 28.7679, 28.80338, 28.83871, 28.87388, 28.9089, 
    28.94377, 28.97848, 29.01305, 29.04745, 29.08171, 29.11581, 29.14976, 
    29.18355, 29.21719, 29.25067, 29.284, 29.31717, 29.35019, 29.38305, 
    29.41575, 29.4483, 29.48069, 29.51293, 29.54501, 29.57693, 29.60869, 
    29.64029, 29.67174, 29.70302, 29.73415, 29.76512, 29.79593, 29.82658, 
    29.85707, 29.8874, 29.91757, 29.94758, 29.97742, 30.00711, 30.03664, 
    30.066, 30.0952, 30.12424, 30.15312, 30.18184, 30.21039, 30.23878, 
    30.26701, 30.29507, 30.32297, 30.3507, 30.37827, 30.40568, 30.43292, 
    30.46, 30.48691, 30.51366, 30.54024, 30.56665, 30.5929, 30.61898, 
    30.6449, 30.67065, 30.69623, 30.72165, 30.74689, 30.77198, 30.79689, 
    30.82163, 30.84621, 30.87062, 30.89486, 30.91892, 30.94283, 30.96656, 
    30.99012, 31.01351, 31.03673, 31.05979, 31.08267, 31.10538, 31.12792, 
    31.15029, 31.17249, 31.19451, 31.21637, 31.23805, 31.25957, 31.2809, 
    31.30207, 31.32306, 31.34389, 31.36454, 31.38501, 31.40531, 31.42544, 
    31.4454, 31.46518, 31.48479, 31.50422, 31.52348, 31.54256, 31.56147, 
    31.58021, 31.59877, 31.61715, 31.63536, 31.65339, 31.67125, 31.68893, 
    31.70644, 31.72377, 31.74092, 31.7579, 31.7747, 31.79132, 31.80776, 
    31.82403, 31.84012, 31.85604, 31.87177, 31.88733, 31.90271, 31.91791, 
    31.93294, 31.94778, 31.96245, 31.97694, 31.99125, 32.00538, 32.01933, 
    32.0331, 32.0467, 32.06011, 32.07334, 32.0864, 32.09927, 32.11197, 
    32.12448, 32.13681, 32.14897, 32.16094, 32.17273, 32.18435, 32.19578, 
    32.20703, 32.2181, 32.22898, 32.23969, 32.25022, 32.26056, 32.27073, 
    32.28071, 32.29051, 32.30013, 32.30956, 32.31882, 32.32789, 32.33678, 
    32.34549, 32.35401, 32.36235, 32.37052, 32.37849, 32.38629, 32.3939, 
    32.40133, 32.40858, 32.41564, 32.42252, 32.42922, 32.43574, 32.44207, 
    32.44822, 32.45418, 32.45996, 32.46556, 32.47097, 32.47621, 32.48125, 
    32.48612, 32.4908, 32.4953, 32.49961, 32.50373, 32.50768, 32.51144, 
    32.51502, 32.51841, 32.52162, 32.52465, 32.52749, 32.53014, 32.53262, 
    32.5349, 32.53701, 32.53893, 32.54067, 32.54222, 32.54359, 32.54477, 
    32.54577, 32.54659, 32.54721, 32.54766, 32.54792, 32.548, 32.54789, 
    32.5476, 32.54713, 32.54647, 32.54562, 32.54459, 32.54338, 32.54198, 
    32.54041, 32.53864, 32.53669, 32.53456, 32.53224, 32.52974, 32.52705, 
    32.52418, 32.52113, 32.51789, 32.51447, 32.51086, 32.50707, 32.50309, 
    32.49894, 32.49459, 32.49007, 32.48536, 32.48047, 32.47539, 32.47013, 
    32.46469, 32.45906, 32.45325, 32.44725, 32.44108, 32.43472, 32.42817, 
    32.42145, 32.41454, 32.40744, 32.40017, 32.39271, 32.38507, 32.37724, 
    32.36924, 32.36105, 32.35268, 32.34412, 32.33538, 32.32647, 32.31736, 
    32.30808, 32.29862, 32.28897, 32.27914, 32.26913, 32.25894, 32.24857, 
    32.23801, 32.22728, 32.21636, 32.20526, 32.19398, 32.18252, 32.17088, 
    32.15906, 32.14706, 32.13488, 32.12251, 32.10997, 32.09724, 32.08434, 
    32.07126, 32.058, 32.04456, 32.03093, 32.01714, 32.00315, 31.98899, 
    31.97466, 31.96014, 31.94545, 31.93057, 31.91552, 31.90029, 31.88488, 
    31.8693, 31.85353, 31.83759, 31.82147, 31.80517, 31.7887, 31.77205, 
    31.75522, 31.73822, 31.72104, 31.70368, 31.68615, 31.66844, 31.65055, 
    31.63249, 31.61426, 31.59584, 31.57726, 31.55849, 31.53956, 31.52044, 
    31.50116, 31.4817, 31.46206, 31.44225, 31.42227, 31.40211, 31.38178, 
    31.36128, 31.3406, 31.31976, 31.29873, 31.27754, 31.25617, 31.23463, 
    31.21292, 31.19104, 31.16899, 31.14676, 31.12436, 31.1018, 31.07906, 
    31.05615, 31.03307, 31.00982, 30.9864, 30.96281, 30.93906, 30.91513, 
    30.89103, 30.86677, 30.84233, 30.81773, 30.79296, 30.76802, 30.74291, 
    30.71764, 30.6922, 30.66659, 30.64081, 30.61487, 30.58876, 30.56248, 
    30.53605, 30.50944, 30.48266, 30.45573, 30.42862, 30.40136, 30.37392, 
    30.34633, 30.31857, 30.29064, 30.26255, 30.2343, 30.20588, 30.17731, 
    30.14856, 30.11966, 30.0906, 30.06137, 30.03198, 30.00243, 29.97271, 
    29.94284, 29.91281,
  26.56002, 26.60389, 26.64761, 26.6912, 26.73466, 26.77798, 26.82116, 
    26.86421, 26.90712, 26.94989, 26.99252, 27.03502, 27.07738, 27.1196, 
    27.16168, 27.20362, 27.24542, 27.28708, 27.3286, 27.36998, 27.41122, 
    27.45232, 27.49328, 27.5341, 27.57477, 27.61531, 27.6557, 27.69595, 
    27.73605, 27.77601, 27.81583, 27.8555, 27.89504, 27.93442, 27.97366, 
    28.01276, 28.05171, 28.09052, 28.12918, 28.16769, 28.20606, 28.24428, 
    28.28236, 28.32028, 28.35806, 28.39569, 28.43318, 28.47051, 28.5077, 
    28.54474, 28.58163, 28.61837, 28.65496, 28.6914, 28.72769, 28.76382, 
    28.79981, 28.83565, 28.87134, 28.90687, 28.94225, 28.97748, 29.01256, 
    29.04749, 29.08226, 29.11688, 29.15134, 29.18565, 29.21981, 29.25381, 
    29.28766, 29.32136, 29.35489, 29.38828, 29.4215, 29.45458, 29.48749, 
    29.52025, 29.55285, 29.5853, 29.61758, 29.64972, 29.68169, 29.7135, 
    29.74516, 29.77666, 29.808, 29.83918, 29.8702, 29.90106, 29.93176, 
    29.9623, 29.99268, 30.0229, 30.05296, 30.08286, 30.1126, 30.14217, 
    30.17159, 30.20084, 30.22993, 30.25886, 30.28762, 30.31622, 30.34466, 
    30.37294, 30.40105, 30.42899, 30.45678, 30.48439, 30.51185, 30.53914, 
    30.56626, 30.59322, 30.62001, 30.64664, 30.6731, 30.69939, 30.72552, 
    30.75148, 30.77728, 30.8029, 30.82836, 30.85365, 30.87878, 30.90373, 
    30.92852, 30.95314, 30.97759, 31.00187, 31.02599, 31.04993, 31.0737, 
    31.0973, 31.12074, 31.144, 31.16709, 31.19002, 31.21277, 31.23535, 
    31.25776, 31.27999, 31.30206, 31.32395, 31.34567, 31.36723, 31.3886, 
    31.40981, 31.43084, 31.4517, 31.47238, 31.4929, 31.51323, 31.5334, 
    31.55339, 31.57321, 31.59285, 31.61232, 31.63161, 31.65073, 31.66967, 
    31.68844, 31.70703, 31.72545, 31.74369, 31.76176, 31.77965, 31.79736, 
    31.8149, 31.83226, 31.84944, 31.86645, 31.88328, 31.89993, 31.91641, 
    31.9327, 31.94882, 31.96477, 31.98053, 31.99612, 32.01152, 32.02676, 
    32.04181, 32.05668, 32.07137, 32.08589, 32.10022, 32.11438, 32.12836, 
    32.14215, 32.15577, 32.16921, 32.18247, 32.19555, 32.20844, 32.22116, 
    32.2337, 32.24606, 32.25823, 32.27023, 32.28204, 32.29367, 32.30513, 
    32.3164, 32.32749, 32.3384, 32.34912, 32.35967, 32.37003, 32.38021, 
    32.39021, 32.40003, 32.40967, 32.41912, 32.42839, 32.43748, 32.44639, 
    32.45511, 32.46365, 32.47201, 32.48019, 32.48818, 32.49599, 32.50362, 
    32.51106, 32.51832, 32.5254, 32.53229, 32.539, 32.54553, 32.55187, 
    32.55803, 32.56401, 32.5698, 32.57541, 32.58083, 32.58607, 32.59113, 
    32.596, 32.60069, 32.6052, 32.60952, 32.61366, 32.61761, 32.62138, 
    32.62496, 32.62836, 32.63157, 32.6346, 32.63745, 32.64011, 32.64259, 
    32.64488, 32.64699, 32.64891, 32.65065, 32.65221, 32.65358, 32.65476, 
    32.65577, 32.65658, 32.65721, 32.65766, 32.65792, 32.658, 32.65789, 
    32.6576, 32.65712, 32.65646, 32.65562, 32.65459, 32.65337, 32.65197, 
    32.65039, 32.64862, 32.64667, 32.64453, 32.64221, 32.6397, 32.63701, 
    32.63414, 32.63108, 32.62783, 32.6244, 32.62079, 32.61699, 32.61301, 
    32.60884, 32.6045, 32.59996, 32.59525, 32.59034, 32.58526, 32.57999, 
    32.57453, 32.56889, 32.56307, 32.55707, 32.55088, 32.54451, 32.53795, 
    32.53121, 32.52429, 32.51719, 32.5099, 32.50242, 32.49477, 32.48693, 
    32.4789, 32.4707, 32.46231, 32.45374, 32.44499, 32.43606, 32.42694, 
    32.41764, 32.40816, 32.39849, 32.38865, 32.37862, 32.3684, 32.35801, 
    32.34744, 32.33668, 32.32574, 32.31463, 32.30333, 32.29185, 32.28019, 
    32.26834, 32.25632, 32.24411, 32.23173, 32.21916, 32.20641, 32.19349, 
    32.18038, 32.1671, 32.15363, 32.13998, 32.12616, 32.11215, 32.09797, 
    32.0836, 32.06906, 32.05434, 32.03944, 32.02436, 32.0091, 31.99366, 
    31.97805, 31.96226, 31.94629, 31.93014, 31.91381, 31.89731, 31.88063, 
    31.86377, 31.84674, 31.82952, 31.81214, 31.79457, 31.77683, 31.75891, 
    31.74082, 31.72255, 31.7041, 31.68548, 31.66669, 31.64772, 31.62857, 
    31.60925, 31.58975, 31.57008, 31.55024, 31.53022, 31.51003, 31.48966, 
    31.46912, 31.44841, 31.42752, 31.40646, 31.38523, 31.36383, 31.34225, 
    31.3205, 31.29858, 31.27649, 31.25422, 31.23179, 31.20918, 31.1864, 
    31.16345, 31.14033, 31.11704, 31.09358, 31.06995, 31.04615, 31.02218, 
    30.99804, 30.97374, 30.94926, 30.92461, 30.8998, 30.87481, 30.84966, 
    30.82435, 30.79886, 30.77321, 30.74739, 30.7214, 30.69525, 30.66892, 
    30.64244, 30.61578, 30.58897, 30.56198, 30.53483, 30.50752, 30.48004, 
    30.45239, 30.42458, 30.39661, 30.36847, 30.34017, 30.31171, 30.28308, 
    30.25429, 30.22534, 30.19622, 30.16695, 30.13751, 30.10791, 30.07814, 
    30.04822, 30.01813,
  26.65983, 26.70376, 26.74755, 26.79121, 26.83473, 26.87812, 26.92137, 
    26.96448, 27.00745, 27.05029, 27.09299, 27.13555, 27.17797, 27.22025, 
    27.2624, 27.3044, 27.34627, 27.38799, 27.42958, 27.47103, 27.51233, 
    27.55349, 27.59451, 27.6354, 27.67613, 27.71673, 27.75718, 27.79749, 
    27.83766, 27.87769, 27.91757, 27.9573, 27.99689, 28.03634, 28.07565, 
    28.11481, 28.15382, 28.19268, 28.23141, 28.26998, 28.30841, 28.34669, 
    28.38483, 28.42281, 28.46065, 28.49835, 28.53589, 28.57328, 28.61053, 
    28.64763, 28.68458, 28.72137, 28.75802, 28.79452, 28.83087, 28.86707, 
    28.90311, 28.93901, 28.97475, 29.01035, 29.04579, 29.08107, 29.11621, 
    29.15119, 29.18602, 29.22069, 29.25522, 29.28958, 29.3238, 29.35786, 
    29.39176, 29.42551, 29.4591, 29.49254, 29.52582, 29.55895, 29.59192, 
    29.62473, 29.65739, 29.68989, 29.72223, 29.75441, 29.78644, 29.81831, 
    29.85002, 29.88157, 29.91296, 29.94419, 29.97527, 30.00618, 30.03693, 
    30.06752, 30.09796, 30.12823, 30.15834, 30.18829, 30.21808, 30.2477, 
    30.27717, 30.30647, 30.33561, 30.36458, 30.3934, 30.42205, 30.45053, 
    30.47886, 30.50702, 30.53501, 30.56284, 30.59051, 30.61801, 30.64534, 
    30.67251, 30.69952, 30.72636, 30.75303, 30.77954, 30.80588, 30.83205, 
    30.85806, 30.8839, 30.90957, 30.93507, 30.96041, 30.98557, 31.01057, 
    31.0354, 31.06007, 31.08456, 31.10888, 31.13304, 31.15702, 31.18084, 
    31.20448, 31.22796, 31.25126, 31.27439, 31.29736, 31.32015, 31.34277, 
    31.36522, 31.38749, 31.4096, 31.43153, 31.45329, 31.47488, 31.49629, 
    31.51754, 31.53861, 31.5595, 31.58022, 31.60077, 31.62115, 31.64135, 
    31.66138, 31.68123, 31.7009, 31.72041, 31.73974, 31.75889, 31.77787, 
    31.79667, 31.81529, 31.83374, 31.85202, 31.87012, 31.88804, 31.90578, 
    31.92335, 31.94074, 31.95796, 31.975, 31.99186, 32.00854, 32.02505, 
    32.04137, 32.05752, 32.07349, 32.08929, 32.1049, 32.12034, 32.13559, 
    32.15067, 32.16557, 32.18029, 32.19484, 32.20919, 32.22338, 32.23738, 
    32.2512, 32.26485, 32.27831, 32.29159, 32.30469, 32.31762, 32.33035, 
    32.34291, 32.35529, 32.36749, 32.37951, 32.39135, 32.403, 32.41447, 
    32.42577, 32.43688, 32.44781, 32.45855, 32.46912, 32.4795, 32.4897, 
    32.49972, 32.50956, 32.51921, 32.52868, 32.53797, 32.54707, 32.556, 
    32.56474, 32.57329, 32.58167, 32.58986, 32.59787, 32.60569, 32.61333, 
    32.62079, 32.62806, 32.63515, 32.64206, 32.64878, 32.65532, 32.66167, 
    32.66785, 32.67383, 32.67963, 32.68525, 32.69069, 32.69594, 32.70101, 
    32.70589, 32.71059, 32.7151, 32.71943, 32.72357, 32.72753, 32.73131, 
    32.7349, 32.7383, 32.74152, 32.74456, 32.74741, 32.75008, 32.75256, 
    32.75486, 32.75697, 32.7589, 32.76064, 32.7622, 32.76357, 32.76476, 
    32.76576, 32.76658, 32.76721, 32.76766, 32.76792, 32.768, 32.76789, 
    32.7676, 32.76712, 32.76646, 32.76561, 32.76458, 32.76337, 32.76196, 
    32.76038, 32.75861, 32.75665, 32.75451, 32.75218, 32.74967, 32.74697, 
    32.74409, 32.74103, 32.73778, 32.73434, 32.73072, 32.72692, 32.72293, 
    32.71875, 32.7144, 32.70985, 32.70513, 32.70022, 32.69512, 32.68984, 
    32.68438, 32.67873, 32.6729, 32.66688, 32.66068, 32.6543, 32.64773, 
    32.64098, 32.63404, 32.62692, 32.61962, 32.61213, 32.60447, 32.59661, 
    32.58857, 32.58035, 32.57195, 32.56337, 32.5546, 32.54565, 32.53651, 
    32.52719, 32.51769, 32.50801, 32.49815, 32.4881, 32.47787, 32.46746, 
    32.45686, 32.44609, 32.43513, 32.42399, 32.41267, 32.40117, 32.38948, 
    32.37762, 32.36557, 32.35335, 32.34094, 32.32835, 32.31558, 32.30263, 
    32.2895, 32.27619, 32.2627, 32.24903, 32.23518, 32.22115, 32.20694, 
    32.19255, 32.17797, 32.16323, 32.1483, 32.13319, 32.11791, 32.10244, 
    32.0868, 32.07098, 32.05498, 32.0388, 32.02245, 32.00591, 31.9892, 
    31.97231, 31.95525, 31.93801, 31.92059, 31.90299, 31.88522, 31.86727, 
    31.84914, 31.83084, 31.81236, 31.7937, 31.77488, 31.75587, 31.73669, 
    31.71733, 31.69781, 31.6781, 31.65822, 31.63816, 31.61794, 31.59753, 
    31.57696, 31.55621, 31.53529, 31.51419, 31.49292, 31.47148, 31.44986, 
    31.42807, 31.40611, 31.38398, 31.36168, 31.3392, 31.31656, 31.29374, 
    31.27075, 31.24759, 31.22425, 31.20075, 31.17708, 31.15324, 31.12923, 
    31.10505, 31.0807, 31.05618, 31.03149, 31.00663, 30.9816, 30.95641, 
    30.93105, 30.90552, 30.87982, 30.85395, 30.82792, 30.80172, 30.77536, 
    30.74882, 30.72212, 30.69526, 30.66823, 30.64103, 30.61367, 30.58614, 
    30.55845, 30.53059, 30.50257, 30.47439, 30.44604, 30.41753, 30.38885, 
    30.36001, 30.33101, 30.30184, 30.27252, 30.24303, 30.21338, 30.18356, 
    30.15359, 30.12345,
  26.75962, 26.80362, 26.84748, 26.8912, 26.93479, 26.97824, 27.02155, 
    27.06473, 27.10777, 27.15067, 27.19343, 27.23606, 27.27855, 27.32089, 
    27.3631, 27.40517, 27.4471, 27.48889, 27.53054, 27.57205, 27.61342, 
    27.65464, 27.69573, 27.73667, 27.77748, 27.81813, 27.85865, 27.89902, 
    27.93925, 27.97934, 28.01929, 28.05908, 28.09874, 28.13825, 28.17761, 
    28.21683, 28.25591, 28.29484, 28.33362, 28.37226, 28.41074, 28.44909, 
    28.48728, 28.52533, 28.56323, 28.60098, 28.63859, 28.67604, 28.71335, 
    28.7505, 28.78751, 28.82437, 28.86108, 28.89763, 28.93404, 28.9703, 
    29.0064, 29.04236, 29.07816, 29.11381, 29.14931, 29.18465, 29.21984, 
    29.25488, 29.28977, 29.3245, 29.35908, 29.3935, 29.42777, 29.46189, 
    29.49585, 29.52965, 29.5633, 29.59679, 29.63013, 29.66331, 29.69634, 
    29.7292, 29.76192, 29.79447, 29.82686, 29.8591, 29.89118, 29.9231, 
    29.95486, 29.98647, 30.01791, 30.0492, 30.08032, 30.11129, 30.14209, 
    30.17274, 30.20322, 30.23355, 30.26371, 30.29371, 30.32354, 30.35322, 
    30.38273, 30.41209, 30.44127, 30.4703, 30.49916, 30.52786, 30.5564, 
    30.58477, 30.61298, 30.64102, 30.6689, 30.69661, 30.72416, 30.75154, 
    30.77876, 30.80581, 30.8327, 30.85942, 30.88597, 30.91235, 30.93857, 
    30.96462, 30.99051, 31.01622, 31.04177, 31.06715, 31.09236, 31.1174, 
    31.14228, 31.16698, 31.19152, 31.21589, 31.24008, 31.26411, 31.28797, 
    31.31165, 31.33517, 31.35851, 31.38169, 31.40469, 31.42752, 31.45018, 
    31.47267, 31.49499, 31.51713, 31.5391, 31.5609, 31.58253, 31.60398, 
    31.62526, 31.64637, 31.6673, 31.68806, 31.70865, 31.72906, 31.74929, 
    31.76936, 31.78925, 31.80896, 31.8285, 31.84786, 31.86704, 31.88606, 
    31.90489, 31.92355, 31.94204, 31.96034, 31.97847, 31.99643, 32.01421, 
    32.03181, 32.04923, 32.06647, 32.08354, 32.10043, 32.11715, 32.13368, 
    32.15004, 32.16622, 32.18222, 32.19804, 32.21368, 32.22915, 32.24443, 
    32.25954, 32.27446, 32.28921, 32.30378, 32.31816, 32.33237, 32.3464, 
    32.36025, 32.37392, 32.38741, 32.40071, 32.41384, 32.42678, 32.43955, 
    32.45213, 32.46453, 32.47675, 32.48879, 32.50065, 32.51233, 32.52382, 
    32.53513, 32.54626, 32.55721, 32.56798, 32.57856, 32.58897, 32.59919, 
    32.60922, 32.61908, 32.62875, 32.63824, 32.64754, 32.65666, 32.6656, 
    32.67436, 32.68293, 32.69132, 32.69953, 32.70755, 32.71539, 32.72304, 
    32.73051, 32.7378, 32.7449, 32.75182, 32.75856, 32.76511, 32.77148, 
    32.77766, 32.78366, 32.78947, 32.7951, 32.80054, 32.80581, 32.81088, 
    32.81577, 32.82048, 32.825, 32.82934, 32.83349, 32.83746, 32.84124, 
    32.84483, 32.84825, 32.85147, 32.85452, 32.85737, 32.86005, 32.86253, 
    32.86483, 32.86695, 32.86888, 32.87062, 32.87218, 32.87356, 32.87475, 
    32.87576, 32.87658, 32.87721, 32.87766, 32.87792, 32.878, 32.87789, 
    32.8776, 32.87712, 32.87646, 32.87561, 32.87458, 32.87336, 32.87195, 
    32.87036, 32.86859, 32.86663, 32.86448, 32.86215, 32.85963, 32.85693, 
    32.85405, 32.85098, 32.84772, 32.84428, 32.84065, 32.83684, 32.83284, 
    32.82866, 32.8243, 32.81975, 32.81501, 32.81009, 32.80499, 32.7997, 
    32.79422, 32.78856, 32.78272, 32.7767, 32.77048, 32.76409, 32.75751, 
    32.75074, 32.74379, 32.73666, 32.72934, 32.72184, 32.71416, 32.70629, 
    32.69824, 32.69001, 32.68159, 32.67299, 32.6642, 32.65523, 32.64608, 
    32.63675, 32.62723, 32.61753, 32.60765, 32.59758, 32.58733, 32.5769, 
    32.56629, 32.55549, 32.54452, 32.53336, 32.52201, 32.51049, 32.49879, 
    32.4869, 32.47483, 32.46258, 32.45015, 32.43754, 32.42475, 32.41177, 
    32.39862, 32.38528, 32.37177, 32.35807, 32.3442, 32.33014, 32.3159, 
    32.30149, 32.28689, 32.27211, 32.25716, 32.24202, 32.22671, 32.21122, 
    32.19555, 32.1797, 32.16367, 32.14746, 32.13108, 32.11451, 32.09777, 
    32.08086, 32.06376, 32.04649, 32.02903, 32.01141, 31.9936, 31.97562, 
    31.95746, 31.93912, 31.92061, 31.90192, 31.88306, 31.86402, 31.84481, 
    31.82542, 31.80585, 31.78611, 31.7662, 31.74611, 31.72584, 31.7054, 
    31.68479, 31.664, 31.64304, 31.62191, 31.6006, 31.57912, 31.55747, 
    31.53564, 31.51364, 31.49147, 31.46913, 31.44661, 31.42392, 31.40106, 
    31.37803, 31.35483, 31.33146, 31.30792, 31.2842, 31.26032, 31.23627, 
    31.21204, 31.18765, 31.16309, 31.13836, 31.11345, 31.08839, 31.06315, 
    31.03774, 31.01217, 30.98642, 30.96051, 30.93443, 30.90819, 30.88178, 
    30.8552, 30.82845, 30.80154, 30.77447, 30.74722, 30.71981, 30.69224, 
    30.6645, 30.63659, 30.60853, 30.58029, 30.5519, 30.52333, 30.49461, 
    30.46572, 30.43667, 30.40745, 30.37808, 30.34854, 30.31883, 30.28897, 
    30.25895, 30.22876,
  26.8594, 26.90346, 26.94738, 26.99117, 27.03483, 27.07834, 27.12172, 
    27.16496, 27.20807, 27.25103, 27.29386, 27.33655, 27.3791, 27.42152, 
    27.46379, 27.50592, 27.54792, 27.58977, 27.63148, 27.67306, 27.71449, 
    27.75578, 27.79693, 27.83794, 27.8788, 27.91952, 27.9601, 28.00054, 
    28.04083, 28.08098, 28.12099, 28.16085, 28.20057, 28.24014, 28.27956, 
    28.31885, 28.35798, 28.39697, 28.43582, 28.47451, 28.51306, 28.55147, 
    28.58972, 28.62783, 28.66579, 28.7036, 28.74127, 28.77878, 28.81615, 
    28.85336, 28.89043, 28.92735, 28.96412, 29.00073, 29.0372, 29.07351, 
    29.10968, 29.14569, 29.18155, 29.21725, 29.25281, 29.28821, 29.32346, 
    29.35856, 29.3935, 29.42829, 29.46293, 29.49741, 29.53173, 29.5659, 
    29.59992, 29.63378, 29.66749, 29.70103, 29.73443, 29.76766, 29.80074, 
    29.83366, 29.86643, 29.89904, 29.93149, 29.96378, 29.99591, 30.02789, 
    30.0597, 30.09136, 30.12285, 30.15419, 30.18537, 30.21639, 30.24724, 
    30.27794, 30.30848, 30.33885, 30.36906, 30.39911, 30.429, 30.45873, 
    30.48829, 30.51769, 30.54693, 30.57601, 30.60492, 30.63367, 30.66225, 
    30.69067, 30.71893, 30.74702, 30.77495, 30.80271, 30.8303, 30.85773, 
    30.885, 30.91209, 30.93903, 30.96579, 30.99239, 31.01882, 31.04509, 
    31.07118, 31.09711, 31.12287, 31.14846, 31.17389, 31.19914, 31.22423, 
    31.24915, 31.2739, 31.29848, 31.32288, 31.34712, 31.37119, 31.39509, 
    31.41882, 31.44238, 31.46576, 31.48898, 31.51202, 31.53489, 31.55759, 
    31.58012, 31.60248, 31.62466, 31.64667, 31.66851, 31.69017, 31.71166, 
    31.73298, 31.75413, 31.7751, 31.79589, 31.81651, 31.83696, 31.85723, 
    31.87733, 31.89726, 31.91701, 31.93658, 31.95597, 31.9752, 31.99424, 
    32.01311, 32.03181, 32.05032, 32.06866, 32.08683, 32.10481, 32.12262, 
    32.14025, 32.15771, 32.17498, 32.19209, 32.20901, 32.22575, 32.24231, 
    32.2587, 32.27491, 32.29094, 32.30679, 32.32246, 32.33795, 32.35326, 
    32.3684, 32.38335, 32.39812, 32.41272, 32.42714, 32.44137, 32.45542, 
    32.4693, 32.48299, 32.4965, 32.50983, 32.52298, 32.53595, 32.54874, 
    32.56134, 32.57377, 32.58601, 32.59807, 32.60995, 32.62165, 32.63317, 
    32.6445, 32.65565, 32.66662, 32.67741, 32.68801, 32.69843, 32.70867, 
    32.71872, 32.7286, 32.73829, 32.74779, 32.75711, 32.76625, 32.77521, 
    32.78398, 32.79257, 32.80098, 32.8092, 32.81723, 32.82508, 32.83276, 
    32.84024, 32.84754, 32.85466, 32.86159, 32.86834, 32.8749, 32.88128, 
    32.88747, 32.89348, 32.89931, 32.90495, 32.9104, 32.91567, 32.92076, 
    32.92566, 32.93037, 32.9349, 32.93925, 32.94341, 32.94738, 32.95117, 
    32.95477, 32.95819, 32.96143, 32.96447, 32.96733, 32.97001, 32.9725, 
    32.97481, 32.97693, 32.97886, 32.98061, 32.98217, 32.98355, 32.98475, 
    32.98575, 32.98657, 32.98721, 32.98766, 32.98792, 32.988, 32.98789, 
    32.9876, 32.98712, 32.98645, 32.9856, 32.98457, 32.98335, 32.98194, 
    32.98035, 32.97857, 32.9766, 32.97446, 32.97212, 32.9696, 32.9669, 
    32.964, 32.96093, 32.95766, 32.95422, 32.95058, 32.94677, 32.94276, 
    32.93857, 32.9342, 32.92964, 32.92489, 32.91996, 32.91485, 32.90955, 
    32.90407, 32.8984, 32.89254, 32.88651, 32.88028, 32.87387, 32.86728, 
    32.8605, 32.85354, 32.8464, 32.83907, 32.83155, 32.82386, 32.81598, 
    32.80791, 32.79966, 32.79122, 32.7826, 32.7738, 32.76482, 32.75565, 
    32.7463, 32.73676, 32.72705, 32.71714, 32.70706, 32.69679, 32.68634, 
    32.67571, 32.6649, 32.6539, 32.64272, 32.63136, 32.61981, 32.60809, 
    32.59618, 32.58409, 32.57182, 32.55936, 32.54673, 32.53391, 32.52091, 
    32.50773, 32.49437, 32.48083, 32.46711, 32.45321, 32.43913, 32.42487, 
    32.41042, 32.3958, 32.381, 32.36602, 32.35085, 32.33551, 32.31999, 
    32.30429, 32.28841, 32.27236, 32.25612, 32.2397, 32.22311, 32.20634, 
    32.18939, 32.17226, 32.15496, 32.13748, 32.11982, 32.10198, 32.08397, 
    32.06577, 32.04741, 32.02886, 32.01014, 31.99124, 31.97217, 31.95292, 
    31.93349, 31.91389, 31.89412, 31.87417, 31.85404, 31.83374, 31.81326, 
    31.79262, 31.77179, 31.75079, 31.72962, 31.70828, 31.68676, 31.66507, 
    31.6432, 31.62116, 31.59895, 31.57657, 31.55401, 31.53129, 31.50839, 
    31.48532, 31.46207, 31.43866, 31.41508, 31.39132, 31.3674, 31.3433, 
    31.31903, 31.2946, 31.26999, 31.24522, 31.22027, 31.19516, 31.16988, 
    31.14443, 31.11881, 31.09302, 31.06706, 31.04094, 31.01465, 30.98819, 
    30.96157, 30.93478, 30.90782, 30.8807, 30.8534, 30.82595, 30.79833, 
    30.77054, 30.74259, 30.71447, 30.68619, 30.65774, 30.62913, 30.60036, 
    30.57142, 30.54232, 30.51305, 30.48363, 30.45404, 30.42429, 30.39437, 
    30.36429, 30.33406,
  26.95915, 27.00328, 27.04727, 27.09113, 27.13484, 27.17843, 27.22187, 
    27.26518, 27.30835, 27.35138, 27.39427, 27.43703, 27.47964, 27.52212, 
    27.56446, 27.60666, 27.64872, 27.69063, 27.73241, 27.77405, 27.81554, 
    27.8569, 27.89811, 27.93918, 27.98011, 28.0209, 28.06154, 28.10204, 
    28.14239, 28.1826, 28.22267, 28.2626, 28.30238, 28.34201, 28.3815, 
    28.42084, 28.46004, 28.49909, 28.538, 28.57676, 28.61537, 28.65383, 
    28.69215, 28.73032, 28.76834, 28.80621, 28.84394, 28.88151, 28.91894, 
    28.95621, 28.99334, 29.03032, 29.06714, 29.10382, 29.14034, 29.17671, 
    29.21294, 29.24901, 29.28492, 29.32069, 29.3563, 29.39176, 29.42707, 
    29.46222, 29.49722, 29.53207, 29.56676, 29.6013, 29.63568, 29.66991, 
    29.70398, 29.7379, 29.77166, 29.80526, 29.83871, 29.872, 29.90514, 
    29.93811, 29.97093, 30.00359, 30.0361, 30.06844, 30.10063, 30.13266, 
    30.16453, 30.19624, 30.22779, 30.25918, 30.29041, 30.32148, 30.35238, 
    30.38313, 30.41372, 30.44415, 30.47441, 30.50451, 30.53445, 30.56423, 
    30.59384, 30.62329, 30.65258, 30.68171, 30.71067, 30.73947, 30.7681, 
    30.79657, 30.82487, 30.85301, 30.88099, 30.90879, 30.93644, 30.96391, 
    30.99122, 31.01837, 31.04535, 31.07216, 31.0988, 31.12528, 31.15159, 
    31.17773, 31.20371, 31.22951, 31.25515, 31.28062, 31.30592, 31.33105, 
    31.35601, 31.3808, 31.40542, 31.42987, 31.45416, 31.47827, 31.50221, 
    31.52598, 31.54958, 31.573, 31.59626, 31.61934, 31.64226, 31.665, 
    31.68756, 31.70996, 31.73218, 31.75423, 31.77611, 31.79781, 31.81934, 
    31.8407, 31.86188, 31.88289, 31.90372, 31.92438, 31.94486, 31.96517, 
    31.98531, 32.00526, 32.02505, 32.04465, 32.06409, 32.08334, 32.10242, 
    32.12133, 32.14005, 32.1586, 32.17698, 32.19518, 32.21319, 32.23103, 
    32.2487, 32.26619, 32.28349, 32.30062, 32.31757, 32.33435, 32.35094, 
    32.36736, 32.3836, 32.39965, 32.41553, 32.43124, 32.44675, 32.4621, 
    32.47726, 32.49224, 32.50704, 32.52166, 32.5361, 32.55036, 32.56444, 
    32.57834, 32.59206, 32.60559, 32.61895, 32.63212, 32.64511, 32.65792, 
    32.67056, 32.683, 32.69527, 32.70735, 32.71925, 32.73097, 32.74251, 
    32.75386, 32.76503, 32.77602, 32.78683, 32.79745, 32.80789, 32.81815, 
    32.82822, 32.83812, 32.84782, 32.85735, 32.86668, 32.87584, 32.88482, 
    32.8936, 32.90221, 32.91063, 32.91887, 32.92691, 32.93478, 32.94247, 
    32.94997, 32.95728, 32.96441, 32.97136, 32.97812, 32.98469, 32.99108, 
    32.99728, 33.00331, 33.00914, 33.01479, 33.02026, 33.02554, 33.03063, 
    33.03554, 33.04026, 33.0448, 33.04916, 33.05332, 33.0573, 33.0611, 
    33.06471, 33.06814, 33.07138, 33.07443, 33.0773, 33.07998, 33.08247, 
    33.08479, 33.08691, 33.08884, 33.0906, 33.09216, 33.09354, 33.09474, 
    33.09575, 33.09657, 33.09721, 33.09766, 33.09792, 33.098, 33.09789, 
    33.0976, 33.09712, 33.09645, 33.0956, 33.09456, 33.09334, 33.09193, 
    33.09033, 33.08855, 33.08659, 33.08443, 33.08209, 33.07957, 33.07685, 
    33.07396, 33.07088, 33.06761, 33.06415, 33.06051, 33.05669, 33.05268, 
    33.04848, 33.0441, 33.03953, 33.03477, 33.02984, 33.02472, 33.01941, 
    33.01391, 33.00823, 33.00237, 32.99632, 32.99008, 32.98366, 32.97706, 
    32.97027, 32.96329, 32.95613, 32.94879, 32.94127, 32.93355, 32.92566, 
    32.91757, 32.90931, 32.90086, 32.89222, 32.88341, 32.8744, 32.86522, 
    32.85585, 32.8463, 32.83656, 32.82664, 32.81654, 32.80626, 32.79578, 
    32.78513, 32.7743, 32.76328, 32.75208, 32.7407, 32.72913, 32.71738, 
    32.70545, 32.69334, 32.68105, 32.66857, 32.65591, 32.64307, 32.63005, 
    32.61685, 32.60346, 32.5899, 32.57615, 32.56223, 32.54811, 32.53383, 
    32.51936, 32.50471, 32.48988, 32.47487, 32.45968, 32.44431, 32.42876, 
    32.41304, 32.39713, 32.38104, 32.36478, 32.34833, 32.33171, 32.31491, 
    32.29792, 32.28077, 32.26343, 32.24591, 32.22823, 32.21035, 32.19231, 
    32.17408, 32.15568, 32.1371, 32.11835, 32.09942, 32.08031, 32.06103, 
    32.04156, 32.02193, 32.00212, 31.98213, 31.96197, 31.94163, 31.92112, 
    31.90044, 31.87957, 31.85854, 31.83733, 31.81595, 31.79439, 31.77266, 
    31.75076, 31.72868, 31.70643, 31.68401, 31.66141, 31.63864, 31.6157, 
    31.59259, 31.56931, 31.54585, 31.52223, 31.49843, 31.47446, 31.45033, 
    31.42602, 31.40154, 31.37689, 31.35207, 31.32708, 31.30193, 31.2766, 
    31.2511, 31.22544, 31.19961, 31.17361, 31.14744, 31.1211, 31.0946, 
    31.06793, 31.04109, 31.01409, 30.98692, 30.95958, 30.93208, 30.90441, 
    30.87657, 30.84857, 30.82041, 30.79208, 30.76358, 30.73492, 30.7061, 
    30.67711, 30.64796, 30.61864, 30.58917, 30.55953, 30.52972, 30.49976, 
    30.46963, 30.43934,
  27.05889, 27.10308, 27.14714, 27.19106, 27.23484, 27.27849, 27.322, 
    27.36537, 27.40861, 27.45171, 27.49467, 27.53749, 27.58017, 27.62271, 
    27.66511, 27.70737, 27.7495, 27.79148, 27.83332, 27.87502, 27.91658, 
    27.958, 27.99928, 28.04041, 28.0814, 28.12225, 28.16295, 28.20352, 
    28.24394, 28.28421, 28.32434, 28.36433, 28.40417, 28.44387, 28.48342, 
    28.52282, 28.56208, 28.60119, 28.64016, 28.67898, 28.71766, 28.75618, 
    28.79456, 28.83279, 28.87087, 28.9088, 28.94659, 28.98422, 29.02171, 
    29.05904, 29.09623, 29.13327, 29.17015, 29.20689, 29.24347, 29.2799, 
    29.31618, 29.35231, 29.38829, 29.42411, 29.45978, 29.4953, 29.53066, 
    29.56588, 29.60093, 29.63584, 29.67058, 29.70518, 29.73962, 29.7739, 
    29.80803, 29.842, 29.87582, 29.90948, 29.94298, 29.97633, 30.00952, 
    30.04255, 30.07542, 30.10814, 30.1407, 30.1731, 30.20534, 30.23742, 
    30.26934, 30.3011, 30.33271, 30.36415, 30.39543, 30.42655, 30.45751, 
    30.48831, 30.51895, 30.54943, 30.57974, 30.6099, 30.63989, 30.66972, 
    30.69938, 30.72888, 30.75822, 30.7874, 30.81641, 30.84525, 30.87394, 
    30.90245, 30.93081, 30.95899, 30.98701, 31.01487, 31.04256, 31.07009, 
    31.09744, 31.12464, 31.15166, 31.17852, 31.20521, 31.23173, 31.25809, 
    31.28428, 31.3103, 31.33615, 31.36183, 31.38734, 31.41268, 31.43786, 
    31.46286, 31.4877, 31.51236, 31.53686, 31.56118, 31.58533, 31.60932, 
    31.63313, 31.65677, 31.68024, 31.70354, 31.72666, 31.74961, 31.77239, 
    31.795, 31.81744, 31.8397, 31.86179, 31.8837, 31.90544, 31.92701, 
    31.94841, 31.96963, 31.99067, 32.01154, 32.03224, 32.05276, 32.0731, 
    32.09327, 32.11327, 32.13309, 32.15273, 32.1722, 32.19149, 32.2106, 
    32.22954, 32.2483, 32.26688, 32.28529, 32.30352, 32.32157, 32.33944, 
    32.35714, 32.37466, 32.392, 32.40916, 32.42614, 32.44294, 32.45957, 
    32.47602, 32.49228, 32.50837, 32.52428, 32.54, 32.55555, 32.57092, 
    32.58611, 32.60112, 32.61595, 32.6306, 32.64506, 32.65935, 32.67345, 
    32.68738, 32.70112, 32.71468, 32.72806, 32.74126, 32.75428, 32.76711, 
    32.77976, 32.79223, 32.80452, 32.81663, 32.82855, 32.84029, 32.85185, 
    32.86322, 32.87442, 32.88543, 32.89625, 32.90689, 32.91735, 32.92763, 
    32.93773, 32.94763, 32.95736, 32.9669, 32.97626, 32.98543, 32.99442, 
    33.00322, 33.01184, 33.02028, 33.02853, 33.0366, 33.04448, 33.05218, 
    33.05969, 33.06702, 33.07416, 33.08112, 33.08789, 33.09448, 33.10088, 
    33.1071, 33.11313, 33.11898, 33.12464, 33.13011, 33.1354, 33.14051, 
    33.14542, 33.15016, 33.15471, 33.15907, 33.16324, 33.16723, 33.17103, 
    33.17465, 33.17808, 33.18132, 33.18438, 33.18726, 33.18995, 33.19244, 
    33.19476, 33.19689, 33.19883, 33.20058, 33.20215, 33.20354, 33.20473, 
    33.20574, 33.20657, 33.20721, 33.20766, 33.20792, 33.208, 33.20789, 
    33.2076, 33.20712, 33.20645, 33.2056, 33.20456, 33.20333, 33.20192, 
    33.20032, 33.19854, 33.19656, 33.1944, 33.19206, 33.18953, 33.18682, 
    33.18391, 33.18082, 33.17755, 33.17409, 33.17044, 33.16661, 33.16259, 
    33.15839, 33.154, 33.14942, 33.14466, 33.13971, 33.13458, 33.12926, 
    33.12375, 33.11806, 33.11219, 33.10613, 33.09988, 33.09345, 33.08683, 
    33.08003, 33.07304, 33.06587, 33.05851, 33.05097, 33.04324, 33.03534, 
    33.02724, 33.01896, 33.01049, 33.00184, 32.99301, 32.98399, 32.97479, 
    32.9654, 32.95583, 32.94608, 32.93614, 32.92602, 32.91571, 32.90522, 
    32.89455, 32.8837, 32.87266, 32.86144, 32.85003, 32.83845, 32.82668, 
    32.81472, 32.80259, 32.79027, 32.77777, 32.76509, 32.75223, 32.73919, 
    32.72596, 32.71255, 32.69896, 32.68519, 32.67123, 32.6571, 32.64279, 
    32.62829, 32.61361, 32.59876, 32.58372, 32.5685, 32.55311, 32.53753, 
    32.52177, 32.50584, 32.48972, 32.47343, 32.45695, 32.4403, 32.42347, 
    32.40646, 32.38927, 32.3719, 32.35435, 32.33663, 32.31873, 32.30065, 
    32.28239, 32.26395, 32.24534, 32.22655, 32.20759, 32.18845, 32.16913, 
    32.14964, 32.12996, 32.11012, 32.0901, 32.0699, 32.04952, 32.02898, 
    32.00825, 31.98735, 31.96628, 31.94503, 31.92361, 31.90202, 31.88025, 
    31.8583, 31.83619, 31.8139, 31.79144, 31.7688, 31.74599, 31.72301, 
    31.69986, 31.67654, 31.65304, 31.62938, 31.60554, 31.58153, 31.55735, 
    31.53299, 31.50847, 31.48378, 31.45892, 31.43389, 31.40869, 31.38331, 
    31.35777, 31.33207, 31.30619, 31.28014, 31.25393, 31.22755, 31.201, 
    31.17428, 31.1474, 31.12035, 31.09313, 31.06574, 31.03819, 31.01048, 
    30.98259, 30.95455, 30.92633, 30.89795, 30.86941, 30.8407, 30.81183, 
    30.78279, 30.75359, 30.72423, 30.6947, 30.66501, 30.63515, 30.60514, 
    30.57496, 30.54462,
  27.15861, 27.20286, 27.24699, 27.29097, 27.33482, 27.37854, 27.42211, 
    27.46555, 27.50885, 27.55201, 27.59504, 27.63792, 27.68067, 27.72328, 
    27.76575, 27.80807, 27.85026, 27.89231, 27.93421, 27.97598, 28.0176, 
    28.05908, 28.10042, 28.14162, 28.18267, 28.22359, 28.26436, 28.30498, 
    28.34546, 28.3858, 28.42599, 28.46604, 28.50595, 28.54571, 28.58532, 
    28.62479, 28.66411, 28.70328, 28.74231, 28.78119, 28.81993, 28.85851, 
    28.89695, 28.93524, 28.97338, 29.01138, 29.04922, 29.08692, 29.12446, 
    29.16186, 29.19911, 29.2362, 29.27315, 29.30994, 29.34658, 29.38307, 
    29.41941, 29.4556, 29.49164, 29.52752, 29.56325, 29.59882, 29.63424, 
    29.66951, 29.70463, 29.73959, 29.77439, 29.80904, 29.84354, 29.87788, 
    29.91207, 29.94609, 29.97997, 30.01368, 30.04724, 30.08064, 30.11389, 
    30.14697, 30.1799, 30.21267, 30.24528, 30.27774, 30.31003, 30.34217, 
    30.37414, 30.40596, 30.43761, 30.46911, 30.50045, 30.53162, 30.56263, 
    30.59348, 30.62418, 30.6547, 30.68507, 30.71527, 30.74532, 30.77519, 
    30.80491, 30.83446, 30.86385, 30.89307, 30.92213, 30.95103, 30.97976, 
    31.00833, 31.03673, 31.06497, 31.09304, 31.12094, 31.14868, 31.17625, 
    31.20366, 31.23089, 31.25797, 31.28487, 31.31161, 31.33818, 31.36458, 
    31.39081, 31.41687, 31.44277, 31.4685, 31.49405, 31.51944, 31.54466, 
    31.56971, 31.59459, 31.6193, 31.64383, 31.6682, 31.6924, 31.71642, 
    31.74027, 31.76396, 31.78747, 31.8108, 31.83397, 31.85696, 31.87979, 
    31.90243, 31.92491, 31.94721, 31.96934, 31.99129, 32.01307, 32.03468, 
    32.05611, 32.07737, 32.09845, 32.11936, 32.14009, 32.16065, 32.18103, 
    32.20124, 32.22127, 32.24112, 32.2608, 32.2803, 32.29963, 32.31878, 
    32.33775, 32.35654, 32.37516, 32.3936, 32.41186, 32.42994, 32.44785, 
    32.46558, 32.48313, 32.5005, 32.51769, 32.5347, 32.55154, 32.56819, 
    32.58467, 32.60096, 32.61708, 32.63302, 32.64878, 32.66435, 32.67975, 
    32.69497, 32.71, 32.72486, 32.73953, 32.75402, 32.76833, 32.78247, 
    32.79642, 32.81018, 32.82377, 32.83717, 32.8504, 32.86344, 32.87629, 
    32.88897, 32.90146, 32.91378, 32.9259, 32.93785, 32.94961, 32.96119, 
    32.97259, 32.9838, 32.99483, 33.00568, 33.01634, 33.02682, 33.03711, 
    33.04722, 33.05715, 33.06689, 33.07645, 33.08583, 33.09502, 33.10402, 
    33.11284, 33.12148, 33.12993, 33.1382, 33.14628, 33.15417, 33.16189, 
    33.16941, 33.17675, 33.18391, 33.19088, 33.19767, 33.20427, 33.21068, 
    33.21691, 33.22295, 33.22881, 33.23448, 33.23997, 33.24527, 33.25038, 
    33.25531, 33.26005, 33.2646, 33.26897, 33.27316, 33.27715, 33.28096, 
    33.28459, 33.28802, 33.29128, 33.29434, 33.29722, 33.29991, 33.30242, 
    33.30473, 33.30687, 33.30881, 33.31057, 33.31214, 33.31353, 33.31473, 
    33.31574, 33.31657, 33.3172, 33.31766, 33.31792, 33.318, 33.31789, 
    33.3176, 33.31712, 33.31645, 33.31559, 33.31455, 33.31332, 33.3119, 
    33.31031, 33.30852, 33.30654, 33.30438, 33.30203, 33.2995, 33.29678, 
    33.29387, 33.29078, 33.28749, 33.28403, 33.28037, 33.27654, 33.27251, 
    33.2683, 33.2639, 33.25931, 33.25454, 33.24958, 33.24444, 33.23911, 
    33.2336, 33.2279, 33.22201, 33.21594, 33.20968, 33.20324, 33.19661, 
    33.18979, 33.18279, 33.17561, 33.16824, 33.16068, 33.15294, 33.14501, 
    33.1369, 33.1286, 33.12012, 33.11146, 33.10261, 33.09357, 33.08435, 
    33.07495, 33.06536, 33.05559, 33.04564, 33.0355, 33.02517, 33.01466, 
    33.00397, 32.9931, 32.98204, 32.97079, 32.95937, 32.94776, 32.93597, 
    32.924, 32.91184, 32.8995, 32.88698, 32.87427, 32.86139, 32.84832, 
    32.83506, 32.82163, 32.80802, 32.79422, 32.78024, 32.76608, 32.75174, 
    32.73722, 32.72252, 32.70763, 32.69257, 32.67733, 32.6619, 32.64629, 
    32.63051, 32.61454, 32.5984, 32.58207, 32.56557, 32.54889, 32.53202, 
    32.51498, 32.49776, 32.48036, 32.46278, 32.44503, 32.42709, 32.40898, 
    32.39069, 32.37222, 32.35358, 32.33475, 32.31576, 32.29658, 32.27723, 
    32.2577, 32.23799, 32.21811, 32.19805, 32.17782, 32.15741, 32.13682, 
    32.11606, 32.09513, 32.07402, 32.05273, 32.03127, 32.00964, 31.98783, 
    31.96585, 31.94369, 31.92136, 31.89886, 31.87619, 31.85334, 31.83032, 
    31.80713, 31.78376, 31.76022, 31.73651, 31.71263, 31.68858, 31.66436, 
    31.63996, 31.6154, 31.59066, 31.56576, 31.54068, 31.51544, 31.49002, 
    31.46444, 31.43868, 31.41276, 31.38667, 31.36041, 31.33398, 31.30739, 
    31.28063, 31.25369, 31.2266, 31.19933, 31.1719, 31.1443, 31.11654, 
    31.08861, 31.06051, 31.03225, 31.00382, 30.97523, 30.94647, 30.91755, 
    30.88846, 30.85921, 30.8298, 30.80022, 30.77048, 30.74057, 30.71051, 
    30.68028, 30.64989,
  27.2583, 27.30263, 27.34682, 27.39087, 27.43479, 27.47856, 27.52221, 
    27.56571, 27.60908, 27.6523, 27.69539, 27.73834, 27.78115, 27.82383, 
    27.86636, 27.90875, 27.951, 27.99311, 28.03509, 28.07691, 28.1186, 
    28.16015, 28.20155, 28.24281, 28.28393, 28.32491, 28.36574, 28.40643, 
    28.44697, 28.48737, 28.52763, 28.56774, 28.60771, 28.64753, 28.6872, 
    28.72673, 28.76612, 28.80536, 28.84444, 28.88339, 28.92218, 28.96083, 
    28.99933, 29.03768, 29.07589, 29.11394, 29.15185, 29.1896, 29.22721, 
    29.26466, 29.30197, 29.33912, 29.37613, 29.41298, 29.44968, 29.48623, 
    29.52263, 29.55888, 29.59497, 29.63091, 29.6667, 29.70233, 29.73781, 
    29.77314, 29.80831, 29.84333, 29.87819, 29.9129, 29.94745, 29.98185, 
    30.01609, 30.05017, 30.0841, 30.11787, 30.15149, 30.18494, 30.21824, 
    30.25138, 30.28437, 30.31719, 30.34986, 30.38237, 30.41471, 30.44691, 
    30.47893, 30.5108, 30.54251, 30.57406, 30.60545, 30.63667, 30.66774, 
    30.69864, 30.72939, 30.75997, 30.79038, 30.82064, 30.85073, 30.88066, 
    30.91043, 30.94003, 30.96947, 30.99874, 31.02785, 31.0568, 31.08558, 
    31.11419, 31.14264, 31.17093, 31.19905, 31.227, 31.25479, 31.28241, 
    31.30986, 31.33714, 31.36426, 31.39121, 31.418, 31.44461, 31.47106, 
    31.49734, 31.52345, 31.54939, 31.57516, 31.60076, 31.62619, 31.65145, 
    31.67655, 31.70147, 31.72622, 31.7508, 31.77521, 31.79945, 31.82352, 
    31.84741, 31.87114, 31.89469, 31.91807, 31.94127, 31.96431, 31.98717, 
    32.00986, 32.03237, 32.05471, 32.07688, 32.09887, 32.12069, 32.14234, 
    32.16381, 32.1851, 32.20622, 32.22717, 32.24794, 32.26853, 32.28895, 
    32.30919, 32.32926, 32.34915, 32.36886, 32.3884, 32.40776, 32.42694, 
    32.44595, 32.46478, 32.48343, 32.5019, 32.5202, 32.53831, 32.55625, 
    32.57401, 32.59159, 32.60899, 32.62622, 32.64326, 32.66013, 32.67681, 
    32.69332, 32.70964, 32.72579, 32.74176, 32.75754, 32.77315, 32.78857, 
    32.80381, 32.81888, 32.83376, 32.84846, 32.86298, 32.87732, 32.89148, 
    32.90545, 32.91924, 32.93285, 32.94629, 32.95953, 32.9726, 32.98548, 
    32.99818, 33.01069, 33.02303, 33.03518, 33.04714, 33.05893, 33.07053, 
    33.08195, 33.09318, 33.10423, 33.11509, 33.12578, 33.13628, 33.14659, 
    33.15672, 33.16666, 33.17643, 33.186, 33.19539, 33.2046, 33.21362, 
    33.22246, 33.23111, 33.23958, 33.24786, 33.25596, 33.26387, 33.2716, 
    33.27914, 33.28649, 33.29366, 33.30064, 33.30744, 33.31406, 33.32048, 
    33.32672, 33.33278, 33.33865, 33.34433, 33.34982, 33.35513, 33.36025, 
    33.36519, 33.36994, 33.3745, 33.37888, 33.38307, 33.38708, 33.3909, 
    33.39452, 33.39797, 33.40123, 33.4043, 33.40718, 33.40988, 33.41239, 
    33.41471, 33.41685, 33.4188, 33.42056, 33.42213, 33.42352, 33.42472, 
    33.42574, 33.42656, 33.4272, 33.42765, 33.42792, 33.428, 33.42789, 
    33.4276, 33.42711, 33.42645, 33.42559, 33.42455, 33.42331, 33.42189, 
    33.42029, 33.4185, 33.41652, 33.41436, 33.412, 33.40946, 33.40674, 
    33.40382, 33.40072, 33.39744, 33.39396, 33.3903, 33.38646, 33.38242, 
    33.3782, 33.37379, 33.3692, 33.36442, 33.35946, 33.35431, 33.34896, 
    33.34344, 33.33773, 33.33183, 33.32575, 33.31948, 33.31302, 33.30638, 
    33.29955, 33.29254, 33.28534, 33.27796, 33.27039, 33.26263, 33.25469, 
    33.24656, 33.23825, 33.22976, 33.22107, 33.21221, 33.20316, 33.19392, 
    33.1845, 33.17489, 33.1651, 33.15513, 33.14497, 33.13463, 33.1241, 
    33.11339, 33.10249, 33.09142, 33.08015, 33.06871, 33.05708, 33.04526, 
    33.03327, 33.02109, 33.00872, 32.99618, 32.98345, 32.97054, 32.95745, 
    32.94417, 32.93071, 32.91708, 32.90325, 32.88925, 32.87506, 32.86069, 
    32.84615, 32.83142, 32.81651, 32.80141, 32.78614, 32.77069, 32.75505, 
    32.73924, 32.72325, 32.70707, 32.69072, 32.67418, 32.65747, 32.64058, 
    32.6235, 32.60625, 32.58882, 32.57121, 32.55342, 32.53546, 32.51731, 
    32.49899, 32.48049, 32.46181, 32.44296, 32.42392, 32.40471, 32.38532, 
    32.36576, 32.34602, 32.3261, 32.306, 32.28573, 32.26529, 32.24466, 
    32.22387, 32.20289, 32.18175, 32.16042, 32.13892, 32.11725, 32.09541, 
    32.07339, 32.05119, 32.02882, 32.00628, 31.98356, 31.96068, 31.93761, 
    31.91438, 31.89097, 31.8674, 31.84365, 31.81972, 31.79563, 31.77136, 
    31.74693, 31.72232, 31.69754, 31.67259, 31.64747, 31.62218, 31.59672, 
    31.57109, 31.5453, 31.51933, 31.49319, 31.46689, 31.44041, 31.41377, 
    31.38696, 31.35999, 31.33284, 31.30553, 31.27805, 31.2504, 31.22259, 
    31.19461, 31.16647, 31.13815, 31.10968, 31.08104, 31.05223, 31.02326, 
    30.99412, 30.96482, 30.93536, 30.90573, 30.87594, 30.84598, 30.81586, 
    30.78559, 30.75514,
  27.35798, 27.40237, 27.44663, 27.49075, 27.53473, 27.57857, 27.62228, 
    27.66585, 27.70928, 27.75257, 27.79573, 27.83875, 27.88162, 27.92436, 
    27.96696, 28.00941, 28.05173, 28.09391, 28.13594, 28.17783, 28.21959, 
    28.2612, 28.30266, 28.34399, 28.38517, 28.42621, 28.46711, 28.50786, 
    28.54847, 28.58893, 28.62925, 28.66942, 28.70945, 28.74934, 28.78907, 
    28.82867, 28.86811, 28.90741, 28.94656, 28.98557, 29.02442, 29.06313, 
    29.10169, 29.14011, 29.17837, 29.21649, 29.25445, 29.29227, 29.32993, 
    29.36745, 29.40482, 29.44203, 29.4791, 29.51601, 29.55277, 29.58938, 
    29.62584, 29.66214, 29.69829, 29.73429, 29.77014, 29.80583, 29.84137, 
    29.87675, 29.91198, 29.94705, 29.98197, 30.01674, 30.05135, 30.0858, 
    30.1201, 30.15424, 30.18822, 30.22205, 30.25572, 30.28923, 30.32259, 
    30.35578, 30.38882, 30.4217, 30.45442, 30.48698, 30.51939, 30.55163, 
    30.58371, 30.61564, 30.6474, 30.679, 30.71044, 30.74172, 30.77284, 
    30.80379, 30.83459, 30.86522, 30.89569, 30.926, 30.95614, 30.98612, 
    31.01594, 31.04559, 31.07508, 31.1044, 31.13356, 31.16256, 31.19139, 
    31.22005, 31.24855, 31.27688, 31.30505, 31.33305, 31.36089, 31.38855, 
    31.41605, 31.44339, 31.47055, 31.49755, 31.52438, 31.55104, 31.57753, 
    31.60386, 31.63001, 31.656, 31.68181, 31.70746, 31.73294, 31.75824, 
    31.78338, 31.80835, 31.83314, 31.85777, 31.88222, 31.9065, 31.93061, 
    31.95455, 31.97831, 32.0019, 32.02533, 32.04857, 32.07165, 32.09455, 
    32.11728, 32.13983, 32.16221, 32.18442, 32.20645, 32.22831, 32.24999, 
    32.2715, 32.29284, 32.31399, 32.33497, 32.35578, 32.37641, 32.39687, 
    32.41714, 32.43725, 32.45717, 32.47692, 32.49649, 32.51589, 32.53511, 
    32.55415, 32.57301, 32.59169, 32.6102, 32.62853, 32.64668, 32.66465, 
    32.68244, 32.70005, 32.71749, 32.73474, 32.75182, 32.76871, 32.78543, 
    32.80196, 32.81832, 32.8345, 32.85049, 32.8663, 32.88194, 32.89739, 
    32.91266, 32.92775, 32.94266, 32.95739, 32.97194, 32.9863, 33.00048, 
    33.01448, 33.0283, 33.04194, 33.05539, 33.06866, 33.08175, 33.09466, 
    33.10738, 33.11992, 33.13227, 33.14445, 33.15644, 33.16824, 33.17986, 
    33.1913, 33.20256, 33.21363, 33.22451, 33.23521, 33.24574, 33.25607, 
    33.26622, 33.27618, 33.28596, 33.29555, 33.30496, 33.31419, 33.32322, 
    33.33208, 33.34075, 33.34923, 33.35753, 33.36564, 33.37357, 33.38131, 
    33.38886, 33.39623, 33.40341, 33.41041, 33.41722, 33.42384, 33.43028, 
    33.43653, 33.4426, 33.44848, 33.45417, 33.45967, 33.465, 33.47013, 
    33.47507, 33.47983, 33.48441, 33.48879, 33.49299, 33.497, 33.50082, 
    33.50446, 33.50791, 33.51118, 33.51425, 33.51714, 33.51984, 33.52236, 
    33.52468, 33.52682, 33.52878, 33.53054, 33.53212, 33.53351, 33.53471, 
    33.53573, 33.53656, 33.5372, 33.53765, 33.53792, 33.538, 33.53789, 
    33.53759, 33.53711, 33.53644, 33.53558, 33.53454, 33.5333, 33.53188, 
    33.53028, 33.52848, 33.5265, 33.52433, 33.52197, 33.51943, 33.5167, 
    33.51378, 33.51067, 33.50738, 33.5039, 33.50023, 33.49638, 33.49234, 
    33.48811, 33.4837, 33.47909, 33.4743, 33.46933, 33.46416, 33.45882, 
    33.45328, 33.44756, 33.44165, 33.43556, 33.42928, 33.42281, 33.41615, 
    33.40931, 33.40229, 33.39508, 33.38768, 33.38009, 33.37232, 33.36437, 
    33.35623, 33.3479, 33.33939, 33.33069, 33.32181, 33.31274, 33.30349, 
    33.29405, 33.28442, 33.27462, 33.26462, 33.25444, 33.24408, 33.23354, 
    33.22281, 33.21189, 33.20079, 33.18951, 33.17804, 33.16639, 33.15455, 
    33.14253, 33.13033, 33.11795, 33.10538, 33.09263, 33.07969, 33.06657, 
    33.05328, 33.03979, 33.02613, 33.01228, 32.99825, 32.98404, 32.96965, 
    32.95507, 32.94032, 32.92538, 32.91026, 32.89496, 32.87948, 32.86382, 
    32.84797, 32.83195, 32.81574, 32.79936, 32.78279, 32.76605, 32.74913, 
    32.73203, 32.71474, 32.69728, 32.67964, 32.66182, 32.64382, 32.62564, 
    32.60728, 32.58875, 32.57004, 32.55115, 32.53208, 32.51283, 32.49341, 
    32.47381, 32.45403, 32.43408, 32.41395, 32.39364, 32.37316, 32.3525, 
    32.33167, 32.31066, 32.28947, 32.26811, 32.24657, 32.22486, 32.20298, 
    32.18092, 32.15868, 32.13628, 32.11369, 32.09094, 32.06801, 32.04491, 
    32.02163, 31.99818, 31.97456, 31.95077, 31.92681, 31.90267, 31.87836, 
    31.85388, 31.82923, 31.80441, 31.77942, 31.75425, 31.72892, 31.70341, 
    31.67774, 31.6519, 31.62589, 31.5997, 31.57335, 31.54683, 31.52015, 
    31.49329, 31.46626, 31.43907, 31.41171, 31.38419, 31.35649, 31.32863, 
    31.30061, 31.27241, 31.24405, 31.21553, 31.18684, 31.15798, 31.12896, 
    31.09978, 31.07043, 31.04091, 31.01123, 30.98139, 30.95138, 30.92121, 
    30.89088, 30.86039,
  27.45764, 27.50209, 27.54642, 27.5906, 27.63465, 27.67856, 27.72234, 
    27.76597, 27.80947, 27.85283, 27.89605, 27.93913, 27.98207, 28.02487, 
    28.06754, 28.11006, 28.15244, 28.19468, 28.23678, 28.27874, 28.32055, 
    28.36223, 28.40376, 28.44515, 28.48639, 28.5275, 28.56846, 28.60927, 
    28.64994, 28.69047, 28.73085, 28.77109, 28.81118, 28.85113, 28.89093, 
    28.93058, 28.97009, 29.00945, 29.04866, 29.08773, 29.12665, 29.16542, 
    29.20404, 29.24252, 29.28084, 29.31902, 29.35704, 29.39492, 29.43265, 
    29.47022, 29.50765, 29.54492, 29.58205, 29.61902, 29.65584, 29.69251, 
    29.72902, 29.76539, 29.8016, 29.83765, 29.87356, 29.90931, 29.9449, 
    29.98035, 30.01563, 30.05077, 30.08574, 30.12057, 30.15523, 30.18974, 
    30.22409, 30.25829, 30.29233, 30.32621, 30.35994, 30.39351, 30.42692, 
    30.46017, 30.49326, 30.5262, 30.55897, 30.59159, 30.62405, 30.65634, 
    30.68848, 30.72046, 30.75227, 30.78393, 30.81542, 30.84675, 30.87792, 
    30.90893, 30.93978, 30.97046, 31.00098, 31.03134, 31.06154, 31.09157, 
    31.12144, 31.15114, 31.18068, 31.21005, 31.23926, 31.26831, 31.29719, 
    31.3259, 31.35445, 31.38283, 31.41104, 31.43909, 31.46697, 31.49469, 
    31.52224, 31.54962, 31.57683, 31.60387, 31.63075, 31.65746, 31.684, 
    31.71037, 31.73657, 31.7626, 31.78846, 31.81415, 31.83967, 31.86502, 
    31.8902, 31.91521, 31.94005, 31.96472, 31.98922, 32.01354, 32.03769, 
    32.06167, 32.08548, 32.10911, 32.13258, 32.15586, 32.17898, 32.20192, 
    32.22469, 32.24728, 32.2697, 32.29195, 32.31402, 32.33592, 32.35764, 
    32.37919, 32.40056, 32.42175, 32.44278, 32.46362, 32.48429, 32.50478, 
    32.52509, 32.54523, 32.56519, 32.58498, 32.60458, 32.62402, 32.64326, 
    32.66234, 32.68124, 32.69995, 32.71849, 32.73685, 32.75504, 32.77304, 
    32.79086, 32.80851, 32.82597, 32.84326, 32.86037, 32.87729, 32.89404, 
    32.91061, 32.92699, 32.9432, 32.95922, 32.97506, 32.99073, 33.00621, 
    33.02151, 33.03662, 33.05156, 33.06631, 33.08089, 33.09528, 33.10949, 
    33.12352, 33.13736, 33.15102, 33.1645, 33.17779, 33.19091, 33.20383, 
    33.21658, 33.22914, 33.24152, 33.25372, 33.26573, 33.27756, 33.2892, 
    33.30066, 33.31194, 33.32302, 33.33393, 33.34465, 33.35519, 33.36554, 
    33.37571, 33.38569, 33.39549, 33.4051, 33.41453, 33.42377, 33.43282, 
    33.4417, 33.45038, 33.45888, 33.46719, 33.47532, 33.48326, 33.49101, 
    33.49858, 33.50597, 33.51316, 33.52017, 33.52699, 33.53363, 33.54008, 
    33.54634, 33.55242, 33.55831, 33.56401, 33.56953, 33.57486, 33.58, 
    33.58496, 33.58973, 33.5943, 33.5987, 33.60291, 33.60692, 33.61076, 
    33.6144, 33.61786, 33.62112, 33.62421, 33.6271, 33.62981, 33.63233, 
    33.63466, 33.6368, 33.63876, 33.64053, 33.64211, 33.64351, 33.64471, 
    33.64573, 33.64656, 33.6472, 33.64766, 33.64792, 33.648, 33.64789, 
    33.64759, 33.64711, 33.64644, 33.64558, 33.64453, 33.6433, 33.64187, 
    33.64026, 33.63846, 33.63648, 33.6343, 33.63194, 33.62939, 33.62666, 
    33.62373, 33.62062, 33.61732, 33.61383, 33.61016, 33.6063, 33.60225, 
    33.59801, 33.59359, 33.58898, 33.58419, 33.5792, 33.57403, 33.56867, 
    33.56313, 33.55739, 33.55147, 33.54536, 33.53907, 33.53259, 33.52593, 
    33.51907, 33.51204, 33.50481, 33.4974, 33.4898, 33.48201, 33.47404, 
    33.46589, 33.45755, 33.44902, 33.4403, 33.4314, 33.42232, 33.41305, 
    33.40359, 33.39395, 33.38412, 33.37411, 33.36392, 33.35353, 33.34297, 
    33.33222, 33.32128, 33.31016, 33.29886, 33.28737, 33.2757, 33.26384, 
    33.2518, 33.23957, 33.22717, 33.21458, 33.2018, 33.18884, 33.1757, 
    33.16238, 33.14887, 33.13518, 33.12131, 33.10725, 33.09302, 33.0786, 
    33.064, 33.04921, 33.03424, 33.0191, 33.00377, 32.98826, 32.97257, 
    32.9567, 32.94064, 32.92441, 32.908, 32.8914, 32.87463, 32.85767, 
    32.84054, 32.82322, 32.80573, 32.78806, 32.77021, 32.75217, 32.73396, 
    32.71557, 32.69701, 32.67826, 32.65934, 32.64023, 32.62095, 32.60149, 
    32.58186, 32.56205, 32.54206, 32.52189, 32.50155, 32.48103, 32.46033, 
    32.43946, 32.41842, 32.39719, 32.37579, 32.35422, 32.33247, 32.31054, 
    32.28844, 32.26617, 32.24372, 32.2211, 32.1983, 32.17533, 32.15219, 
    32.12888, 32.10538, 32.08172, 32.05789, 32.03388, 32.0097, 31.98535, 
    31.96083, 31.93613, 31.91127, 31.88623, 31.86102, 31.83565, 31.8101, 
    31.78438, 31.75849, 31.73243, 31.70621, 31.67981, 31.65324, 31.62651, 
    31.59961, 31.57254, 31.5453, 31.51789, 31.49032, 31.46258, 31.43467, 
    31.40659, 31.37835, 31.34994, 31.32137, 31.29263, 31.26372, 31.23465, 
    31.20542, 31.17602, 31.14645, 31.11672, 31.08683, 31.05677, 31.02655, 
    30.99617, 30.96562,
  27.55728, 27.6018, 27.64619, 27.69044, 27.73455, 27.77853, 27.82237, 
    27.86607, 27.90964, 27.95306, 27.99635, 28.03949, 28.0825, 28.12537, 
    28.16809, 28.21068, 28.25313, 28.29543, 28.3376, 28.37962, 28.4215, 
    28.46324, 28.50484, 28.54629, 28.5876, 28.62877, 28.66979, 28.71067, 
    28.7514, 28.79199, 28.83244, 28.87274, 28.91289, 28.9529, 28.99276, 
    29.03248, 29.07205, 29.11147, 29.15075, 29.18988, 29.22886, 29.26769, 
    29.30637, 29.34491, 29.3833, 29.42153, 29.45962, 29.49755, 29.53534, 
    29.57298, 29.61046, 29.6478, 29.68498, 29.72202, 29.75889, 29.79562, 
    29.8322, 29.86862, 29.90489, 29.94101, 29.97697, 30.01278, 30.04843, 
    30.08393, 30.11927, 30.15446, 30.1895, 30.22438, 30.2591, 30.29367, 
    30.32808, 30.36233, 30.39643, 30.43037, 30.46415, 30.49777, 30.53124, 
    30.56454, 30.59769, 30.63068, 30.66351, 30.69618, 30.72869, 30.76105, 
    30.79324, 30.82527, 30.85714, 30.88885, 30.92039, 30.95178, 30.983, 
    31.01406, 31.04496, 31.0757, 31.10627, 31.13668, 31.16692, 31.197, 
    31.22692, 31.25668, 31.28627, 31.31569, 31.34495, 31.37404, 31.40297, 
    31.43174, 31.46033, 31.48876, 31.51703, 31.54513, 31.57306, 31.60082, 
    31.62841, 31.65584, 31.6831, 31.71019, 31.73711, 31.76387, 31.79045, 
    31.81687, 31.84311, 31.86919, 31.8951, 31.92084, 31.9464, 31.9718, 
    31.99702, 32.02208, 32.04696, 32.07167, 32.09621, 32.12057, 32.14477, 
    32.16879, 32.19264, 32.21632, 32.23982, 32.26315, 32.2863, 32.30929, 
    32.3321, 32.35473, 32.37719, 32.39948, 32.42159, 32.44352, 32.46528, 
    32.48687, 32.50828, 32.52951, 32.55057, 32.57145, 32.59216, 32.61269, 
    32.63304, 32.65321, 32.67321, 32.69303, 32.71267, 32.73214, 32.75142, 
    32.77053, 32.78946, 32.80821, 32.82679, 32.84518, 32.8634, 32.88143, 
    32.89929, 32.91697, 32.93446, 32.95178, 32.96891, 32.98587, 33.00265, 
    33.01925, 33.03566, 33.0519, 33.06795, 33.08382, 33.09951, 33.11502, 
    33.13035, 33.14549, 33.16046, 33.17524, 33.18984, 33.20426, 33.21849, 
    33.23254, 33.24641, 33.2601, 33.2736, 33.28692, 33.30006, 33.31301, 
    33.32578, 33.33836, 33.35077, 33.36298, 33.37502, 33.38687, 33.39853, 
    33.41002, 33.42131, 33.43242, 33.44335, 33.45409, 33.46465, 33.47502, 
    33.4852, 33.4952, 33.50502, 33.51465, 33.52409, 33.53335, 33.54242, 
    33.55131, 33.56001, 33.56852, 33.57685, 33.585, 33.59295, 33.60072, 
    33.6083, 33.6157, 33.62291, 33.62993, 33.63677, 33.64342, 33.64988, 
    33.65615, 33.66224, 33.66814, 33.67385, 33.67938, 33.68472, 33.68987, 
    33.69484, 33.69962, 33.7042, 33.70861, 33.71282, 33.71685, 33.72068, 
    33.72434, 33.7278, 33.73108, 33.73417, 33.73706, 33.73978, 33.7423, 
    33.74464, 33.74678, 33.74874, 33.75051, 33.7521, 33.75349, 33.7547, 
    33.75572, 33.75655, 33.7572, 33.75765, 33.75792, 33.758, 33.75789, 
    33.7576, 33.75711, 33.75644, 33.75557, 33.75452, 33.75329, 33.75186, 
    33.75025, 33.74845, 33.74646, 33.74428, 33.74191, 33.73936, 33.73662, 
    33.73369, 33.73057, 33.72726, 33.72377, 33.72009, 33.71622, 33.71217, 
    33.70792, 33.70349, 33.69887, 33.69407, 33.68907, 33.68389, 33.67852, 
    33.67297, 33.66722, 33.66129, 33.65517, 33.64887, 33.64238, 33.6357, 
    33.62883, 33.62178, 33.61454, 33.60712, 33.5995, 33.59171, 33.58372, 
    33.57555, 33.56719, 33.55865, 33.54992, 33.541, 33.5319, 33.52261, 
    33.51314, 33.50348, 33.49363, 33.4836, 33.47339, 33.46299, 33.4524, 
    33.44163, 33.43068, 33.41954, 33.40821, 33.3967, 33.38501, 33.37313, 
    33.36106, 33.34882, 33.33639, 33.32377, 33.31097, 33.29799, 33.28483, 
    33.27148, 33.25795, 33.24423, 33.23033, 33.21625, 33.20199, 33.18754, 
    33.17291, 33.1581, 33.14311, 33.12794, 33.11258, 33.09704, 33.08132, 
    33.06542, 33.04934, 33.03308, 33.01663, 33.00001, 32.9832, 32.96622, 
    32.94905, 32.93171, 32.91418, 32.89647, 32.87859, 32.86052, 32.84228, 
    32.82386, 32.80526, 32.78648, 32.76752, 32.74838, 32.72907, 32.70958, 
    32.6899, 32.67006, 32.65003, 32.62983, 32.60945, 32.58889, 32.56816, 
    32.54725, 32.52617, 32.5049, 32.48347, 32.46185, 32.44006, 32.4181, 
    32.39596, 32.37365, 32.35116, 32.3285, 32.30566, 32.28265, 32.25947, 
    32.23611, 32.21258, 32.18888, 32.165, 32.14095, 32.11673, 32.09233, 
    32.06777, 32.04303, 32.01812, 31.99304, 31.96779, 31.94237, 31.91677, 
    31.89101, 31.86508, 31.83898, 31.8127, 31.78626, 31.75965, 31.73287, 
    31.70592, 31.6788, 31.65151, 31.62406, 31.59644, 31.56865, 31.54069, 
    31.51257, 31.48428, 31.45582, 31.4272, 31.39841, 31.36945, 31.34033, 
    31.31105, 31.2816, 31.25198, 31.2222, 31.19226, 31.16215, 31.13188, 
    31.10144, 31.07084,
  27.65689, 27.70148, 27.74594, 27.79026, 27.83444, 27.87848, 27.92239, 
    27.96615, 28.00978, 28.05327, 28.09663, 28.13984, 28.18291, 28.22584, 
    28.26864, 28.31129, 28.3538, 28.39617, 28.4384, 28.48049, 28.52243, 
    28.56423, 28.60589, 28.64741, 28.68879, 28.73001, 28.7711, 28.81205, 
    28.85284, 28.8935, 28.93401, 28.97437, 29.01459, 29.05466, 29.09458, 
    29.13436, 29.17399, 29.21348, 29.25282, 29.29201, 29.33105, 29.36994, 
    29.40869, 29.44728, 29.48573, 29.52403, 29.56218, 29.60018, 29.63802, 
    29.67572, 29.71327, 29.75066, 29.7879, 29.825, 29.86194, 29.89872, 
    29.93536, 29.97184, 30.00817, 30.04434, 30.08036, 30.11623, 30.15194, 
    30.1875, 30.2229, 30.25815, 30.29324, 30.32818, 30.36296, 30.39758, 
    30.43205, 30.46636, 30.50051, 30.53451, 30.56834, 30.60202, 30.63555, 
    30.66891, 30.70211, 30.73516, 30.76804, 30.80077, 30.83333, 30.86574, 
    30.89798, 30.93007, 30.96199, 30.99375, 31.02535, 31.05679, 31.08806, 
    31.11918, 31.15013, 31.18092, 31.21154, 31.242, 31.2723, 31.30243, 
    31.3324, 31.36221, 31.39185, 31.42132, 31.45063, 31.47977, 31.50875, 
    31.53757, 31.56621, 31.59469, 31.623, 31.65115, 31.67913, 31.70694, 
    31.73458, 31.76206, 31.78936, 31.8165, 31.84347, 31.87027, 31.8969, 
    31.92336, 31.94966, 31.97578, 32.00173, 32.02751, 32.05312, 32.07856, 
    32.10383, 32.12893, 32.15385, 32.17861, 32.20319, 32.2276, 32.25183, 
    32.2759, 32.29979, 32.32351, 32.34705, 32.37043, 32.39362, 32.41665, 
    32.4395, 32.46217, 32.48467, 32.507, 32.52915, 32.55112, 32.57292, 
    32.59454, 32.61599, 32.63726, 32.65836, 32.67928, 32.70002, 32.72058, 
    32.74097, 32.76118, 32.78122, 32.80107, 32.82075, 32.84025, 32.85957, 
    32.87872, 32.89768, 32.91647, 32.93507, 32.9535, 32.97175, 32.98981, 
    33.00771, 33.02541, 33.04294, 33.06029, 33.07746, 33.09445, 33.11126, 
    33.12788, 33.14433, 33.16059, 33.17667, 33.19257, 33.20829, 33.22383, 
    33.23919, 33.25436, 33.26935, 33.28416, 33.29879, 33.31323, 33.32749, 
    33.34157, 33.35546, 33.36917, 33.3827, 33.39605, 33.40921, 33.42218, 
    33.43498, 33.44759, 33.46001, 33.47225, 33.48431, 33.49618, 33.50787, 
    33.51937, 33.53068, 33.54181, 33.55276, 33.56352, 33.5741, 33.58449, 
    33.5947, 33.60471, 33.61455, 33.6242, 33.63366, 33.64293, 33.65202, 
    33.66092, 33.66964, 33.67817, 33.68652, 33.69467, 33.70264, 33.71043, 
    33.71803, 33.72543, 33.73266, 33.73969, 33.74654, 33.7532, 33.75968, 
    33.76596, 33.77206, 33.77797, 33.7837, 33.78924, 33.79459, 33.79975, 
    33.80472, 33.80951, 33.8141, 33.81852, 33.82273, 33.82677, 33.83062, 
    33.83427, 33.83775, 33.84103, 33.84412, 33.84702, 33.84974, 33.85227, 
    33.85461, 33.85676, 33.85873, 33.8605, 33.86209, 33.86349, 33.8647, 
    33.86572, 33.86655, 33.8672, 33.86765, 33.86792, 33.868, 33.86789, 
    33.86759, 33.86711, 33.86643, 33.86557, 33.86452, 33.86328, 33.86185, 
    33.86023, 33.85843, 33.85643, 33.85425, 33.85188, 33.84932, 33.84658, 
    33.84364, 33.84052, 33.83721, 33.83371, 33.83002, 33.82615, 33.82208, 
    33.81783, 33.81339, 33.80876, 33.80395, 33.79894, 33.79375, 33.78837, 
    33.78281, 33.77705, 33.77111, 33.76498, 33.75867, 33.75216, 33.74547, 
    33.73859, 33.73153, 33.72427, 33.71684, 33.70921, 33.70139, 33.69339, 
    33.68521, 33.67683, 33.66827, 33.65953, 33.6506, 33.64148, 33.63217, 
    33.62268, 33.613, 33.60314, 33.59309, 33.58286, 33.57244, 33.56183, 
    33.55104, 33.54007, 33.5289, 33.51756, 33.50603, 33.49431, 33.48241, 
    33.47033, 33.45806, 33.4456, 33.43296, 33.42014, 33.40714, 33.39395, 
    33.38057, 33.36702, 33.35328, 33.33936, 33.32525, 33.31096, 33.29649, 
    33.28183, 33.26699, 33.25197, 33.23677, 33.22139, 33.20582, 33.19007, 
    33.17414, 33.15803, 33.14174, 33.12526, 33.10861, 33.09177, 33.07476, 
    33.05756, 33.04018, 33.02262, 33.00489, 32.98697, 32.96887, 32.9506, 
    32.93214, 32.91351, 32.89469, 32.8757, 32.85653, 32.83718, 32.81765, 
    32.79794, 32.77806, 32.758, 32.73776, 32.71734, 32.69675, 32.67598, 
    32.65503, 32.63391, 32.61261, 32.59114, 32.56948, 32.54766, 32.52565, 
    32.50348, 32.48112, 32.4586, 32.43589, 32.41302, 32.38997, 32.36674, 
    32.34334, 32.31977, 32.29602, 32.27211, 32.24801, 32.22375, 32.19931, 
    32.1747, 32.14992, 32.12497, 32.09985, 32.07455, 32.04908, 32.02345, 
    31.99763, 31.97166, 31.94551, 31.91919, 31.8927, 31.86604, 31.83922, 
    31.81222, 31.78506, 31.75772, 31.73022, 31.70255, 31.67471, 31.64671, 
    31.61854, 31.5902, 31.56169, 31.53302, 31.50418, 31.47518, 31.446, 
    31.41667, 31.38717, 31.3575, 31.32767, 31.29768, 31.26752, 31.23719, 
    31.20671, 31.17606,
  27.75649, 27.80115, 27.84567, 27.89006, 27.9343, 27.97841, 28.02238, 
    28.06622, 28.10991, 28.15347, 28.19689, 28.24016, 28.2833, 28.3263, 
    28.36916, 28.41188, 28.45445, 28.49689, 28.53918, 28.58133, 28.62334, 
    28.66521, 28.70693, 28.74852, 28.78996, 28.83125, 28.8724, 28.91341, 
    28.95427, 28.99498, 29.03556, 29.07598, 29.11626, 29.1564, 29.19639, 
    29.23623, 29.27592, 29.31547, 29.35487, 29.39412, 29.43323, 29.47218, 
    29.51099, 29.54965, 29.58815, 29.62651, 29.66472, 29.70278, 29.74069, 
    29.77845, 29.81605, 29.85351, 29.89081, 29.92796, 29.96496, 30.00181, 
    30.0385, 30.07504, 30.11143, 30.14766, 30.18374, 30.21967, 30.25544, 
    30.29106, 30.32652, 30.36182, 30.39697, 30.43196, 30.4668, 30.50148, 
    30.53601, 30.57037, 30.60458, 30.63863, 30.67253, 30.70626, 30.73984, 
    30.77326, 30.80652, 30.83962, 30.87256, 30.90534, 30.93796, 30.97042, 
    31.00271, 31.03485, 31.06683, 31.09864, 31.1303, 31.16179, 31.19312, 
    31.22428, 31.25529, 31.28613, 31.3168, 31.34731, 31.37766, 31.40785, 
    31.43787, 31.46772, 31.49742, 31.52694, 31.5563, 31.58549, 31.61452, 
    31.64338, 31.67208, 31.70061, 31.72897, 31.75716, 31.78519, 31.81305, 
    31.84074, 31.86826, 31.89562, 31.9228, 31.94982, 31.97667, 32.00334, 
    32.02985, 32.05619, 32.08236, 32.10835, 32.13418, 32.15984, 32.18532, 
    32.21063, 32.23577, 32.26074, 32.28554, 32.31017, 32.33462, 32.3589, 
    32.383, 32.40694, 32.4307, 32.45428, 32.4777, 32.50093, 32.524, 32.54689, 
    32.56961, 32.59214, 32.61451, 32.6367, 32.65871, 32.68055, 32.70221, 
    32.7237, 32.74501, 32.76614, 32.7871, 32.80788, 32.82848, 32.84891, 
    32.86915, 32.88922, 32.90911, 32.92883, 32.94836, 32.96772, 32.9869, 
    33.00589, 33.02472, 33.04335, 33.06181, 33.0801, 33.0982, 33.11612, 
    33.13386, 33.15142, 33.1688, 33.186, 33.20302, 33.21986, 33.23652, 
    33.25299, 33.26928, 33.28539, 33.30132, 33.31707, 33.33264, 33.34802, 
    33.36322, 33.37824, 33.39308, 33.40773, 33.4222, 33.43649, 33.45059, 
    33.46451, 33.47825, 33.4918, 33.50517, 33.51836, 33.53136, 33.54417, 
    33.5568, 33.56925, 33.58152, 33.59359, 33.60549, 33.6172, 33.62872, 
    33.64006, 33.65121, 33.66217, 33.67295, 33.68355, 33.69396, 33.70419, 
    33.71422, 33.72408, 33.73374, 33.74322, 33.75251, 33.76162, 33.77054, 
    33.77927, 33.78782, 33.79618, 33.80435, 33.81234, 33.82013, 33.82774, 
    33.83517, 33.8424, 33.84945, 33.85632, 33.86299, 33.86947, 33.87577, 
    33.88189, 33.88781, 33.89354, 33.89909, 33.90445, 33.90962, 33.9146, 
    33.9194, 33.924, 33.92842, 33.93265, 33.93669, 33.94055, 33.94421, 
    33.94769, 33.95097, 33.95407, 33.95699, 33.95971, 33.96224, 33.96458, 
    33.96674, 33.96871, 33.97049, 33.97208, 33.97348, 33.97469, 33.97572, 
    33.97655, 33.9772, 33.97765, 33.97792, 33.978, 33.97789, 33.97759, 
    33.9771, 33.97643, 33.97556, 33.97451, 33.97327, 33.97184, 33.97022, 
    33.96841, 33.96641, 33.96423, 33.96185, 33.95929, 33.95654, 33.9536, 
    33.95047, 33.94715, 33.94365, 33.93995, 33.93607, 33.932, 33.92773, 
    33.92329, 33.91865, 33.91383, 33.90881, 33.90361, 33.89822, 33.89265, 
    33.88688, 33.88093, 33.87479, 33.86846, 33.86195, 33.85524, 33.84835, 
    33.84127, 33.83401, 33.82655, 33.81891, 33.81108, 33.80307, 33.79487, 
    33.78648, 33.7779, 33.76914, 33.76019, 33.75105, 33.74173, 33.73222, 
    33.72253, 33.71265, 33.70258, 33.69233, 33.68189, 33.67126, 33.66045, 
    33.64946, 33.63828, 33.62691, 33.61535, 33.60362, 33.59169, 33.57959, 
    33.5673, 33.55482, 33.54216, 33.52931, 33.51628, 33.50307, 33.48967, 
    33.47609, 33.46232, 33.44837, 33.43424, 33.41993, 33.40543, 33.39074, 
    33.37588, 33.36083, 33.3456, 33.33019, 33.31459, 33.29882, 33.28286, 
    33.26672, 33.25039, 33.23389, 33.21721, 33.20034, 33.18329, 33.16607, 
    33.14865, 33.13107, 33.1133, 33.09534, 33.07722, 33.05891, 33.04042, 
    33.02175, 33.0029, 32.98388, 32.96467, 32.94528, 32.92572, 32.90598, 
    32.88606, 32.86596, 32.84569, 32.82523, 32.8046, 32.7838, 32.76281, 
    32.74165, 32.72031, 32.6988, 32.67711, 32.65524, 32.6332, 32.61098, 
    32.58859, 32.56602, 32.54328, 32.52036, 32.49727, 32.47401, 32.45057, 
    32.42695, 32.40316, 32.3792, 32.35507, 32.33076, 32.30628, 32.28163, 
    32.25681, 32.23181, 32.20664, 32.1813, 32.15579, 32.1301, 32.10425, 
    32.07823, 32.05203, 32.02567, 31.99913, 31.97243, 31.94555, 31.91851, 
    31.8913, 31.86392, 31.83637, 31.80865, 31.78077, 31.75271, 31.72449, 
    31.69611, 31.66755, 31.63883, 31.60994, 31.58089, 31.55167, 31.52228, 
    31.49273, 31.46301, 31.43313, 31.40309, 31.37287, 31.3425, 31.31196, 
    31.28126,
  27.85607, 27.90079, 27.94538, 27.98983, 28.03415, 28.07832, 28.12236, 
    28.16626, 28.21002, 28.25364, 28.29713, 28.34047, 28.38368, 28.42674, 
    28.46966, 28.51245, 28.55509, 28.59759, 28.63995, 28.68216, 28.72424, 
    28.76617, 28.80796, 28.8496, 28.89111, 28.93246, 28.97368, 29.01475, 
    29.05567, 29.09645, 29.13709, 29.17758, 29.21792, 29.25812, 29.29817, 
    29.33808, 29.37783, 29.41744, 29.45691, 29.49622, 29.53539, 29.5744, 
    29.61327, 29.65199, 29.69056, 29.72898, 29.76725, 29.80537, 29.84334, 
    29.88116, 29.91883, 29.95634, 29.9937, 30.03091, 30.06797, 30.10488, 
    30.14163, 30.17823, 30.21468, 30.25097, 30.28711, 30.32309, 30.35892, 
    30.3946, 30.43011, 30.46548, 30.50068, 30.53574, 30.57063, 30.60537, 
    30.63995, 30.67437, 30.70864, 30.74275, 30.7767, 30.81049, 30.84412, 
    30.87759, 30.91091, 30.94406, 30.97706, 31.00989, 31.04257, 31.07508, 
    31.10744, 31.13963, 31.17166, 31.20353, 31.23523, 31.26678, 31.29816, 
    31.32938, 31.36043, 31.39132, 31.42205, 31.45262, 31.48302, 31.51325, 
    31.54333, 31.57323, 31.60297, 31.63255, 31.66196, 31.6912, 31.72028, 
    31.74919, 31.77794, 31.80651, 31.83492, 31.86317, 31.89124, 31.91915, 
    31.94689, 31.97446, 32.00186, 32.02909, 32.05616, 32.08305, 32.10978, 
    32.13633, 32.16271, 32.18892, 32.21497, 32.24084, 32.26654, 32.29207, 
    32.31742, 32.34261, 32.36763, 32.39247, 32.41713, 32.44163, 32.46595, 
    32.4901, 32.51408, 32.53788, 32.56151, 32.58496, 32.60824, 32.63135, 
    32.65428, 32.67703, 32.69962, 32.72202, 32.74425, 32.7663, 32.78818, 
    32.80988, 32.83141, 32.85275, 32.87392, 32.89492, 32.91573, 32.93637, 
    32.95683, 32.97712, 32.99722, 33.01715, 33.0369, 33.05647, 33.07586, 
    33.09507, 33.11411, 33.13296, 33.15163, 33.17013, 33.18844, 33.20657, 
    33.22453, 33.2423, 33.2599, 33.27731, 33.29454, 33.31159, 33.32846, 
    33.34514, 33.36165, 33.37797, 33.39411, 33.41007, 33.42585, 33.44144, 
    33.45686, 33.47208, 33.48713, 33.502, 33.51667, 33.53117, 33.54548, 
    33.55961, 33.57356, 33.58732, 33.6009, 33.61429, 33.6275, 33.64053, 
    33.65337, 33.66602, 33.67849, 33.69078, 33.70288, 33.71479, 33.72652, 
    33.73807, 33.74942, 33.7606, 33.77159, 33.78239, 33.793, 33.80343, 
    33.81367, 33.82373, 33.8336, 33.84328, 33.85278, 33.86209, 33.87122, 
    33.88015, 33.8889, 33.89746, 33.90584, 33.91402, 33.92202, 33.92984, 
    33.93746, 33.9449, 33.95215, 33.95921, 33.96609, 33.97277, 33.97927, 
    33.98558, 33.9917, 33.99764, 34.00338, 34.00894, 34.01431, 34.01949, 
    34.02448, 34.02929, 34.0339, 34.03833, 34.04257, 34.04662, 34.05048, 
    34.05415, 34.05763, 34.06092, 34.06403, 34.06694, 34.06967, 34.07221, 
    34.07456, 34.07672, 34.07869, 34.08047, 34.08207, 34.08347, 34.08468, 
    34.08571, 34.08654, 34.08719, 34.08765, 34.08792, 34.088, 34.08789, 
    34.08759, 34.0871, 34.08643, 34.08556, 34.0845, 34.08326, 34.08183, 
    34.0802, 34.07839, 34.07639, 34.0742, 34.07182, 34.06925, 34.0665, 
    34.06355, 34.06042, 34.05709, 34.05358, 34.04988, 34.04599, 34.04191, 
    34.03764, 34.03318, 34.02854, 34.0237, 34.01868, 34.01347, 34.00808, 
    34.00249, 33.99671, 33.99075, 33.9846, 33.97826, 33.97173, 33.96501, 
    33.95811, 33.95102, 33.94374, 33.93627, 33.92862, 33.92077, 33.91274, 
    33.90453, 33.89612, 33.88753, 33.87875, 33.86979, 33.86063, 33.85129, 
    33.84177, 33.83205, 33.82215, 33.81207, 33.80179, 33.79134, 33.78069, 
    33.76986, 33.75884, 33.74764, 33.73625, 33.72468, 33.71292, 33.70098, 
    33.68885, 33.67653, 33.66403, 33.65135, 33.63848, 33.62542, 33.61219, 
    33.59876, 33.58516, 33.57137, 33.55739, 33.54323, 33.52889, 33.51436, 
    33.49966, 33.48476, 33.46969, 33.45443, 33.43899, 33.42337, 33.40756, 
    33.39157, 33.3754, 33.35905, 33.34251, 33.3258, 33.3089, 33.29182, 
    33.27456, 33.25712, 33.2395, 33.2217, 33.20372, 33.18555, 33.16721, 
    33.14869, 33.12999, 33.11111, 33.09204, 33.0728, 33.05338, 33.03379, 
    33.01401, 32.99405, 32.97392, 32.95361, 32.93312, 32.91245, 32.89161, 
    32.87059, 32.84939, 32.82801, 32.80646, 32.78473, 32.76283, 32.74074, 
    32.71849, 32.69605, 32.67345, 32.65066, 32.6277, 32.60457, 32.58126, 
    32.55778, 32.53413, 32.5103, 32.48629, 32.46212, 32.43777, 32.41324, 
    32.38855, 32.36368, 32.33864, 32.31343, 32.28804, 32.26249, 32.23676, 
    32.21086, 32.18479, 32.15855, 32.13214, 32.10556, 32.07881, 32.05189, 
    32.0248, 31.99754, 31.97011, 31.94251, 31.91475, 31.88681, 31.85871, 
    31.83044, 31.80201, 31.7734, 31.74463, 31.71569, 31.68659, 31.65732, 
    31.62788, 31.59828, 31.56851, 31.53858, 31.50848, 31.47822, 31.44779, 
    31.4172, 31.38645,
  27.95563, 28.00042, 28.04507, 28.08959, 28.13397, 28.17822, 28.22232, 
    28.26629, 28.31011, 28.3538, 28.39735, 28.44076, 28.48403, 28.52716, 
    28.57015, 28.613, 28.6557, 28.69827, 28.74069, 28.78297, 28.82511, 
    28.86711, 28.90896, 28.95067, 28.99224, 29.03366, 29.07494, 29.11607, 
    29.15706, 29.19791, 29.23861, 29.27916, 29.31957, 29.35983, 29.39994, 
    29.43991, 29.47973, 29.5194, 29.55893, 29.5983, 29.63753, 29.67661, 
    29.71554, 29.75432, 29.79295, 29.83143, 29.86976, 29.90794, 29.94597, 
    29.98385, 30.02158, 30.05916, 30.09658, 30.13385, 30.17097, 30.20794, 
    30.24475, 30.28141, 30.31791, 30.35427, 30.39046, 30.4265, 30.46239, 
    30.49812, 30.5337, 30.56912, 30.60439, 30.6395, 30.67445, 30.70924, 
    30.74388, 30.77836, 30.81268, 30.84685, 30.88085, 30.9147, 30.94839, 
    30.98192, 31.01529, 31.0485, 31.08155, 31.11444, 31.14717, 31.17974, 
    31.21214, 31.24439, 31.27647, 31.3084, 31.34016, 31.37175, 31.40319, 
    31.43446, 31.46557, 31.49651, 31.52729, 31.55791, 31.58836, 31.61865, 
    31.64877, 31.67873, 31.70852, 31.73815, 31.76761, 31.7969, 31.82603, 
    31.85499, 31.88379, 31.91241, 31.94087, 31.96916, 31.99729, 32.02524, 
    32.05303, 32.08065, 32.1081, 32.13538, 32.16249, 32.18943, 32.2162, 
    32.2428, 32.26923, 32.29549, 32.32158, 32.34749, 32.37324, 32.39881, 
    32.42421, 32.44944, 32.4745, 32.49939, 32.5241, 32.54863, 32.573, 
    32.59719, 32.62121, 32.64505, 32.66872, 32.69222, 32.71554, 32.73869, 
    32.76166, 32.78445, 32.80708, 32.82952, 32.85179, 32.87388, 32.8958, 
    32.91754, 32.9391, 32.96049, 32.9817, 33.00273, 33.02358, 33.04426, 
    33.06475, 33.08508, 33.10522, 33.12518, 33.14497, 33.16457, 33.184, 
    33.20324, 33.22231, 33.2412, 33.25991, 33.27843, 33.29678, 33.31495, 
    33.33294, 33.35074, 33.36837, 33.38581, 33.40307, 33.42015, 33.43705, 
    33.45377, 33.4703, 33.48666, 33.50283, 33.51882, 33.53462, 33.55024, 
    33.56569, 33.58094, 33.59602, 33.61091, 33.62561, 33.64014, 33.65448, 
    33.66863, 33.6826, 33.69639, 33.70999, 33.72341, 33.73664, 33.74969, 
    33.76256, 33.77523, 33.78773, 33.80004, 33.81216, 33.8241, 33.83585, 
    33.84742, 33.8588, 33.86999, 33.881, 33.89182, 33.90245, 33.9129, 
    33.92316, 33.93324, 33.94313, 33.95283, 33.96234, 33.97167, 33.98081, 
    33.98976, 33.99853, 34.00711, 34.0155, 34.0237, 34.03172, 34.03954, 
    34.04718, 34.05463, 34.0619, 34.06897, 34.07586, 34.08256, 34.08907, 
    34.09539, 34.10152, 34.10747, 34.11322, 34.11879, 34.12417, 34.12936, 
    34.13437, 34.13918, 34.1438, 34.14824, 34.15248, 34.15654, 34.1604, 
    34.16409, 34.16757, 34.17087, 34.17398, 34.17691, 34.17964, 34.18218, 
    34.18454, 34.1867, 34.18867, 34.19046, 34.19205, 34.19346, 34.19468, 
    34.19571, 34.19654, 34.19719, 34.19765, 34.19792, 34.198, 34.19789, 
    34.19759, 34.1971, 34.19642, 34.19556, 34.1945, 34.19325, 34.19181, 
    34.19019, 34.18837, 34.18637, 34.18417, 34.18179, 34.17922, 34.17646, 
    34.1735, 34.17036, 34.16703, 34.16351, 34.15981, 34.15591, 34.15182, 
    34.14754, 34.14308, 34.13843, 34.13359, 34.12856, 34.12333, 34.11792, 
    34.11233, 34.10654, 34.10057, 34.0944, 34.08805, 34.08151, 34.07478, 
    34.06786, 34.06076, 34.05347, 34.04599, 34.03831, 34.03046, 34.02242, 
    34.01418, 34.00576, 33.99715, 33.98836, 33.97937, 33.97021, 33.96085, 
    33.95131, 33.94157, 33.93166, 33.92155, 33.91126, 33.90078, 33.89012, 
    33.87926, 33.86823, 33.85701, 33.8456, 33.834, 33.82222, 33.81025, 
    33.7981, 33.78577, 33.77324, 33.76054, 33.74764, 33.73456, 33.7213, 
    33.70786, 33.69422, 33.6804, 33.6664, 33.65222, 33.63785, 33.6233, 
    33.60856, 33.59364, 33.57854, 33.56326, 33.54779, 33.53214, 33.5163, 
    33.50028, 33.48408, 33.4677, 33.45114, 33.43439, 33.41746, 33.40035, 
    33.38306, 33.36559, 33.34793, 33.3301, 33.31209, 33.29389, 33.27552, 
    33.25696, 33.23822, 33.21931, 33.20021, 33.18093, 33.16148, 33.14185, 
    33.12204, 33.10204, 33.08187, 33.06152, 33.041, 33.02029, 32.99941, 
    32.97835, 32.95712, 32.9357, 32.91411, 32.89235, 32.8704, 32.84828, 
    32.82598, 32.80351, 32.78086, 32.75804, 32.73504, 32.71186, 32.68851, 
    32.66499, 32.6413, 32.61742, 32.59338, 32.56916, 32.54477, 32.5202, 
    32.49546, 32.47055, 32.44546, 32.4202, 32.39478, 32.36917, 32.3434, 
    32.31746, 32.29134, 32.26506, 32.2386, 32.21198, 32.18518, 32.15821, 
    32.13107, 32.10377, 32.07629, 32.04865, 32.02083, 31.99285, 31.9647, 
    31.93638, 31.9079, 31.87924, 31.85042, 31.82143, 31.79228, 31.76296, 
    31.73347, 31.70382, 31.674, 31.64402, 31.61387, 31.58356, 31.55308, 
    31.52244, 31.49163,
  28.05517, 28.10003, 28.14475, 28.18933, 28.23378, 28.27809, 28.32226, 
    28.36629, 28.41018, 28.45394, 28.49755, 28.54103, 28.58436, 28.62756, 
    28.67061, 28.71353, 28.7563, 28.79893, 28.84142, 28.88376, 28.92597, 
    28.96803, 29.00995, 29.05172, 29.09335, 29.13484, 29.17618, 29.21738, 
    29.25843, 29.29934, 29.34011, 29.38072, 29.42119, 29.46152, 29.50169, 
    29.54172, 29.58161, 29.62134, 29.66093, 29.70037, 29.73966, 29.7788, 
    29.81779, 29.85663, 29.89532, 29.93387, 29.97226, 30.0105, 30.04859, 
    30.08653, 30.12432, 30.16196, 30.19944, 30.23677, 30.27395, 30.31098, 
    30.34785, 30.38457, 30.42113, 30.45754, 30.4938, 30.5299, 30.56585, 
    30.60164, 30.63727, 30.67275, 30.70807, 30.74324, 30.77825, 30.8131, 
    30.8478, 30.88234, 30.91671, 30.95094, 30.985, 31.0189, 31.05265, 
    31.08623, 31.11966, 31.15292, 31.18603, 31.21897, 31.25176, 31.28438, 
    31.31684, 31.34914, 31.38128, 31.41326, 31.44507, 31.47672, 31.50821, 
    31.53953, 31.57069, 31.60169, 31.63252, 31.66319, 31.6937, 31.72404, 
    31.75421, 31.78422, 31.81406, 31.84374, 31.87325, 31.90259, 31.93177, 
    31.96078, 31.98963, 32.0183, 32.04681, 32.07515, 32.10332, 32.13132, 
    32.15916, 32.18682, 32.21432, 32.24165, 32.26881, 32.2958, 32.32261, 
    32.34926, 32.37573, 32.40204, 32.42817, 32.45414, 32.47993, 32.50554, 
    32.53099, 32.55626, 32.58137, 32.6063, 32.63105, 32.65563, 32.68004, 
    32.70428, 32.72834, 32.75222, 32.77594, 32.79947, 32.82283, 32.84602, 
    32.86903, 32.89187, 32.91453, 32.93702, 32.95932, 32.98146, 33.00341, 
    33.02519, 33.04679, 33.06822, 33.08947, 33.11053, 33.13142, 33.15214, 
    33.17267, 33.19303, 33.21321, 33.23321, 33.25303, 33.27267, 33.29213, 
    33.31141, 33.33051, 33.34943, 33.36818, 33.38674, 33.40512, 33.42332, 
    33.44134, 33.45918, 33.47683, 33.49431, 33.5116, 33.52871, 33.54564, 
    33.56239, 33.57896, 33.59534, 33.61154, 33.62756, 33.64339, 33.65904, 
    33.67451, 33.6898, 33.7049, 33.71982, 33.73455, 33.7491, 33.76347, 
    33.77765, 33.79165, 33.80546, 33.81908, 33.83253, 33.84579, 33.85886, 
    33.87175, 33.88445, 33.89697, 33.90929, 33.92144, 33.9334, 33.94518, 
    33.95676, 33.96816, 33.97937, 33.9904, 34.00124, 34.0119, 34.02237, 
    34.03265, 34.04274, 34.05265, 34.06237, 34.0719, 34.08125, 34.0904, 
    34.09937, 34.10815, 34.11675, 34.12516, 34.13337, 34.1414, 34.14925, 
    34.1569, 34.16436, 34.17164, 34.17873, 34.18563, 34.19234, 34.19886, 
    34.2052, 34.21134, 34.2173, 34.22306, 34.22865, 34.23404, 34.23923, 
    34.24424, 34.24907, 34.2537, 34.25814, 34.26239, 34.26646, 34.27034, 
    34.27402, 34.27752, 34.28082, 34.28394, 34.28687, 34.2896, 34.29215, 
    34.29451, 34.29668, 34.29866, 34.30045, 34.30204, 34.30345, 34.30467, 
    34.3057, 34.30654, 34.30719, 34.30765, 34.30792, 34.308, 34.30789, 
    34.30759, 34.3071, 34.30642, 34.30555, 34.30449, 34.30324, 34.3018, 
    34.30017, 34.29836, 34.29635, 34.29415, 34.29176, 34.28918, 34.28642, 
    34.28346, 34.28031, 34.27698, 34.27345, 34.26973, 34.26583, 34.26173, 
    34.25745, 34.25298, 34.24832, 34.24347, 34.23842, 34.23319, 34.22778, 
    34.22217, 34.21637, 34.21038, 34.20421, 34.19785, 34.19129, 34.18455, 
    34.17762, 34.1705, 34.1632, 34.1557, 34.14802, 34.14014, 34.13208, 
    34.12384, 34.1154, 34.10678, 34.09797, 34.08897, 34.07978, 34.0704, 
    34.06084, 34.05109, 34.04116, 34.03104, 34.02073, 34.01023, 33.99954, 
    33.98867, 33.97762, 33.96637, 33.95494, 33.94333, 33.93152, 33.91953, 
    33.90736, 33.895, 33.88245, 33.86972, 33.8568, 33.8437, 33.83041, 
    33.81694, 33.80328, 33.78944, 33.77542, 33.76121, 33.74681, 33.73223, 
    33.71747, 33.70252, 33.68739, 33.67208, 33.65658, 33.6409, 33.62503, 
    33.60899, 33.59276, 33.57635, 33.55975, 33.54298, 33.52602, 33.50888, 
    33.49155, 33.47405, 33.45636, 33.4385, 33.42045, 33.40222, 33.38381, 
    33.36522, 33.34645, 33.3275, 33.30837, 33.28906, 33.26957, 33.2499, 
    33.23006, 33.21003, 33.18982, 33.16944, 33.14887, 33.12813, 33.10721, 
    33.08612, 33.06484, 33.04339, 33.02176, 32.99995, 32.97797, 32.95581, 
    32.93347, 32.91096, 32.88827, 32.86541, 32.84237, 32.81915, 32.79576, 
    32.7722, 32.74846, 32.72454, 32.70045, 32.67619, 32.65176, 32.62715, 
    32.60236, 32.57741, 32.55228, 32.52698, 32.5015, 32.47586, 32.45004, 
    32.42405, 32.39789, 32.37156, 32.34505, 32.31838, 32.29154, 32.26452, 
    32.23734, 32.20998, 32.18246, 32.15477, 32.12691, 32.09888, 32.07068, 
    32.04231, 32.01377, 31.98507, 31.9562, 31.92717, 31.89796, 31.86859, 
    31.83905, 31.80935, 31.77948, 31.74945, 31.71925, 31.68888, 31.65835, 
    31.62766, 31.5968,
  28.15468, 28.19961, 28.2444, 28.28905, 28.33356, 28.37794, 28.42218, 
    28.46627, 28.51023, 28.55406, 28.59774, 28.64128, 28.68468, 28.72794, 
    28.77106, 28.81404, 28.85688, 28.89957, 28.94213, 28.98454, 29.02681, 
    29.06893, 29.11092, 29.15276, 29.19445, 29.236, 29.27741, 29.31867, 
    29.35979, 29.40076, 29.44159, 29.48227, 29.5228, 29.56319, 29.60343, 
    29.64352, 29.68347, 29.72326, 29.76291, 29.80241, 29.84177, 29.88097, 
    29.92002, 29.95893, 29.99768, 30.03629, 30.07474, 30.11304, 30.1512, 
    30.1892, 30.22705, 30.26474, 30.30229, 30.33968, 30.37692, 30.414, 
    30.45093, 30.48771, 30.52434, 30.56081, 30.59712, 30.63328, 30.66929, 
    30.70514, 30.74083, 30.77637, 30.81175, 30.84697, 30.88204, 30.91695, 
    30.9517, 30.9863, 31.02073, 31.05501, 31.08913, 31.12309, 31.15689, 
    31.19053, 31.22401, 31.25733, 31.29049, 31.32349, 31.35633, 31.38901, 
    31.42153, 31.45388, 31.48607, 31.5181, 31.54997, 31.58167, 31.61321, 
    31.64459, 31.67581, 31.70686, 31.73774, 31.76846, 31.79902, 31.82941, 
    31.85963, 31.88969, 31.91959, 31.94932, 31.97888, 32.00827, 32.0375, 
    32.06656, 32.09546, 32.12418, 32.15274, 32.18113, 32.20935, 32.2374, 
    32.26528, 32.293, 32.32054, 32.34792, 32.37512, 32.40215, 32.42902, 
    32.45571, 32.48223, 32.50858, 32.53476, 32.56077, 32.58661, 32.61227, 
    32.63776, 32.66308, 32.68822, 32.7132, 32.738, 32.76262, 32.78708, 
    32.81135, 32.83546, 32.85938, 32.88314, 32.90672, 32.93012, 32.95335, 
    32.9764, 32.99928, 33.02198, 33.04451, 33.06686, 33.08903, 33.11102, 
    33.13284, 33.15448, 33.17594, 33.19723, 33.21833, 33.23926, 33.26001, 
    33.28059, 33.30098, 33.32119, 33.34123, 33.36108, 33.38076, 33.40026, 
    33.41957, 33.43871, 33.45766, 33.47644, 33.49504, 33.51345, 33.53168, 
    33.54974, 33.5676, 33.58529, 33.6028, 33.62012, 33.63727, 33.65423, 
    33.67101, 33.6876, 33.70402, 33.72025, 33.73629, 33.75216, 33.76784, 
    33.78334, 33.79865, 33.81378, 33.82872, 33.84348, 33.85806, 33.87245, 
    33.88666, 33.90068, 33.91452, 33.92817, 33.94164, 33.95493, 33.96802, 
    33.98093, 33.99366, 34.0062, 34.01855, 34.03072, 34.0427, 34.0545, 
    34.0661, 34.07753, 34.08876, 34.09981, 34.11067, 34.12135, 34.13183, 
    34.14214, 34.15225, 34.16217, 34.17191, 34.18146, 34.19082, 34.2, 
    34.20898, 34.21778, 34.22639, 34.23481, 34.24305, 34.25109, 34.25895, 
    34.26662, 34.27409, 34.28138, 34.28849, 34.2954, 34.30212, 34.30866, 
    34.31501, 34.32116, 34.32713, 34.33291, 34.3385, 34.34389, 34.34911, 
    34.35413, 34.35896, 34.3636, 34.36805, 34.37231, 34.37638, 34.38026, 
    34.38396, 34.38746, 34.39077, 34.39389, 34.39683, 34.39957, 34.40212, 
    34.40448, 34.40666, 34.40864, 34.41043, 34.41203, 34.41344, 34.41467, 
    34.4157, 34.41654, 34.41719, 34.41765, 34.41792, 34.418, 34.41789, 
    34.41759, 34.4171, 34.41642, 34.41555, 34.41449, 34.41323, 34.41179, 
    34.41016, 34.40834, 34.40633, 34.40412, 34.40173, 34.39915, 34.39637, 
    34.39341, 34.39026, 34.38692, 34.38338, 34.37966, 34.37575, 34.37165, 
    34.36736, 34.36288, 34.3582, 34.35334, 34.34829, 34.34305, 34.33762, 
    34.332, 34.3262, 34.3202, 34.31401, 34.30764, 34.30107, 34.29432, 
    34.28738, 34.28024, 34.27292, 34.26542, 34.25772, 34.24983, 34.24176, 
    34.23349, 34.22504, 34.2164, 34.20757, 34.19856, 34.18935, 34.17996, 
    34.17038, 34.16061, 34.15066, 34.14052, 34.13019, 34.11967, 34.10897, 
    34.09808, 34.087, 34.07573, 34.06428, 34.05264, 34.04082, 34.02881, 
    34.01661, 34.00423, 33.99166, 33.9789, 33.96596, 33.95284, 33.93953, 
    33.92603, 33.91235, 33.89848, 33.88443, 33.87019, 33.85577, 33.84116, 
    33.82637, 33.8114, 33.79624, 33.7809, 33.76537, 33.74966, 33.73377, 
    33.71769, 33.70144, 33.68499, 33.66837, 33.65156, 33.63457, 33.6174, 
    33.60004, 33.58251, 33.56479, 33.54689, 33.52881, 33.51055, 33.49211, 
    33.47348, 33.45468, 33.4357, 33.41653, 33.39718, 33.37766, 33.35796, 
    33.33807, 33.31801, 33.29776, 33.27734, 33.25674, 33.23597, 33.21501, 
    33.19387, 33.17256, 33.15107, 33.1294, 33.10756, 33.08553, 33.06333, 
    33.04095, 33.0184, 32.99567, 32.97277, 32.94969, 32.92643, 32.903, 
    32.87939, 32.85561, 32.83165, 32.80752, 32.78322, 32.75874, 32.73409, 
    32.70926, 32.68426, 32.65909, 32.63374, 32.60822, 32.58253, 32.55667, 
    32.53063, 32.50443, 32.47805, 32.4515, 32.42478, 32.39789, 32.37083, 
    32.3436, 32.3162, 32.28862, 32.26088, 32.23298, 32.2049, 32.17665, 
    32.14823, 32.11965, 32.0909, 32.06197, 32.03289, 32.00364, 31.97421, 
    31.94462, 31.91487, 31.88495, 31.85486, 31.82461, 31.7942, 31.76361, 
    31.73287, 31.70195,
  28.25418, 28.29917, 28.34403, 28.38875, 28.43333, 28.47777, 28.52207, 
    28.56624, 28.61027, 28.65415, 28.6979, 28.74151, 28.78498, 28.8283, 
    28.87149, 28.91453, 28.95744, 29.0002, 29.04282, 29.08529, 29.12763, 
    29.16982, 29.21186, 29.25377, 29.29553, 29.33714, 29.37862, 29.41994, 
    29.46112, 29.50216, 29.54305, 29.58379, 29.62439, 29.66484, 29.70514, 
    29.7453, 29.78531, 29.82517, 29.86488, 29.90445, 29.94386, 29.98313, 
    30.02224, 30.06121, 30.10003, 30.13869, 30.17721, 30.21557, 30.25378, 
    30.29184, 30.32975, 30.36751, 30.40512, 30.44257, 30.47987, 30.51701, 
    30.554, 30.59084, 30.62753, 30.66405, 30.70043, 30.73665, 30.77271, 
    30.80862, 30.84437, 30.87997, 30.91541, 30.95069, 30.98581, 31.02078, 
    31.05559, 31.09024, 31.12473, 31.15907, 31.19324, 31.22726, 31.26112, 
    31.29482, 31.32835, 31.36173, 31.39495, 31.428, 31.4609, 31.49363, 
    31.5262, 31.55861, 31.59085, 31.62294, 31.65486, 31.68661, 31.71821, 
    31.74964, 31.78091, 31.81201, 31.84295, 31.87372, 31.90433, 31.93477, 
    31.96505, 31.99516, 32.0251, 32.05489, 32.0845, 32.11394, 32.14322, 
    32.17233, 32.20127, 32.23005, 32.25866, 32.28709, 32.31536, 32.34346, 
    32.3714, 32.39916, 32.42675, 32.45417, 32.48142, 32.5085, 32.53542, 
    32.56216, 32.58872, 32.61512, 32.64135, 32.6674, 32.69328, 32.71899, 
    32.74453, 32.76989, 32.79508, 32.8201, 32.84494, 32.86961, 32.8941, 
    32.91842, 32.94257, 32.96654, 32.99033, 33.01395, 33.0374, 33.06067, 
    33.08377, 33.10668, 33.12943, 33.15199, 33.17438, 33.19659, 33.21862, 
    33.24048, 33.26216, 33.28366, 33.30499, 33.32613, 33.3471, 33.36788, 
    33.38849, 33.40892, 33.42917, 33.44925, 33.46914, 33.48885, 33.50838, 
    33.52773, 33.5469, 33.56589, 33.5847, 33.60333, 33.62178, 33.64005, 
    33.65813, 33.67603, 33.69375, 33.71129, 33.72865, 33.74582, 33.76281, 
    33.77962, 33.79625, 33.81269, 33.82895, 33.84503, 33.86092, 33.87663, 
    33.89216, 33.9075, 33.92266, 33.93763, 33.95242, 33.96702, 33.98144, 
    33.99567, 34.00972, 34.02358, 34.03726, 34.05075, 34.06406, 34.07718, 
    34.09012, 34.10287, 34.11543, 34.12781, 34.14, 34.152, 34.16382, 
    34.17545, 34.18689, 34.19815, 34.20922, 34.2201, 34.23079, 34.2413, 
    34.25162, 34.26175, 34.27169, 34.28145, 34.29102, 34.3004, 34.30959, 
    34.31859, 34.3274, 34.33603, 34.34447, 34.35272, 34.36078, 34.36865, 
    34.37633, 34.38382, 34.39113, 34.39824, 34.40517, 34.41191, 34.41845, 
    34.42481, 34.43098, 34.43696, 34.44275, 34.44835, 34.45375, 34.45898, 
    34.464, 34.46885, 34.4735, 34.47795, 34.48222, 34.48631, 34.49019, 
    34.49389, 34.4974, 34.50072, 34.50385, 34.50679, 34.50953, 34.51209, 
    34.51446, 34.51664, 34.51862, 34.52042, 34.52202, 34.52343, 34.52466, 
    34.52569, 34.52654, 34.52719, 34.52765, 34.52792, 34.528, 34.52789, 
    34.52759, 34.5271, 34.52641, 34.52554, 34.52448, 34.52322, 34.52178, 
    34.52015, 34.51832, 34.5163, 34.5141, 34.5117, 34.50911, 34.50634, 
    34.50337, 34.50021, 34.49686, 34.49332, 34.48959, 34.48567, 34.48156, 
    34.47726, 34.47277, 34.46809, 34.46322, 34.45816, 34.45291, 34.44747, 
    34.44184, 34.43602, 34.43002, 34.42382, 34.41743, 34.41085, 34.40409, 
    34.39713, 34.38999, 34.38265, 34.37513, 34.36742, 34.35952, 34.35143, 
    34.34315, 34.33468, 34.32602, 34.31718, 34.30815, 34.29892, 34.28952, 
    34.27992, 34.27013, 34.26016, 34.25, 34.23965, 34.22911, 34.21839, 
    34.20748, 34.19638, 34.18509, 34.17362, 34.16196, 34.15012, 34.13808, 
    34.12586, 34.11346, 34.10086, 34.08809, 34.07512, 34.06197, 34.04863, 
    34.03511, 34.0214, 34.00751, 33.99343, 33.97917, 33.96472, 33.95009, 
    33.93527, 33.92027, 33.90508, 33.88971, 33.87416, 33.85842, 33.8425, 
    33.82639, 33.8101, 33.79363, 33.77698, 33.76014, 33.74312, 33.72591, 
    33.70853, 33.69096, 33.67321, 33.65528, 33.63717, 33.61887, 33.6004, 
    33.58174, 33.5629, 33.54388, 33.52468, 33.5053, 33.48574, 33.466, 
    33.44608, 33.42598, 33.4057, 33.38524, 33.3646, 33.34379, 33.3228, 
    33.30162, 33.28027, 33.25874, 33.23703, 33.21515, 33.19309, 33.17085, 
    33.14843, 33.12584, 33.10307, 33.08012, 33.057, 33.0337, 33.01023, 
    32.98658, 32.96276, 32.93876, 32.91459, 32.89024, 32.86572, 32.84102, 
    32.81615, 32.7911, 32.76589, 32.7405, 32.71494, 32.6892, 32.66329, 
    32.63721, 32.61096, 32.58453, 32.55794, 32.53117, 32.50423, 32.47712, 
    32.44984, 32.4224, 32.39478, 32.36699, 32.33903, 32.3109, 32.28261, 
    32.25414, 32.22551, 32.1967, 32.16774, 32.1386, 32.10929, 32.07982, 
    32.05019, 32.02038, 31.99041, 31.96027, 31.92997, 31.8995, 31.86886, 
    31.83806, 31.8071,
  28.35366, 28.39872, 28.44364, 28.48843, 28.53307, 28.57758, 28.62195, 
    28.66619, 28.71028, 28.75423, 28.79804, 28.84172, 28.88525, 28.92864, 
    28.9719, 29.01501, 29.05797, 29.1008, 29.14349, 29.18603, 29.22843, 
    29.27068, 29.3128, 29.35476, 29.39659, 29.43827, 29.4798, 29.5212, 
    29.56244, 29.60354, 29.6445, 29.6853, 29.72596, 29.76648, 29.80684, 
    29.84706, 29.88713, 29.92706, 29.96683, 30.00646, 30.04594, 30.08526, 
    30.12444, 30.16347, 30.20235, 30.24108, 30.27965, 30.31808, 30.35635, 
    30.39448, 30.43245, 30.47026, 30.50793, 30.54544, 30.5828, 30.62001, 
    30.65706, 30.69396, 30.7307, 30.76729, 30.80372, 30.84, 30.87612, 
    30.91209, 30.9479, 30.98355, 31.01905, 31.05439, 31.08957, 31.1246, 
    31.15947, 31.19418, 31.22873, 31.26312, 31.29735, 31.33142, 31.36534, 
    31.39909, 31.43268, 31.46611, 31.49939, 31.5325, 31.56544, 31.59823, 
    31.63086, 31.66332, 31.69562, 31.72776, 31.75974, 31.79155, 31.82319, 
    31.85468, 31.886, 31.91715, 31.94814, 31.97897, 32.00963, 32.04012, 
    32.07045, 32.10062, 32.13061, 32.16044, 32.19011, 32.2196, 32.24893, 
    32.27809, 32.30708, 32.33591, 32.36456, 32.39305, 32.42137, 32.44952, 
    32.4775, 32.50531, 32.53295, 32.56042, 32.58772, 32.61485, 32.6418, 
    32.66859, 32.69521, 32.72165, 32.74792, 32.77402, 32.79995, 32.8257, 
    32.85128, 32.87669, 32.90192, 32.92698, 32.95187, 32.97658, 33.00112, 
    33.02548, 33.04967, 33.07368, 33.09752, 33.12119, 33.14468, 33.16799, 
    33.19112, 33.21408, 33.23686, 33.25947, 33.28189, 33.30415, 33.32622, 
    33.34811, 33.36983, 33.39137, 33.41273, 33.43392, 33.45492, 33.47575, 
    33.4964, 33.51686, 33.53715, 33.55725, 33.57718, 33.59693, 33.6165, 
    33.63588, 33.65509, 33.67411, 33.69296, 33.71162, 33.7301, 33.7484, 
    33.76652, 33.78445, 33.80221, 33.81978, 33.83717, 33.85437, 33.8714, 
    33.88824, 33.90489, 33.92136, 33.93766, 33.95376, 33.96968, 33.98542, 
    34.00098, 34.01635, 34.03153, 34.04653, 34.06134, 34.07597, 34.09042, 
    34.10468, 34.11876, 34.13264, 34.14635, 34.15987, 34.17319, 34.18634, 
    34.1993, 34.21207, 34.22466, 34.23706, 34.24927, 34.2613, 34.27314, 
    34.28479, 34.29625, 34.30753, 34.31862, 34.32952, 34.34024, 34.35076, 
    34.3611, 34.37125, 34.38121, 34.39099, 34.40057, 34.40997, 34.41918, 
    34.4282, 34.43703, 34.44567, 34.45412, 34.46239, 34.47046, 34.47835, 
    34.48605, 34.49355, 34.50087, 34.508, 34.51494, 34.52169, 34.52825, 
    34.53462, 34.5408, 34.54679, 34.55259, 34.5582, 34.56362, 34.56884, 
    34.57388, 34.57874, 34.58339, 34.58786, 34.59214, 34.59623, 34.60012, 
    34.60383, 34.60735, 34.61067, 34.6138, 34.61674, 34.6195, 34.62206, 
    34.62443, 34.62661, 34.6286, 34.6304, 34.63201, 34.63343, 34.63465, 
    34.63569, 34.63653, 34.63718, 34.63765, 34.63792, 34.638, 34.63789, 
    34.63759, 34.6371, 34.63641, 34.63554, 34.63447, 34.63322, 34.63177, 
    34.63013, 34.6283, 34.62628, 34.62407, 34.62167, 34.61908, 34.61629, 
    34.61332, 34.61016, 34.6068, 34.60326, 34.59952, 34.59559, 34.59147, 
    34.58717, 34.58267, 34.57798, 34.5731, 34.56803, 34.56277, 34.55732, 
    34.55168, 34.54585, 34.53983, 34.53362, 34.52722, 34.52063, 34.51385, 
    34.50689, 34.49973, 34.49238, 34.48484, 34.47712, 34.4692, 34.46109, 
    34.4528, 34.44432, 34.43565, 34.42678, 34.41774, 34.4085, 34.39907, 
    34.38945, 34.37965, 34.36966, 34.35948, 34.34911, 34.33855, 34.32781, 
    34.31688, 34.30576, 34.29445, 34.28296, 34.27128, 34.25941, 34.24735, 
    34.23511, 34.22268, 34.21006, 34.19726, 34.18427, 34.1711, 34.15774, 
    34.14419, 34.13046, 34.11654, 34.10244, 34.08815, 34.07367, 34.05901, 
    34.04417, 34.02914, 34.01392, 33.99853, 33.98294, 33.96718, 33.95123, 
    33.93509, 33.91877, 33.90227, 33.88559, 33.86871, 33.85166, 33.83443, 
    33.81701, 33.79941, 33.78163, 33.76366, 33.74552, 33.72719, 33.70868, 
    33.68999, 33.67112, 33.65206, 33.63283, 33.61341, 33.59382, 33.57404, 
    33.55408, 33.53395, 33.51363, 33.49314, 33.47247, 33.45161, 33.43058, 
    33.40937, 33.38798, 33.36641, 33.34467, 33.32274, 33.30064, 33.27836, 
    33.25591, 33.23327, 33.21046, 33.18747, 33.16431, 33.14097, 33.11745, 
    33.09377, 33.0699, 33.04586, 33.02164, 32.99725, 32.97268, 32.94794, 
    32.92303, 32.89794, 32.87268, 32.84724, 32.82164, 32.79586, 32.7699, 
    32.74377, 32.71748, 32.69101, 32.66436, 32.63755, 32.61057, 32.58341, 
    32.55608, 32.52859, 32.50092, 32.47308, 32.44508, 32.4169, 32.38856, 
    32.36004, 32.33136, 32.30251, 32.27349, 32.2443, 32.21495, 32.18542, 
    32.15574, 32.12588, 32.09586, 32.06567, 32.03531, 32.00479, 31.9741, 
    31.94325, 31.91224,
  28.45311, 28.49824, 28.54323, 28.58808, 28.6328, 28.67737, 28.72181, 
    28.76611, 28.81027, 28.85429, 28.89817, 28.94191, 28.98551, 29.02897, 
    29.07228, 29.11546, 29.15849, 29.20139, 29.24414, 29.28675, 29.32921, 
    29.37153, 29.41371, 29.45574, 29.49763, 29.53938, 29.58098, 29.62243, 
    29.66374, 29.7049, 29.74592, 29.78679, 29.82752, 29.8681, 29.90853, 
    29.94881, 29.98894, 30.02893, 30.06877, 30.10846, 30.14799, 30.18739, 
    30.22663, 30.26572, 30.30466, 30.34345, 30.38209, 30.42057, 30.45891, 
    30.49709, 30.53512, 30.573, 30.61073, 30.6483, 30.68572, 30.72299, 
    30.7601, 30.79706, 30.83386, 30.87051, 30.907, 30.94334, 30.97952, 
    31.01555, 31.05141, 31.08713, 31.12268, 31.15808, 31.19332, 31.2284, 
    31.26333, 31.2981, 31.3327, 31.36715, 31.40144, 31.43557, 31.46954, 
    31.50335, 31.537, 31.57049, 31.60381, 31.63698, 31.66998, 31.70283, 
    31.73551, 31.76802, 31.80038, 31.83257, 31.8646, 31.89647, 31.92817, 
    31.9597, 31.99108, 32.02229, 32.05333, 32.08421, 32.11492, 32.14547, 
    32.17585, 32.20606, 32.23611, 32.26599, 32.2957, 32.32525, 32.35463, 
    32.38384, 32.41288, 32.44176, 32.47046, 32.499, 32.52737, 32.55556, 
    32.58359, 32.61145, 32.63914, 32.66666, 32.694, 32.72118, 32.74818, 
    32.77502, 32.80168, 32.82817, 32.85448, 32.88063, 32.9066, 32.9324, 
    32.95803, 32.98348, 33.00876, 33.03386, 33.05879, 33.08355, 33.10813, 
    33.13254, 33.15677, 33.18082, 33.20471, 33.22841, 33.25194, 33.2753, 
    33.29847, 33.32147, 33.34429, 33.36694, 33.38941, 33.4117, 33.43381, 
    33.45575, 33.4775, 33.49908, 33.52048, 33.5417, 33.56274, 33.58361, 
    33.60429, 33.62479, 33.64512, 33.66526, 33.68523, 33.70501, 33.72461, 
    33.74403, 33.76327, 33.78233, 33.80121, 33.81991, 33.83842, 33.85675, 
    33.8749, 33.89287, 33.91066, 33.92826, 33.94568, 33.96292, 33.97997, 
    33.99685, 34.01353, 34.03003, 34.04635, 34.06249, 34.07844, 34.09421, 
    34.10979, 34.12519, 34.1404, 34.15543, 34.17027, 34.18493, 34.1994, 
    34.21369, 34.22779, 34.2417, 34.25543, 34.26897, 34.28233, 34.2955, 
    34.30848, 34.32128, 34.33389, 34.34631, 34.35855, 34.37059, 34.38245, 
    34.39413, 34.40561, 34.41691, 34.42802, 34.43895, 34.44968, 34.46022, 
    34.47058, 34.48075, 34.49073, 34.50052, 34.51013, 34.51954, 34.52877, 
    34.5378, 34.54665, 34.55531, 34.56378, 34.57206, 34.58015, 34.58805, 
    34.59576, 34.60328, 34.61061, 34.61776, 34.62471, 34.63147, 34.63804, 
    34.64442, 34.65062, 34.65662, 34.66243, 34.66805, 34.67348, 34.67871, 
    34.68377, 34.68862, 34.69329, 34.69777, 34.70205, 34.70615, 34.71005, 
    34.71376, 34.71729, 34.72062, 34.72376, 34.72671, 34.72947, 34.73203, 
    34.73441, 34.73659, 34.73859, 34.74039, 34.742, 34.74342, 34.74465, 
    34.74568, 34.74653, 34.74718, 34.74765, 34.74792, 34.748, 34.74789, 
    34.74759, 34.74709, 34.74641, 34.74553, 34.74446, 34.74321, 34.74176, 
    34.74012, 34.73828, 34.73626, 34.73404, 34.73164, 34.72904, 34.72625, 
    34.72327, 34.7201, 34.71674, 34.71319, 34.70945, 34.70551, 34.70139, 
    34.69707, 34.69256, 34.68787, 34.68298, 34.6779, 34.67263, 34.66717, 
    34.66152, 34.65568, 34.64965, 34.64342, 34.63702, 34.63041, 34.62362, 
    34.61664, 34.60947, 34.6021, 34.59455, 34.58681, 34.57888, 34.57076, 
    34.56245, 34.55396, 34.54527, 34.53639, 34.52732, 34.51807, 34.50862, 
    34.49899, 34.48917, 34.47916, 34.46896, 34.45857, 34.44799, 34.43723, 
    34.42628, 34.41514, 34.40381, 34.39229, 34.38059, 34.3687, 34.35662, 
    34.34436, 34.33191, 34.31927, 34.30644, 34.29343, 34.28023, 34.26684, 
    34.25327, 34.23951, 34.22557, 34.21144, 34.19712, 34.18262, 34.16793, 
    34.15306, 34.138, 34.12276, 34.10734, 34.09172, 34.07593, 34.05995, 
    34.04379, 34.02744, 34.0109, 33.99419, 33.97729, 33.96021, 33.94294, 
    33.92549, 33.90786, 33.89004, 33.87204, 33.85387, 33.8355, 33.81696, 
    33.79824, 33.77933, 33.76024, 33.74097, 33.72152, 33.70189, 33.68208, 
    33.66209, 33.64191, 33.62156, 33.60103, 33.58032, 33.55943, 33.53836, 
    33.51711, 33.49568, 33.47407, 33.45229, 33.43032, 33.40818, 33.38586, 
    33.36337, 33.34069, 33.31784, 33.29482, 33.27161, 33.24823, 33.22467, 
    33.20094, 33.17703, 33.15295, 33.12869, 33.10426, 33.07965, 33.05486, 
    33.0299, 33.00477, 32.97947, 32.95398, 32.92833, 32.9025, 32.87651, 
    32.85033, 32.82399, 32.79747, 32.77078, 32.74392, 32.71689, 32.68969, 
    32.66232, 32.63477, 32.60706, 32.57917, 32.55112, 32.52289, 32.4945, 
    32.46593, 32.4372, 32.4083, 32.37923, 32.34999, 32.32059, 32.29102, 
    32.26127, 32.23137, 32.20129, 32.17105, 32.14064, 32.11007, 32.07933, 
    32.04843, 32.01736,
  28.55255, 28.59774, 28.6428, 28.68772, 28.7325, 28.77714, 28.82165, 
    28.86601, 28.91024, 28.95433, 28.99827, 29.04208, 29.08574, 29.12927, 
    29.17265, 29.21589, 29.259, 29.30195, 29.34477, 29.38744, 29.42997, 
    29.47236, 29.5146, 29.5567, 29.59865, 29.64046, 29.68213, 29.72365, 
    29.76502, 29.80625, 29.84733, 29.88827, 29.92905, 29.9697, 30.01019, 
    30.05054, 30.09073, 30.13078, 30.17068, 30.21044, 30.25004, 30.28949, 
    30.32879, 30.36795, 30.40695, 30.4458, 30.4845, 30.52305, 30.56145, 
    30.59969, 30.63778, 30.67572, 30.71351, 30.75114, 30.78863, 30.82595, 
    30.86312, 30.90014, 30.937, 30.97371, 31.01027, 31.04666, 31.0829, 
    31.11899, 31.15491, 31.19069, 31.2263, 31.26176, 31.29705, 31.3322, 
    31.36718, 31.402, 31.43667, 31.47117, 31.50552, 31.5397, 31.57373, 
    31.6076, 31.6413, 31.67484, 31.70823, 31.74145, 31.77451, 31.80741, 
    31.84014, 31.87271, 31.90512, 31.93737, 31.96945, 32.00137, 32.03313, 
    32.06472, 32.09615, 32.12741, 32.1585, 32.18943, 32.2202, 32.2508, 
    32.28123, 32.31149, 32.34159, 32.37152, 32.40129, 32.43089, 32.46032, 
    32.48958, 32.51867, 32.5476, 32.57635, 32.60494, 32.63335, 32.6616, 
    32.68968, 32.71758, 32.74532, 32.77288, 32.80028, 32.8275, 32.85456, 
    32.88144, 32.90814, 32.93468, 32.96104, 32.98723, 33.01325, 33.0391, 
    33.06477, 33.09026, 33.11559, 33.14074, 33.16571, 33.19051, 33.21513, 
    33.23959, 33.26386, 33.28796, 33.31188, 33.33563, 33.3592, 33.3826, 
    33.40581, 33.42885, 33.45172, 33.4744, 33.49691, 33.51924, 33.54139, 
    33.56337, 33.58517, 33.60678, 33.62822, 33.64948, 33.67056, 33.69146, 
    33.71218, 33.73272, 33.75308, 33.77326, 33.79326, 33.81308, 33.83272, 
    33.85218, 33.87145, 33.89054, 33.90946, 33.92819, 33.94674, 33.9651, 
    33.98329, 34.00129, 34.0191, 34.03674, 34.05419, 34.07146, 34.08855, 
    34.10545, 34.12217, 34.1387, 34.15505, 34.17122, 34.18719, 34.20299, 
    34.2186, 34.23403, 34.24927, 34.26432, 34.27919, 34.29388, 34.30838, 
    34.32269, 34.33681, 34.35076, 34.36451, 34.37808, 34.39146, 34.40465, 
    34.41766, 34.43048, 34.44311, 34.45556, 34.46782, 34.47989, 34.49177, 
    34.50346, 34.51497, 34.52629, 34.53742, 34.54837, 34.55912, 34.56968, 
    34.58006, 34.59025, 34.60025, 34.61006, 34.61968, 34.62911, 34.63836, 
    34.64741, 34.65627, 34.66495, 34.67344, 34.68173, 34.68983, 34.69775, 
    34.70547, 34.71301, 34.72036, 34.72751, 34.73448, 34.74125, 34.74783, 
    34.75423, 34.76043, 34.76645, 34.77227, 34.7779, 34.78334, 34.78859, 
    34.79364, 34.79851, 34.80319, 34.80767, 34.81197, 34.81607, 34.81998, 
    34.8237, 34.82723, 34.83057, 34.83371, 34.83667, 34.83943, 34.842, 
    34.84438, 34.84657, 34.84857, 34.85037, 34.85199, 34.85341, 34.85464, 
    34.85568, 34.85653, 34.85718, 34.85765, 34.85792, 34.858, 34.85789, 
    34.85759, 34.85709, 34.85641, 34.85553, 34.85446, 34.8532, 34.85175, 
    34.8501, 34.84826, 34.84624, 34.84402, 34.84161, 34.839, 34.83621, 
    34.83323, 34.83005, 34.82668, 34.82312, 34.81937, 34.81543, 34.8113, 
    34.80698, 34.80246, 34.79775, 34.79285, 34.78777, 34.78249, 34.77702, 
    34.77136, 34.76551, 34.75946, 34.75323, 34.74681, 34.74019, 34.73339, 
    34.72639, 34.71921, 34.71183, 34.70427, 34.69651, 34.68856, 34.68043, 
    34.6721, 34.66359, 34.65488, 34.64599, 34.63691, 34.62763, 34.61817, 
    34.60852, 34.59868, 34.58865, 34.57843, 34.56803, 34.55743, 34.54665, 
    34.53568, 34.52451, 34.51316, 34.50163, 34.4899, 34.47799, 34.46589, 
    34.4536, 34.44113, 34.42846, 34.41562, 34.40258, 34.38935, 34.37594, 
    34.36235, 34.34856, 34.33459, 34.32044, 34.3061, 34.29157, 34.27686, 
    34.26196, 34.24687, 34.2316, 34.21614, 34.2005, 34.18468, 34.16867, 
    34.15247, 34.1361, 34.11953, 34.10279, 34.08586, 34.06874, 34.05145, 
    34.03396, 34.0163, 33.99845, 33.98042, 33.96221, 33.94381, 33.92524, 
    33.90648, 33.88754, 33.86842, 33.84911, 33.82962, 33.80996, 33.79011, 
    33.77008, 33.74987, 33.72948, 33.70892, 33.68817, 33.66724, 33.64613, 
    33.62484, 33.60337, 33.58173, 33.55991, 33.5379, 33.51572, 33.49336, 
    33.47083, 33.44811, 33.42522, 33.40215, 33.37891, 33.35548, 33.33189, 
    33.30811, 33.28416, 33.26003, 33.23573, 33.21125, 33.1866, 33.16177, 
    33.13677, 33.11159, 33.08624, 33.06072, 33.03502, 33.00915, 32.9831, 
    32.95688, 32.93049, 32.90393, 32.87719, 32.85029, 32.82321, 32.79596, 
    32.76854, 32.74094, 32.71318, 32.68525, 32.65714, 32.62887, 32.60043, 
    32.57181, 32.54303, 32.51408, 32.48496, 32.45567, 32.42622, 32.3966, 
    32.3668, 32.33684, 32.30672, 32.27642, 32.24597, 32.21534, 32.18455, 
    32.15359, 32.12247,
  28.65196, 28.69722, 28.74235, 28.78733, 28.83218, 28.87689, 28.92146, 
    28.9659, 29.01019, 29.05434, 29.09836, 29.14223, 29.18596, 29.22955, 
    29.273, 29.31631, 29.35948, 29.4025, 29.44538, 29.48812, 29.53072, 
    29.57317, 29.61547, 29.65764, 29.69966, 29.74153, 29.78326, 29.82485, 
    29.86628, 29.90758, 29.94872, 29.98972, 30.03057, 30.07128, 30.11184, 
    30.15224, 30.19251, 30.23262, 30.27258, 30.3124, 30.35206, 30.39158, 
    30.43094, 30.47016, 30.50922, 30.54814, 30.5869, 30.62551, 30.66397, 
    30.70228, 30.74043, 30.77843, 30.81628, 30.85397, 30.89151, 30.9289, 
    30.96613, 31.00321, 31.04013, 31.0769, 31.11351, 31.14997, 31.18627, 
    31.22241, 31.2584, 31.29423, 31.3299, 31.36542, 31.40077, 31.43597, 
    31.47101, 31.50589, 31.54062, 31.57518, 31.60958, 31.64382, 31.67791, 
    31.71183, 31.74559, 31.77919, 31.81263, 31.84591, 31.87902, 31.91198, 
    31.94477, 31.97739, 32.00986, 32.04216, 32.0743, 32.10627, 32.13808, 
    32.16972, 32.2012, 32.23251, 32.26366, 32.29465, 32.32546, 32.35611, 
    32.3866, 32.41692, 32.44707, 32.47705, 32.50687, 32.53651, 32.56599, 
    32.59531, 32.62445, 32.65342, 32.68223, 32.71087, 32.73933, 32.76763, 
    32.79575, 32.82371, 32.85149, 32.8791, 32.90655, 32.93382, 32.96092, 
    32.98785, 33.0146, 33.04118, 33.06759, 33.09383, 33.11989, 33.14578, 
    33.1715, 33.19704, 33.22241, 33.2476, 33.27262, 33.29746, 33.32213, 
    33.34663, 33.37094, 33.39508, 33.41905, 33.44284, 33.46645, 33.48989, 
    33.51315, 33.53623, 33.55914, 33.58186, 33.60441, 33.62678, 33.64897, 
    33.67099, 33.69282, 33.71448, 33.73595, 33.75725, 33.77837, 33.79931, 
    33.82006, 33.84064, 33.86104, 33.88126, 33.90129, 33.92115, 33.94082, 
    33.96032, 33.97963, 33.99875, 34.0177, 34.03646, 34.05505, 34.07345, 
    34.09166, 34.1097, 34.12755, 34.14521, 34.1627, 34.18, 34.19712, 
    34.21405, 34.2308, 34.24736, 34.26374, 34.27993, 34.29594, 34.31177, 
    34.32741, 34.34286, 34.35813, 34.37321, 34.38811, 34.40282, 34.41735, 
    34.43169, 34.44584, 34.45981, 34.47359, 34.48718, 34.50059, 34.51381, 
    34.52684, 34.53968, 34.55234, 34.5648, 34.57709, 34.58918, 34.60109, 
    34.6128, 34.62433, 34.63567, 34.64682, 34.65778, 34.66856, 34.67914, 
    34.68954, 34.69975, 34.70977, 34.71959, 34.72923, 34.73868, 34.74794, 
    34.75702, 34.7659, 34.77459, 34.78309, 34.7914, 34.79952, 34.80745, 
    34.81519, 34.82274, 34.8301, 34.83727, 34.84424, 34.85103, 34.85763, 
    34.86403, 34.87025, 34.87627, 34.8821, 34.88774, 34.8932, 34.89845, 
    34.90352, 34.9084, 34.91308, 34.91758, 34.92188, 34.92599, 34.92991, 
    34.93364, 34.93717, 34.94051, 34.94366, 34.94662, 34.94939, 34.95197, 
    34.95436, 34.95655, 34.95855, 34.96036, 34.96198, 34.9634, 34.96463, 
    34.96568, 34.96652, 34.96718, 34.96765, 34.96792, 34.968, 34.96789, 
    34.96759, 34.96709, 34.9664, 34.96552, 34.96445, 34.96319, 34.96173, 
    34.96009, 34.95824, 34.95621, 34.95399, 34.95158, 34.94897, 34.94617, 
    34.94318, 34.94, 34.93662, 34.93306, 34.9293, 34.92535, 34.92121, 
    34.91688, 34.91235, 34.90764, 34.90273, 34.89764, 34.89235, 34.88686, 
    34.8812, 34.87533, 34.86928, 34.86303, 34.8566, 34.84997, 34.84315, 
    34.83614, 34.82895, 34.82156, 34.81398, 34.80621, 34.79825, 34.7901, 
    34.78175, 34.77322, 34.7645, 34.75559, 34.74649, 34.7372, 34.72772, 
    34.71805, 34.70819, 34.69815, 34.68791, 34.67748, 34.66687, 34.65606, 
    34.64507, 34.63389, 34.62252, 34.61096, 34.59921, 34.58728, 34.57516, 
    34.56285, 34.55035, 34.53766, 34.52479, 34.51173, 34.49848, 34.48504, 
    34.47142, 34.45761, 34.44361, 34.42944, 34.41507, 34.40051, 34.38577, 
    34.37084, 34.35573, 34.34043, 34.32495, 34.30928, 34.29343, 34.27739, 
    34.26116, 34.24475, 34.22816, 34.21138, 34.19442, 34.17728, 34.15995, 
    34.14243, 34.12474, 34.10686, 34.08879, 34.07055, 34.05212, 34.03351, 
    34.01472, 33.99574, 33.97658, 33.95724, 33.93772, 33.91802, 33.89814, 
    33.87807, 33.85783, 33.8374, 33.8168, 33.79601, 33.77504, 33.75389, 
    33.73257, 33.71106, 33.68938, 33.66751, 33.64547, 33.62325, 33.60086, 
    33.57828, 33.55552, 33.53259, 33.50948, 33.48619, 33.46273, 33.43909, 
    33.41527, 33.39128, 33.36711, 33.34276, 33.31824, 33.29354, 33.26867, 
    33.24363, 33.21841, 33.19301, 33.16744, 33.1417, 33.11578, 33.08969, 
    33.06343, 33.03699, 33.01038, 32.9836, 32.95664, 32.92952, 32.90222, 
    32.87475, 32.84711, 32.8193, 32.79131, 32.76316, 32.73484, 32.70635, 
    32.67768, 32.64885, 32.61985, 32.59068, 32.56134, 32.53184, 32.50216, 
    32.47232, 32.44231, 32.41213, 32.38179, 32.35128, 32.3206, 32.28976, 
    32.25875, 32.22757,
  28.75135, 28.79668, 28.84188, 28.88693, 28.93185, 28.97662, 29.02126, 
    29.06576, 29.11012, 29.15434, 29.19842, 29.24236, 29.28616, 29.32981, 
    29.37333, 29.41671, 29.45994, 29.50303, 29.54597, 29.58878, 29.63144, 
    29.67396, 29.71633, 29.75856, 29.80064, 29.84258, 29.88438, 29.92603, 
    29.96753, 30.00888, 30.05009, 30.09116, 30.13207, 30.17284, 30.21346, 
    30.25394, 30.29426, 30.33444, 30.37447, 30.41434, 30.45407, 30.49365, 
    30.53308, 30.57236, 30.61148, 30.65046, 30.68928, 30.72795, 30.76647, 
    30.80484, 30.84306, 30.88112, 30.91903, 30.95679, 30.99439, 31.03183, 
    31.06913, 31.10626, 31.14325, 31.18007, 31.21675, 31.25326, 31.28962, 
    31.32582, 31.36187, 31.39776, 31.43349, 31.46906, 31.50448, 31.53973, 
    31.57483, 31.60977, 31.64455, 31.67917, 31.71363, 31.74793, 31.78207, 
    31.81605, 31.84987, 31.88352, 31.91702, 31.95035, 31.98352, 32.01653, 
    32.04938, 32.08206, 32.11458, 32.14693, 32.17912, 32.21115, 32.24301, 
    32.27471, 32.30624, 32.33761, 32.36881, 32.39985, 32.43072, 32.46142, 
    32.49196, 32.52233, 32.55253, 32.58257, 32.61243, 32.64213, 32.67167, 
    32.70103, 32.73022, 32.75924, 32.7881, 32.81678, 32.8453, 32.87364, 
    32.90182, 32.92982, 32.95765, 32.98532, 33.01281, 33.04012, 33.06727, 
    33.09425, 33.12105, 33.14767, 33.17413, 33.20041, 33.22652, 33.25246, 
    33.27822, 33.30381, 33.32922, 33.35446, 33.37952, 33.40441, 33.42912, 
    33.45366, 33.47802, 33.5022, 33.52621, 33.55005, 33.5737, 33.59718, 
    33.62048, 33.6436, 33.66655, 33.68931, 33.7119, 33.73431, 33.75655, 
    33.7786, 33.80047, 33.82217, 33.84369, 33.86502, 33.88617, 33.90715, 
    33.92795, 33.94856, 33.96899, 33.98925, 34.00932, 34.02921, 34.04892, 
    34.06845, 34.0878, 34.10696, 34.12594, 34.14474, 34.16335, 34.18179, 
    34.20004, 34.21811, 34.23599, 34.25368, 34.2712, 34.28854, 34.30568, 
    34.32265, 34.33942, 34.35602, 34.37243, 34.38865, 34.40469, 34.42055, 
    34.43621, 34.4517, 34.467, 34.48211, 34.49703, 34.51177, 34.52632, 
    34.54069, 34.55487, 34.56886, 34.58266, 34.59628, 34.60971, 34.62296, 
    34.63601, 34.64888, 34.66156, 34.67405, 34.68636, 34.69847, 34.7104, 
    34.72213, 34.73368, 34.74504, 34.75622, 34.7672, 34.778, 34.7886, 
    34.79902, 34.80924, 34.81928, 34.82913, 34.83878, 34.84825, 34.85753, 
    34.86662, 34.87551, 34.88422, 34.89274, 34.90107, 34.9092, 34.91714, 
    34.9249, 34.93246, 34.93984, 34.94702, 34.95401, 34.96081, 34.96742, 
    34.97384, 34.98006, 34.9861, 34.99194, 34.99759, 35.00306, 35.00832, 
    35.0134, 35.01829, 35.02298, 35.02748, 35.03179, 35.03591, 35.03984, 
    35.04357, 35.04711, 35.05046, 35.05362, 35.05659, 35.05936, 35.06194, 
    35.06433, 35.06653, 35.06853, 35.07034, 35.07196, 35.07339, 35.07463, 
    35.07567, 35.07652, 35.07718, 35.07764, 35.07792, 35.078, 35.07789, 
    35.07758, 35.07709, 35.0764, 35.07552, 35.07444, 35.07318, 35.07172, 
    35.07007, 35.06823, 35.06619, 35.06396, 35.06155, 35.05893, 35.05613, 
    35.05313, 35.04995, 35.04657, 35.04299, 35.03923, 35.03527, 35.03112, 
    35.02678, 35.02225, 35.01752, 35.01261, 35.0075, 35.0022, 34.99671, 
    34.99103, 34.98516, 34.97909, 34.97284, 34.96639, 34.95975, 34.95292, 
    34.9459, 34.93868, 34.93128, 34.92369, 34.9159, 34.90793, 34.89976, 
    34.8914, 34.88286, 34.87412, 34.86519, 34.85608, 34.84677, 34.83727, 
    34.82758, 34.81771, 34.80764, 34.79738, 34.78694, 34.7763, 34.76548, 
    34.75446, 34.74326, 34.73187, 34.72029, 34.70852, 34.69656, 34.68442, 
    34.67208, 34.65956, 34.64685, 34.63396, 34.62087, 34.6076, 34.59414, 
    34.58049, 34.56666, 34.55264, 34.53843, 34.52403, 34.50945, 34.49468, 
    34.47973, 34.46459, 34.44926, 34.43375, 34.41805, 34.40217, 34.3861, 
    34.36985, 34.3534, 34.33678, 34.31998, 34.30298, 34.2858, 34.26844, 
    34.2509, 34.23317, 34.21526, 34.19716, 34.17888, 34.16042, 34.14178, 
    34.12295, 34.10394, 34.08475, 34.06537, 34.04581, 34.02608, 34.00616, 
    33.98606, 33.96577, 33.94531, 33.92467, 33.90385, 33.88284, 33.86166, 
    33.84029, 33.81875, 33.79702, 33.77512, 33.75304, 33.73078, 33.70834, 
    33.68572, 33.66293, 33.63995, 33.6168, 33.59348, 33.56997, 33.54629, 
    33.52243, 33.49839, 33.47418, 33.44979, 33.42522, 33.40048, 33.37557, 
    33.35048, 33.32521, 33.29977, 33.27416, 33.24837, 33.2224, 33.19627, 
    33.16996, 33.14347, 33.11682, 33.08999, 33.06299, 33.03582, 33.00847, 
    32.98095, 32.95326, 32.9254, 32.89737, 32.86917, 32.8408, 32.81226, 
    32.78355, 32.75467, 32.72561, 32.69639, 32.667, 32.63745, 32.60772, 
    32.57783, 32.54776, 32.51754, 32.48714, 32.45658, 32.42585, 32.39495, 
    32.36389, 32.33266,
  28.85073, 28.89612, 28.94138, 28.9865, 29.03149, 29.07633, 29.12104, 
    29.1656, 29.21003, 29.25432, 29.29846, 29.34247, 29.38634, 29.43006, 
    29.47364, 29.51708, 29.56038, 29.60353, 29.64655, 29.68942, 29.73214, 
    29.77473, 29.81717, 29.85946, 29.90161, 29.94361, 29.98547, 30.02719, 
    30.06875, 30.11017, 30.15145, 30.19258, 30.23356, 30.27439, 30.31507, 
    30.35561, 30.396, 30.43624, 30.47633, 30.51627, 30.55606, 30.5957, 
    30.63519, 30.67453, 30.71372, 30.75276, 30.79165, 30.83038, 30.86896, 
    30.90739, 30.94567, 30.98379, 31.02176, 31.05958, 31.09724, 31.13475, 
    31.1721, 31.2093, 31.24635, 31.28323, 31.31996, 31.35654, 31.39296, 
    31.42922, 31.46532, 31.50127, 31.53706, 31.57269, 31.60817, 31.64348, 
    31.67864, 31.71363, 31.74847, 31.78315, 31.81767, 31.85202, 31.88622, 
    31.92026, 31.95413, 31.98784, 32.02139, 32.05478, 32.08801, 32.12107, 
    32.15397, 32.18671, 32.21928, 32.25169, 32.28394, 32.31602, 32.34794, 
    32.37969, 32.41128, 32.4427, 32.47395, 32.50504, 32.53596, 32.56672, 
    32.59731, 32.62773, 32.65799, 32.68807, 32.71799, 32.74774, 32.77732, 
    32.80674, 32.83598, 32.86505, 32.89396, 32.92269, 32.95126, 32.97965, 
    33.00787, 33.03593, 33.06381, 33.09152, 33.11906, 33.14642, 33.17361, 
    33.20064, 33.22749, 33.25416, 33.28066, 33.30699, 33.33315, 33.35913, 
    33.38493, 33.41057, 33.43602, 33.46131, 33.48642, 33.51135, 33.5361, 
    33.56068, 33.58509, 33.60931, 33.63337, 33.65724, 33.68094, 33.70446, 
    33.7278, 33.75097, 33.77395, 33.79676, 33.81939, 33.84184, 33.86411, 
    33.8862, 33.90812, 33.92985, 33.9514, 33.97278, 33.99397, 34.01499, 
    34.03582, 34.05647, 34.07695, 34.09723, 34.11734, 34.13727, 34.15702, 
    34.17658, 34.19596, 34.21516, 34.23417, 34.25301, 34.27166, 34.29012, 
    34.30841, 34.32651, 34.34442, 34.36215, 34.3797, 34.39706, 34.41425, 
    34.43124, 34.44805, 34.46468, 34.48111, 34.49737, 34.51344, 34.52932, 
    34.54502, 34.56053, 34.57586, 34.59099, 34.60595, 34.62071, 34.63529, 
    34.64968, 34.66389, 34.67791, 34.69174, 34.70538, 34.71883, 34.7321, 
    34.74518, 34.75808, 34.77078, 34.78329, 34.79562, 34.80776, 34.81971, 
    34.83147, 34.84304, 34.85442, 34.86562, 34.87662, 34.88743, 34.89806, 
    34.90849, 34.91874, 34.92879, 34.93866, 34.94833, 34.95782, 34.96711, 
    34.97622, 34.98513, 34.99386, 35.00239, 35.01073, 35.01888, 35.02684, 
    35.03461, 35.04219, 35.04958, 35.05677, 35.06378, 35.07059, 35.07721, 
    35.08364, 35.08988, 35.09592, 35.10178, 35.10744, 35.11291, 35.11819, 
    35.12328, 35.12817, 35.13288, 35.13739, 35.1417, 35.14583, 35.14977, 
    35.1535, 35.15705, 35.16041, 35.16357, 35.16655, 35.16932, 35.17191, 
    35.1743, 35.17651, 35.17851, 35.18033, 35.18195, 35.18338, 35.18462, 
    35.18567, 35.18652, 35.18718, 35.18764, 35.18792, 35.188, 35.18789, 
    35.18758, 35.18709, 35.1864, 35.18551, 35.18444, 35.18317, 35.18171, 
    35.18005, 35.17821, 35.17617, 35.17394, 35.17152, 35.1689, 35.16609, 
    35.16309, 35.15989, 35.15651, 35.15293, 35.14915, 35.14519, 35.14103, 
    35.13668, 35.13214, 35.12741, 35.12249, 35.11737, 35.11206, 35.10656, 
    35.10086, 35.09498, 35.08891, 35.08264, 35.07618, 35.06953, 35.06268, 
    35.05565, 35.04842, 35.041, 35.0334, 35.0256, 35.0176, 35.00943, 
    35.00105, 34.99249, 34.98374, 34.97479, 34.96566, 34.95633, 34.94682, 
    34.93711, 34.92722, 34.91713, 34.90686, 34.89639, 34.88573, 34.87489, 
    34.86386, 34.85263, 34.84122, 34.82962, 34.81783, 34.80585, 34.79368, 
    34.78133, 34.76878, 34.75605, 34.74313, 34.73001, 34.71672, 34.70324, 
    34.68956, 34.6757, 34.66166, 34.64742, 34.633, 34.61839, 34.60359, 
    34.58861, 34.57344, 34.55809, 34.54255, 34.52682, 34.51091, 34.49481, 
    34.47853, 34.46206, 34.4454, 34.42856, 34.41154, 34.39433, 34.37694, 
    34.35936, 34.3416, 34.32365, 34.30553, 34.28721, 34.26872, 34.25004, 
    34.23118, 34.21213, 34.19291, 34.1735, 34.1539, 34.13413, 34.11417, 
    34.09404, 34.07372, 34.05322, 34.03254, 34.01168, 33.99063, 33.96941, 
    33.94801, 33.92643, 33.90466, 33.88272, 33.8606, 33.8383, 33.81582, 
    33.79316, 33.77032, 33.74731, 33.72412, 33.70075, 33.6772, 33.65348, 
    33.62957, 33.6055, 33.58124, 33.55681, 33.5322, 33.50742, 33.48246, 
    33.45732, 33.43201, 33.40652, 33.38086, 33.35503, 33.32902, 33.30284, 
    33.27648, 33.24995, 33.22325, 33.19637, 33.16933, 33.14211, 33.11471, 
    33.08715, 33.05941, 33.0315, 33.00342, 32.97517, 32.94675, 32.91816, 
    32.8894, 32.86047, 32.83136, 32.80209, 32.77265, 32.74305, 32.71327, 
    32.68332, 32.65321, 32.62293, 32.59248, 32.56187, 32.53108, 32.50013, 
    32.46902, 32.43774,
  28.95008, 28.99554, 29.04087, 29.08606, 29.13111, 29.17602, 29.22079, 
    29.26542, 29.30992, 29.35427, 29.39849, 29.44256, 29.48649, 29.53028, 
    29.57393, 29.61744, 29.6608, 29.70402, 29.7471, 29.79004, 29.83283, 
    29.87548, 29.91798, 29.96034, 30.00256, 30.04462, 30.08655, 30.12833, 
    30.16996, 30.21144, 30.25278, 30.29398, 30.33502, 30.37592, 30.41667, 
    30.45727, 30.49772, 30.53802, 30.57818, 30.61818, 30.65804, 30.69774, 
    30.73729, 30.7767, 30.81595, 30.85505, 30.894, 30.93279, 30.97144, 
    31.00993, 31.04827, 31.08645, 31.12448, 31.16236, 31.20008, 31.23765, 
    31.27506, 31.31232, 31.34943, 31.38638, 31.42317, 31.4598, 31.49628, 
    31.5326, 31.56877, 31.60477, 31.64062, 31.67631, 31.71184, 31.74722, 
    31.78243, 31.81749, 31.85238, 31.88712, 31.92169, 31.9561, 31.99036, 
    32.02445, 32.05838, 32.09215, 32.12576, 32.1592, 32.19248, 32.2256, 
    32.25856, 32.29135, 32.32398, 32.35645, 32.38874, 32.42088, 32.45285, 
    32.48466, 32.5163, 32.54777, 32.57908, 32.61022, 32.6412, 32.672, 
    32.70265, 32.73312, 32.76343, 32.79356, 32.82354, 32.85334, 32.88297, 
    32.91243, 32.94173, 32.97085, 32.99981, 33.02859, 33.05721, 33.08565, 
    33.11392, 33.14202, 33.16995, 33.19771, 33.2253, 33.25271, 33.27995, 
    33.30702, 33.33392, 33.36064, 33.38719, 33.41356, 33.43976, 33.46579, 
    33.49164, 33.51732, 33.54282, 33.56815, 33.5933, 33.61828, 33.64308, 
    33.6677, 33.69215, 33.71642, 33.74051, 33.76443, 33.78817, 33.81173, 
    33.83511, 33.85832, 33.88135, 33.9042, 33.92687, 33.94936, 33.97167, 
    33.9938, 34.01575, 34.03753, 34.05912, 34.08054, 34.10177, 34.12282, 
    34.14369, 34.16438, 34.18489, 34.20522, 34.22536, 34.24532, 34.2651, 
    34.2847, 34.30412, 34.32335, 34.3424, 34.36127, 34.37996, 34.39845, 
    34.41677, 34.4349, 34.45285, 34.47062, 34.4882, 34.50559, 34.5228, 
    34.53983, 34.55667, 34.57333, 34.58979, 34.60608, 34.62218, 34.63809, 
    34.65382, 34.66936, 34.68471, 34.69988, 34.71486, 34.72965, 34.74426, 
    34.75867, 34.77291, 34.78695, 34.80081, 34.81448, 34.82796, 34.84125, 
    34.85435, 34.86727, 34.87999, 34.89253, 34.90488, 34.91705, 34.92902, 
    34.9408, 34.95239, 34.96379, 34.97501, 34.98603, 34.99687, 35.00751, 
    35.01797, 35.02823, 35.03831, 35.04819, 35.05788, 35.06739, 35.0767, 
    35.08582, 35.09475, 35.10349, 35.11204, 35.1204, 35.12856, 35.13654, 
    35.14433, 35.15192, 35.15932, 35.16653, 35.17354, 35.18037, 35.187, 
    35.19344, 35.19969, 35.20575, 35.21162, 35.21729, 35.22277, 35.22806, 
    35.23316, 35.23806, 35.24277, 35.24729, 35.25162, 35.25575, 35.25969, 
    35.26344, 35.26699, 35.27036, 35.27353, 35.2765, 35.27929, 35.28188, 
    35.28428, 35.28648, 35.2885, 35.29031, 35.29194, 35.29337, 35.29461, 
    35.29566, 35.29652, 35.29718, 35.29765, 35.29792, 35.298, 35.29789, 
    35.29758, 35.29708, 35.29639, 35.29551, 35.29443, 35.29316, 35.2917, 
    35.29004, 35.28819, 35.28615, 35.28391, 35.28148, 35.27886, 35.27605, 
    35.27304, 35.26984, 35.26645, 35.26286, 35.25908, 35.25511, 35.25095, 
    35.24659, 35.24204, 35.2373, 35.23236, 35.22724, 35.22192, 35.2164, 
    35.2107, 35.20481, 35.19872, 35.19244, 35.18597, 35.1793, 35.17245, 
    35.1654, 35.15816, 35.15073, 35.1431, 35.13529, 35.12729, 35.11909, 
    35.1107, 35.10212, 35.09335, 35.08439, 35.07524, 35.0659, 35.05636, 
    35.04664, 35.03672, 35.02662, 35.01633, 35.00584, 34.99517, 34.9843, 
    34.97325, 34.962, 34.95057, 34.93895, 34.92714, 34.91513, 34.90294, 
    34.89056, 34.87799, 34.86524, 34.85229, 34.83916, 34.82584, 34.81232, 
    34.79863, 34.78474, 34.77067, 34.75641, 34.74196, 34.72732, 34.7125, 
    34.69749, 34.68229, 34.66691, 34.65134, 34.63559, 34.61964, 34.60352, 
    34.5872, 34.5707, 34.55402, 34.53715, 34.52009, 34.50285, 34.48543, 
    34.46782, 34.45003, 34.43205, 34.41389, 34.39554, 34.37701, 34.3583, 
    34.3394, 34.32032, 34.30106, 34.28162, 34.26199, 34.24218, 34.22219, 
    34.20201, 34.18166, 34.16112, 34.1404, 34.1195, 34.09842, 34.07716, 
    34.05572, 34.0341, 34.01229, 33.99031, 33.96815, 33.94581, 33.92329, 
    33.9006, 33.87772, 33.85466, 33.83143, 33.80802, 33.78443, 33.76066, 
    33.73671, 33.71259, 33.68829, 33.66382, 33.63917, 33.61434, 33.58933, 
    33.56416, 33.5388, 33.51327, 33.48756, 33.46169, 33.43563, 33.4094, 
    33.383, 33.35642, 33.32967, 33.30275, 33.27565, 33.24839, 33.22094, 
    33.19333, 33.16555, 33.13759, 33.10946, 33.08116, 33.05269, 33.02405, 
    32.99524, 32.96626, 32.9371, 32.90778, 32.87829, 32.84863, 32.81881, 
    32.78881, 32.75864, 32.72831, 32.69781, 32.66714, 32.63631, 32.6053, 
    32.57414, 32.5428,
  29.0494, 29.09494, 29.14033, 29.18559, 29.23071, 29.27569, 29.32053, 
    29.36523, 29.40979, 29.45421, 29.49849, 29.54263, 29.58663, 29.63048, 
    29.6742, 29.71777, 29.7612, 29.80449, 29.84764, 29.89064, 29.93349, 
    29.97621, 30.01878, 30.0612, 30.10348, 30.14562, 30.18761, 30.22945, 
    30.27115, 30.3127, 30.3541, 30.39536, 30.43647, 30.47743, 30.51824, 
    30.5589, 30.59942, 30.63979, 30.68, 30.72007, 30.75999, 30.79976, 
    30.83937, 30.87884, 30.91815, 30.95732, 30.99633, 31.03518, 31.07389, 
    31.11244, 31.15084, 31.18909, 31.22718, 31.26512, 31.30291, 31.34054, 
    31.37801, 31.41533, 31.45249, 31.4895, 31.52635, 31.56305, 31.59959, 
    31.63597, 31.67219, 31.70826, 31.74416, 31.77991, 31.8155, 31.85093, 
    31.88621, 31.92132, 31.95627, 31.99107, 32.0257, 32.06017, 32.09448, 
    32.12863, 32.16262, 32.19644, 32.23011, 32.26361, 32.29694, 32.33012, 
    32.36313, 32.39598, 32.42866, 32.46118, 32.49354, 32.52573, 32.55775, 
    32.58961, 32.6213, 32.65283, 32.6842, 32.71539, 32.74642, 32.77728, 
    32.80797, 32.8385, 32.86886, 32.89905, 32.92907, 32.95892, 32.98861, 
    33.01812, 33.04746, 33.07664, 33.10564, 33.13448, 33.16314, 33.19164, 
    33.21996, 33.24811, 33.27608, 33.30389, 33.33153, 33.35899, 33.38628, 
    33.41339, 33.44033, 33.46711, 33.4937, 33.52012, 33.54637, 33.57244, 
    33.59834, 33.62406, 33.64961, 33.67498, 33.70018, 33.7252, 33.75004, 
    33.77471, 33.7992, 33.82352, 33.84765, 33.87161, 33.89539, 33.919, 
    33.94242, 33.96567, 33.98874, 34.01163, 34.03434, 34.05687, 34.07922, 
    34.1014, 34.12339, 34.1452, 34.16683, 34.18829, 34.20956, 34.23064, 
    34.25155, 34.27228, 34.29283, 34.31319, 34.33337, 34.35337, 34.37319, 
    34.39282, 34.41227, 34.43154, 34.45063, 34.46953, 34.48825, 34.50678, 
    34.52513, 34.5433, 34.56128, 34.57907, 34.59669, 34.61412, 34.63136, 
    34.64841, 34.66529, 34.68197, 34.69847, 34.71479, 34.73092, 34.74686, 
    34.76261, 34.77818, 34.79356, 34.80876, 34.82376, 34.83859, 34.85322, 
    34.86766, 34.88192, 34.89599, 34.90987, 34.92357, 34.93708, 34.95039, 
    34.96352, 34.97646, 34.98921, 35.00177, 35.01414, 35.02633, 35.03832, 
    35.05013, 35.06174, 35.07317, 35.0844, 35.09545, 35.1063, 35.11697, 
    35.12744, 35.13773, 35.14782, 35.15772, 35.16743, 35.17695, 35.18628, 
    35.19542, 35.20437, 35.21312, 35.22169, 35.23006, 35.23824, 35.24623, 
    35.25403, 35.26164, 35.26905, 35.27628, 35.28331, 35.29015, 35.29679, 
    35.30325, 35.30951, 35.31558, 35.32145, 35.32714, 35.33263, 35.33793, 
    35.34303, 35.34795, 35.35267, 35.35719, 35.36153, 35.36567, 35.36962, 
    35.37337, 35.37694, 35.38031, 35.38348, 35.38646, 35.38926, 35.39185, 
    35.39425, 35.39646, 35.39848, 35.4003, 35.40193, 35.40337, 35.40461, 
    35.40566, 35.40651, 35.40717, 35.40764, 35.40792, 35.408, 35.40789, 
    35.40758, 35.40708, 35.40639, 35.40551, 35.40443, 35.40315, 35.40168, 
    35.40002, 35.39817, 35.39613, 35.39389, 35.39145, 35.38882, 35.38601, 
    35.38299, 35.37979, 35.37638, 35.3728, 35.36901, 35.36503, 35.36086, 
    35.35649, 35.35193, 35.34718, 35.34224, 35.3371, 35.33177, 35.32625, 
    35.32054, 35.31463, 35.30853, 35.30224, 35.29575, 35.28908, 35.28221, 
    35.27515, 35.26789, 35.26045, 35.25281, 35.24498, 35.23697, 35.22875, 
    35.22035, 35.21175, 35.20296, 35.19399, 35.18482, 35.17546, 35.16591, 
    35.15617, 35.14623, 35.13611, 35.1258, 35.11529, 35.1046, 35.09371, 
    35.08264, 35.07137, 35.05992, 35.04827, 35.03644, 35.02441, 35.0122, 
    34.9998, 34.98721, 34.97443, 34.96146, 34.9483, 34.93495, 34.92142, 
    34.90769, 34.89378, 34.87968, 34.86539, 34.85092, 34.83625, 34.8214, 
    34.80637, 34.79114, 34.77573, 34.76013, 34.74435, 34.72838, 34.71222, 
    34.69588, 34.67935, 34.66263, 34.64573, 34.62864, 34.61137, 34.59391, 
    34.57627, 34.55845, 34.54044, 34.52224, 34.50386, 34.4853, 34.46655, 
    34.44762, 34.4285, 34.40921, 34.38973, 34.37006, 34.35022, 34.33019, 
    34.30998, 34.28959, 34.26902, 34.24826, 34.22732, 34.2062, 34.1849, 
    34.16343, 34.14176, 34.11992, 34.0979, 34.0757, 34.05332, 34.03076, 
    34.00802, 33.9851, 33.96201, 33.93873, 33.91528, 33.89164, 33.86784, 
    33.84385, 33.81968, 33.79534, 33.77082, 33.74612, 33.72125, 33.69621, 
    33.67098, 33.64558, 33.62001, 33.59425, 33.56833, 33.54223, 33.51595, 
    33.48951, 33.46288, 33.43608, 33.40911, 33.38197, 33.35466, 33.32717, 
    33.2995, 33.27167, 33.24366, 33.21549, 33.18714, 33.15862, 33.12993, 
    33.10107, 33.07204, 33.04284, 33.01346, 32.98392, 32.95421, 32.92433, 
    32.89428, 32.86407, 32.83368, 32.80313, 32.77241, 32.74152, 32.71047, 
    32.67924, 32.64786,
  29.14871, 29.19431, 29.23977, 29.2851, 29.33028, 29.37533, 29.42024, 
    29.46501, 29.50963, 29.55412, 29.59847, 29.64268, 29.68674, 29.73067, 
    29.77445, 29.81809, 29.86158, 29.90494, 29.94815, 29.99122, 30.03414, 
    30.07692, 30.11956, 30.16205, 30.20439, 30.24659, 30.28865, 30.33055, 
    30.37232, 30.41393, 30.4554, 30.49672, 30.53789, 30.57892, 30.6198, 
    30.66052, 30.70111, 30.74154, 30.78182, 30.82195, 30.86193, 30.90176, 
    30.94144, 30.98097, 31.02034, 31.05957, 31.09864, 31.13756, 31.17633, 
    31.21494, 31.25341, 31.29172, 31.32987, 31.36787, 31.40571, 31.44341, 
    31.48094, 31.51832, 31.55555, 31.59261, 31.62952, 31.66628, 31.70288, 
    31.73932, 31.7756, 31.81173, 31.84769, 31.8835, 31.91915, 31.95464, 
    31.98997, 32.02514, 32.06015, 32.095, 32.12969, 32.16422, 32.19859, 
    32.2328, 32.26684, 32.30072, 32.33444, 32.368, 32.40139, 32.43462, 
    32.46769, 32.5006, 32.53333, 32.56591, 32.59832, 32.63056, 32.66264, 
    32.69455, 32.7263, 32.75788, 32.7893, 32.82055, 32.85163, 32.88254, 
    32.91329, 32.94387, 32.97428, 33.00452, 33.03459, 33.0645, 33.09423, 
    33.12379, 33.15319, 33.18242, 33.21147, 33.24036, 33.26907, 33.29761, 
    33.32598, 33.35418, 33.38221, 33.41006, 33.43775, 33.46526, 33.4926, 
    33.51976, 33.54675, 33.57356, 33.60021, 33.62667, 33.65297, 33.67909, 
    33.70503, 33.7308, 33.75639, 33.78181, 33.80705, 33.83212, 33.857, 
    33.88171, 33.90625, 33.93061, 33.95478, 33.97879, 34.00261, 34.02626, 
    34.04972, 34.07301, 34.09612, 34.11906, 34.14181, 34.16438, 34.18677, 
    34.20898, 34.23101, 34.25287, 34.27454, 34.29603, 34.31734, 34.33847, 
    34.35941, 34.38018, 34.40076, 34.42116, 34.44138, 34.46141, 34.48127, 
    34.50094, 34.52042, 34.53973, 34.55885, 34.57778, 34.59653, 34.6151, 
    34.63349, 34.65169, 34.6697, 34.68753, 34.70518, 34.72264, 34.73991, 
    34.757, 34.7739, 34.79062, 34.80715, 34.82349, 34.83965, 34.85562, 
    34.87141, 34.887, 34.90241, 34.91764, 34.93267, 34.94752, 34.96218, 
    34.97665, 34.99094, 35.00503, 35.01894, 35.03266, 35.04619, 35.05953, 
    35.07269, 35.08565, 35.09842, 35.11101, 35.12341, 35.13561, 35.14763, 
    35.15945, 35.17109, 35.18254, 35.19379, 35.20486, 35.21573, 35.22642, 
    35.23691, 35.24722, 35.25733, 35.26725, 35.27698, 35.28652, 35.29586, 
    35.30502, 35.31398, 35.32276, 35.33134, 35.33973, 35.34792, 35.35593, 
    35.36374, 35.37136, 35.37879, 35.38603, 35.39307, 35.39993, 35.40658, 
    35.41305, 35.41932, 35.4254, 35.43129, 35.43699, 35.44249, 35.4478, 
    35.45291, 35.45783, 35.46256, 35.4671, 35.47144, 35.47559, 35.47955, 
    35.48331, 35.48688, 35.49025, 35.49343, 35.49643, 35.49922, 35.50182, 
    35.50423, 35.50644, 35.50846, 35.51029, 35.51192, 35.51336, 35.5146, 
    35.51565, 35.51651, 35.51717, 35.51764, 35.51792, 35.518, 35.51789, 
    35.51758, 35.51708, 35.51639, 35.5155, 35.51442, 35.51314, 35.51167, 
    35.51001, 35.50815, 35.5061, 35.50386, 35.50142, 35.49879, 35.49596, 
    35.49295, 35.48973, 35.48633, 35.48273, 35.47894, 35.47495, 35.47077, 
    35.46639, 35.46183, 35.45707, 35.45211, 35.44697, 35.44163, 35.4361, 
    35.43037, 35.42445, 35.41834, 35.41204, 35.40554, 35.39885, 35.39197, 
    35.3849, 35.37763, 35.37017, 35.36252, 35.35468, 35.34664, 35.33841, 
    35.32999, 35.32138, 35.31258, 35.30359, 35.2944, 35.28502, 35.27545, 
    35.26569, 35.25574, 35.2456, 35.23526, 35.22474, 35.21403, 35.20312, 
    35.19202, 35.18074, 35.16926, 35.1576, 35.14574, 35.13369, 35.12146, 
    35.10903, 35.09642, 35.08361, 35.07062, 35.05743, 35.04406, 35.0305, 
    35.01675, 35.00282, 34.98869, 34.97438, 34.95987, 34.94518, 34.93031, 
    34.91524, 34.89999, 34.88455, 34.86892, 34.85311, 34.83711, 34.82092, 
    34.80455, 34.78799, 34.77124, 34.75431, 34.73719, 34.71989, 34.7024, 
    34.68472, 34.66686, 34.64882, 34.63059, 34.61218, 34.59358, 34.5748, 
    34.55584, 34.53669, 34.51735, 34.49784, 34.47814, 34.45826, 34.43819, 
    34.41795, 34.39751, 34.3769, 34.35611, 34.33514, 34.31398, 34.29264, 
    34.27112, 34.24942, 34.22754, 34.20548, 34.18324, 34.16082, 34.13822, 
    34.11544, 34.09248, 34.06934, 34.04602, 34.02253, 33.99886, 33.975, 
    33.95097, 33.92677, 33.90238, 33.87782, 33.85308, 33.82816, 33.80307, 
    33.7778, 33.75235, 33.72673, 33.70094, 33.67497, 33.64882, 33.6225, 
    33.596, 33.56934, 33.54249, 33.51547, 33.48828, 33.46092, 33.43338, 
    33.40567, 33.37779, 33.34974, 33.32151, 33.29311, 33.26454, 33.2358, 
    33.20689, 33.17781, 33.14855, 33.11913, 33.08954, 33.05978, 33.02985, 
    32.99974, 32.96948, 32.93904, 32.90844, 32.87766, 32.84672, 32.81562, 
    32.78434, 32.7529,
  29.24799, 29.29366, 29.33919, 29.38459, 29.42984, 29.47495, 29.51993, 
    29.56477, 29.60946, 29.65402, 29.69843, 29.7427, 29.78684, 29.83083, 
    29.87468, 29.91838, 29.96194, 30.00537, 30.04864, 30.09178, 30.13477, 
    30.17761, 30.22031, 30.26287, 30.30528, 30.34755, 30.38967, 30.43164, 
    30.47347, 30.51515, 30.55668, 30.59806, 30.6393, 30.68039, 30.72133, 
    30.76213, 30.80277, 30.84326, 30.88361, 30.9238, 30.96385, 31.00374, 
    31.04348, 31.08307, 31.12251, 31.1618, 31.20094, 31.23992, 31.27875, 
    31.31743, 31.35595, 31.39432, 31.43254, 31.4706, 31.50851, 31.54626, 
    31.58385, 31.6213, 31.65858, 31.69571, 31.73268, 31.7695, 31.80615, 
    31.84265, 31.879, 31.91518, 31.95121, 31.98707, 32.02278, 32.05833, 
    32.09372, 32.12895, 32.16402, 32.19893, 32.23367, 32.26826, 32.30268, 
    32.33695, 32.37105, 32.40499, 32.43876, 32.47238, 32.50583, 32.53911, 
    32.57224, 32.60519, 32.63799, 32.67062, 32.70308, 32.73538, 32.76752, 
    32.79948, 32.83129, 32.86292, 32.89439, 32.92569, 32.95683, 32.98779, 
    33.01859, 33.04922, 33.07969, 33.10998, 33.1401, 33.17006, 33.19984, 
    33.22946, 33.25891, 33.28819, 33.31729, 33.34623, 33.37499, 33.40358, 
    33.432, 33.46025, 33.48832, 33.51623, 33.54396, 33.57152, 33.5989, 
    33.62611, 33.65315, 33.68002, 33.7067, 33.73322, 33.75956, 33.78572, 
    33.81171, 33.83752, 33.86316, 33.88863, 33.91391, 33.93902, 33.96395, 
    33.98871, 34.01329, 34.03769, 34.06191, 34.08596, 34.10982, 34.13351, 
    34.15702, 34.18035, 34.2035, 34.22647, 34.24927, 34.27188, 34.29431, 
    34.31657, 34.33864, 34.36053, 34.38224, 34.40377, 34.42511, 34.44628, 
    34.46727, 34.48807, 34.50869, 34.52913, 34.54938, 34.56945, 34.58934, 
    34.60905, 34.62857, 34.64791, 34.66706, 34.68604, 34.70482, 34.72342, 
    34.74184, 34.76007, 34.77812, 34.79598, 34.81366, 34.83115, 34.84846, 
    34.86558, 34.88251, 34.89926, 34.91582, 34.93219, 34.94838, 34.96438, 
    34.98019, 34.99582, 35.01126, 35.02651, 35.04158, 35.05645, 35.07114, 
    35.08564, 35.09995, 35.11407, 35.12801, 35.14175, 35.1553, 35.16867, 
    35.18185, 35.19484, 35.20763, 35.22025, 35.23266, 35.24489, 35.25693, 
    35.26878, 35.28044, 35.2919, 35.30318, 35.31427, 35.32516, 35.33587, 
    35.34638, 35.3567, 35.36684, 35.37677, 35.38652, 35.39608, 35.40545, 
    35.41462, 35.4236, 35.43239, 35.44099, 35.44939, 35.4576, 35.46562, 
    35.47345, 35.48109, 35.48853, 35.49578, 35.50283, 35.5097, 35.51637, 
    35.52285, 35.52914, 35.53523, 35.54113, 35.54683, 35.55235, 35.55766, 
    35.56279, 35.56772, 35.57246, 35.577, 35.58135, 35.58551, 35.58947, 
    35.59324, 35.59682, 35.6002, 35.60339, 35.60638, 35.60918, 35.61179, 
    35.6142, 35.61642, 35.61844, 35.62027, 35.62191, 35.62335, 35.6246, 
    35.62565, 35.62651, 35.62717, 35.62764, 35.62792, 35.628, 35.62789, 
    35.62758, 35.62708, 35.62638, 35.6255, 35.62441, 35.62313, 35.62166, 
    35.62, 35.61813, 35.61608, 35.61383, 35.61139, 35.60875, 35.60592, 
    35.6029, 35.59968, 35.59627, 35.59266, 35.58886, 35.58487, 35.58068, 
    35.5763, 35.57172, 35.56695, 35.56199, 35.55684, 35.55148, 35.54594, 
    35.54021, 35.53428, 35.52815, 35.52184, 35.51533, 35.50863, 35.50173, 
    35.49464, 35.48737, 35.47989, 35.47223, 35.46437, 35.45632, 35.44807, 
    35.43964, 35.43101, 35.42219, 35.41318, 35.40398, 35.39458, 35.38499, 
    35.37522, 35.36525, 35.35508, 35.34473, 35.33419, 35.32345, 35.31253, 
    35.30141, 35.2901, 35.27861, 35.26692, 35.25504, 35.24297, 35.23071, 
    35.21826, 35.20562, 35.19279, 35.17978, 35.16657, 35.15317, 35.13959, 
    35.12581, 35.11185, 35.0977, 35.08335, 35.06883, 35.05411, 35.0392, 
    35.02411, 35.00883, 34.99336, 34.97771, 34.96186, 34.94583, 34.92962, 
    34.91321, 34.89662, 34.87984, 34.86288, 34.84573, 34.8284, 34.81087, 
    34.79317, 34.77528, 34.7572, 34.73894, 34.72049, 34.70186, 34.68304, 
    34.66404, 34.64486, 34.62549, 34.60594, 34.58621, 34.56629, 34.54619, 
    34.52591, 34.50544, 34.48479, 34.46396, 34.44294, 34.42175, 34.40038, 
    34.37881, 34.35708, 34.33516, 34.31306, 34.29078, 34.26831, 34.24567, 
    34.22285, 34.19985, 34.17667, 34.15331, 34.12978, 34.10606, 34.08216, 
    34.05809, 34.03384, 34.00941, 33.98481, 33.96002, 33.93506, 33.90992, 
    33.88461, 33.85912, 33.83345, 33.80761, 33.7816, 33.7554, 33.72903, 
    33.70249, 33.67578, 33.64889, 33.62182, 33.59458, 33.56717, 33.53959, 
    33.51183, 33.48389, 33.45579, 33.42752, 33.39907, 33.37045, 33.34166, 
    33.3127, 33.28357, 33.25426, 33.22479, 33.19514, 33.16533, 33.13535, 
    33.1052, 33.07488, 33.04439, 33.01373, 32.98291, 32.95191, 32.92075, 
    32.88942, 32.85793,
  29.34726, 29.39299, 29.43859, 29.48405, 29.52938, 29.57456, 29.6196, 
    29.6645, 29.70927, 29.75389, 29.79837, 29.84271, 29.88691, 29.93097, 
    29.97488, 30.01866, 30.06229, 30.10577, 30.14912, 30.19232, 30.23537, 
    30.27828, 30.32105, 30.36367, 30.40615, 30.44848, 30.49067, 30.5327, 
    30.5746, 30.61634, 30.65794, 30.69939, 30.74069, 30.78185, 30.82285, 
    30.86371, 30.90442, 30.94497, 30.98538, 31.02564, 31.06575, 31.10571, 
    31.14551, 31.18517, 31.22467, 31.26402, 31.30322, 31.34226, 31.38116, 
    31.4199, 31.45848, 31.49691, 31.53519, 31.57331, 31.61128, 31.6491, 
    31.68675, 31.72425, 31.7616, 31.79879, 31.83582, 31.8727, 31.90941, 
    31.94597, 31.98238, 32.01862, 32.0547, 32.09063, 32.1264, 32.16201, 
    32.19745, 32.23274, 32.26787, 32.30283, 32.33764, 32.37228, 32.40676, 
    32.44109, 32.47524, 32.50924, 32.54307, 32.57674, 32.61025, 32.64359, 
    32.67677, 32.70979, 32.74263, 32.77532, 32.80784, 32.84019, 32.87238, 
    32.9044, 32.93626, 32.96795, 32.99947, 33.03083, 33.06201, 33.09303, 
    33.12389, 33.15457, 33.18508, 33.21543, 33.24561, 33.27561, 33.30545, 
    33.33512, 33.36462, 33.39394, 33.4231, 33.45208, 33.4809, 33.50954, 
    33.53801, 33.5663, 33.59443, 33.62238, 33.65016, 33.67777, 33.7052, 
    33.73246, 33.75954, 33.78646, 33.81319, 33.83975, 33.86614, 33.89235, 
    33.91838, 33.94424, 33.96993, 33.99544, 34.02077, 34.04592, 34.0709, 
    34.0957, 34.12032, 34.14476, 34.16903, 34.19312, 34.21703, 34.24076, 
    34.26431, 34.28768, 34.31087, 34.33389, 34.35672, 34.37938, 34.40185, 
    34.42414, 34.44625, 34.46818, 34.48993, 34.5115, 34.53289, 34.55409, 
    34.57511, 34.59595, 34.61661, 34.63708, 34.65738, 34.67749, 34.69741, 
    34.71715, 34.73671, 34.75608, 34.77527, 34.79428, 34.8131, 34.83174, 
    34.85019, 34.86845, 34.88654, 34.90443, 34.92214, 34.93966, 34.957, 
    34.97415, 34.99112, 35.0079, 35.02449, 35.04089, 35.05711, 35.07314, 
    35.08898, 35.10464, 35.12011, 35.13538, 35.15047, 35.16538, 35.18009, 
    35.19462, 35.20896, 35.22311, 35.23706, 35.25084, 35.26442, 35.27781, 
    35.29101, 35.30402, 35.31684, 35.32948, 35.34192, 35.35417, 35.36623, 
    35.3781, 35.38978, 35.40127, 35.41257, 35.42368, 35.43459, 35.44532, 
    35.45585, 35.46619, 35.47634, 35.4863, 35.49607, 35.50564, 35.51503, 
    35.52422, 35.53321, 35.54202, 35.55063, 35.55905, 35.56728, 35.57532, 
    35.58316, 35.59081, 35.59827, 35.60553, 35.6126, 35.61948, 35.62616, 
    35.63265, 35.63895, 35.64505, 35.65096, 35.65668, 35.6622, 35.66753, 
    35.67266, 35.6776, 35.68235, 35.6869, 35.69127, 35.69543, 35.6994, 
    35.70318, 35.70676, 35.71015, 35.71334, 35.71634, 35.71915, 35.72176, 
    35.72417, 35.72639, 35.72842, 35.73026, 35.7319, 35.73334, 35.73459, 
    35.73565, 35.7365, 35.73717, 35.73764, 35.73792, 35.738, 35.73789, 
    35.73758, 35.73708, 35.73638, 35.73549, 35.73441, 35.73312, 35.73165, 
    35.72998, 35.72812, 35.72606, 35.7238, 35.72136, 35.71872, 35.71588, 
    35.71285, 35.70963, 35.70621, 35.70259, 35.69878, 35.69478, 35.69059, 
    35.6862, 35.68161, 35.67684, 35.67186, 35.6667, 35.66134, 35.65578, 
    35.65004, 35.6441, 35.63797, 35.63164, 35.62511, 35.6184, 35.61149, 
    35.60439, 35.5971, 35.58961, 35.58193, 35.57406, 35.56599, 35.55774, 
    35.54928, 35.54064, 35.5318, 35.52277, 35.51355, 35.50414, 35.49453, 
    35.48474, 35.47475, 35.46457, 35.4542, 35.44363, 35.43288, 35.42193, 
    35.41079, 35.39947, 35.38795, 35.37624, 35.36433, 35.35225, 35.33996, 
    35.32749, 35.31483, 35.30198, 35.28893, 35.2757, 35.26228, 35.24867, 
    35.23487, 35.22088, 35.2067, 35.19233, 35.17778, 35.16303, 35.1481, 
    35.13298, 35.11767, 35.10217, 35.08649, 35.07062, 35.05456, 35.03831, 
    35.02187, 35.00525, 34.98845, 34.97145, 34.95427, 34.9369, 34.91935, 
    34.90161, 34.88369, 34.86558, 34.84728, 34.8288, 34.81013, 34.79129, 
    34.77225, 34.75303, 34.73363, 34.71404, 34.69427, 34.67432, 34.65418, 
    34.63386, 34.61335, 34.59267, 34.5718, 34.55075, 34.52951, 34.5081, 
    34.4865, 34.46473, 34.44276, 34.42062, 34.3983, 34.3758, 34.35312, 
    34.33026, 34.30722, 34.284, 34.26059, 34.23701, 34.21326, 34.18932, 
    34.1652, 34.14091, 34.11644, 34.09179, 34.06696, 34.04195, 34.01677, 
    33.99141, 33.96588, 33.94017, 33.91428, 33.88821, 33.86198, 33.83556, 
    33.80898, 33.78221, 33.75527, 33.72816, 33.70087, 33.67341, 33.64578, 
    33.61797, 33.58999, 33.56184, 33.53352, 33.50502, 33.47635, 33.44751, 
    33.4185, 33.38931, 33.35996, 33.33044, 33.30074, 33.27088, 33.24084, 
    33.21064, 33.18027, 33.14973, 33.11901, 33.08814, 33.05709, 33.02588, 
    32.9945, 32.96295,
  29.4465, 29.4923, 29.53797, 29.5835, 29.62889, 29.67414, 29.71925, 
    29.76422, 29.80905, 29.85374, 29.89829, 29.9427, 29.98696, 30.03109, 
    30.07507, 30.11891, 30.16261, 30.20616, 30.24957, 30.29284, 30.33596, 
    30.37893, 30.42177, 30.46446, 30.507, 30.5494, 30.59165, 30.63375, 
    30.67571, 30.71752, 30.75918, 30.8007, 30.84206, 30.88328, 30.92435, 
    30.96527, 31.00605, 31.04667, 31.08714, 31.12746, 31.16763, 31.20765, 
    31.24752, 31.28724, 31.32681, 31.36622, 31.40548, 31.44459, 31.48354, 
    31.52235, 31.56099, 31.59949, 31.63783, 31.67601, 31.71404, 31.75191, 
    31.78963, 31.8272, 31.8646, 31.90185, 31.93894, 31.97588, 32.01266, 
    32.04928, 32.08574, 32.12204, 32.15819, 32.19417, 32.23, 32.26567, 
    32.30117, 32.33652, 32.3717, 32.40673, 32.44159, 32.47629, 32.51083, 
    32.54521, 32.57943, 32.61348, 32.64737, 32.6811, 32.71466, 32.74805, 
    32.78129, 32.81436, 32.84727, 32.88, 32.91258, 32.94499, 32.97723, 
    33.00931, 33.04122, 33.07296, 33.10454, 33.13595, 33.16719, 33.19826, 
    33.22916, 33.2599, 33.29047, 33.32087, 33.3511, 33.38115, 33.41105, 
    33.44076, 33.47031, 33.49969, 33.5289, 33.55793, 33.58679, 33.61549, 
    33.644, 33.67235, 33.70053, 33.72853, 33.75636, 33.78401, 33.81149, 
    33.8388, 33.86593, 33.89289, 33.91967, 33.94628, 33.97271, 33.99897, 
    34.02505, 34.05096, 34.07668, 34.10224, 34.12761, 34.15281, 34.17783, 
    34.20267, 34.22734, 34.25183, 34.27614, 34.30027, 34.32422, 34.348, 
    34.37159, 34.395, 34.41824, 34.44129, 34.46417, 34.48686, 34.50938, 
    34.53171, 34.55386, 34.57583, 34.59762, 34.61922, 34.64065, 34.66189, 
    34.68295, 34.70383, 34.72453, 34.74504, 34.76537, 34.78551, 34.80547, 
    34.82525, 34.84484, 34.86425, 34.88348, 34.90252, 34.92138, 34.94004, 
    34.95853, 34.97683, 34.99495, 35.01287, 35.03061, 35.04817, 35.06554, 
    35.08272, 35.09972, 35.11653, 35.13315, 35.14959, 35.16583, 35.18189, 
    35.19777, 35.21345, 35.22895, 35.24426, 35.25937, 35.2743, 35.28905, 
    35.3036, 35.31796, 35.33214, 35.34612, 35.35992, 35.37352, 35.38694, 
    35.40017, 35.4132, 35.42605, 35.43871, 35.45117, 35.46345, 35.47553, 
    35.48742, 35.49913, 35.51064, 35.52195, 35.53308, 35.54402, 35.55476, 
    35.56532, 35.57568, 35.58585, 35.59583, 35.60561, 35.6152, 35.6246, 
    35.63381, 35.64283, 35.65165, 35.66028, 35.66871, 35.67696, 35.68501, 
    35.69287, 35.70053, 35.708, 35.71528, 35.72236, 35.72925, 35.73595, 
    35.74245, 35.74876, 35.75488, 35.7608, 35.76653, 35.77206, 35.7774, 
    35.78254, 35.78749, 35.79225, 35.79681, 35.80117, 35.80535, 35.80933, 
    35.81311, 35.8167, 35.8201, 35.8233, 35.8263, 35.82911, 35.83173, 
    35.83415, 35.83638, 35.83841, 35.84024, 35.84188, 35.84333, 35.84458, 
    35.84564, 35.8465, 35.84717, 35.84764, 35.84792, 35.848, 35.84789, 
    35.84758, 35.84708, 35.84638, 35.84549, 35.8444, 35.84312, 35.84164, 
    35.83997, 35.8381, 35.83604, 35.83378, 35.83133, 35.82868, 35.82584, 
    35.8228, 35.81957, 35.81615, 35.81253, 35.80871, 35.8047, 35.8005, 
    35.7961, 35.79151, 35.78672, 35.78174, 35.77657, 35.77119, 35.76563, 
    35.75987, 35.75392, 35.74778, 35.74144, 35.7349, 35.72818, 35.72125, 
    35.71414, 35.70683, 35.69933, 35.69164, 35.68375, 35.67567, 35.66739, 
    35.65892, 35.65026, 35.64141, 35.63237, 35.62313, 35.6137, 35.60408, 
    35.59426, 35.58425, 35.57405, 35.56366, 35.55308, 35.5423, 35.53133, 
    35.52018, 35.50883, 35.49729, 35.48555, 35.47363, 35.46152, 35.44921, 
    35.43672, 35.42403, 35.41116, 35.39809, 35.38483, 35.37138, 35.35775, 
    35.34392, 35.32991, 35.3157, 35.30131, 35.28673, 35.27195, 35.25699, 
    35.24184, 35.22651, 35.21098, 35.19527, 35.17936, 35.16328, 35.147, 
    35.13054, 35.11388, 35.09704, 35.08002, 35.06281, 35.04541, 35.02782, 
    35.01005, 34.99209, 34.97395, 34.95562, 34.9371, 34.9184, 34.89952, 
    34.88045, 34.86119, 34.84176, 34.82214, 34.80233, 34.78234, 34.76217, 
    34.74181, 34.72126, 34.70054, 34.67963, 34.65855, 34.63727, 34.61582, 
    34.59418, 34.57236, 34.55037, 34.52819, 34.50583, 34.48328, 34.46056, 
    34.43766, 34.41457, 34.39131, 34.36787, 34.34425, 34.32045, 34.29646, 
    34.2723, 34.24797, 34.22345, 34.19876, 34.17389, 34.14884, 34.12361, 
    34.09821, 34.07263, 34.04687, 34.02094, 33.99483, 33.96854, 33.94208, 
    33.91545, 33.88863, 33.86165, 33.83449, 33.80716, 33.77965, 33.75196, 
    33.72411, 33.69608, 33.66788, 33.6395, 33.61096, 33.58224, 33.55335, 
    33.52428, 33.49505, 33.46565, 33.43607, 33.40633, 33.37641, 33.34632, 
    33.31607, 33.28564, 33.25505, 33.22429, 33.19336, 33.16226, 33.13099, 
    33.09956, 33.06795,
  29.54572, 29.59159, 29.63733, 29.68292, 29.72838, 29.7737, 29.81887, 
    29.86391, 29.90881, 29.95357, 29.99819, 30.04266, 30.08699, 30.13119, 
    30.17523, 30.21914, 30.26291, 30.30653, 30.35, 30.39334, 30.43652, 
    30.47957, 30.52247, 30.56522, 30.60783, 30.65029, 30.69261, 30.73478, 
    30.7768, 30.81867, 30.8604, 30.90198, 30.94341, 30.9847, 31.02583, 
    31.06682, 31.10765, 31.14834, 31.18888, 31.22926, 31.2695, 31.30958, 
    31.34952, 31.3893, 31.42892, 31.4684, 31.50773, 31.5469, 31.58591, 
    31.62478, 31.66349, 31.70204, 31.74045, 31.77869, 31.81678, 31.85472, 
    31.8925, 31.93012, 31.96759, 32.0049, 32.04205, 32.07905, 32.11589, 
    32.15257, 32.18909, 32.22545, 32.26165, 32.2977, 32.33358, 32.36931, 
    32.40488, 32.44028, 32.47552, 32.51061, 32.54553, 32.58029, 32.61489, 
    32.64932, 32.68359, 32.7177, 32.75165, 32.78543, 32.81905, 32.8525, 
    32.8858, 32.91892, 32.95189, 32.98468, 33.01731, 33.04977, 33.08207, 
    33.1142, 33.14617, 33.17796, 33.20959, 33.24105, 33.27235, 33.30348, 
    33.33443, 33.36522, 33.39584, 33.42629, 33.45657, 33.48669, 33.51662, 
    33.5464, 33.576, 33.60542, 33.63468, 33.66377, 33.69268, 33.72142, 
    33.74999, 33.77839, 33.80661, 33.83466, 33.86254, 33.89024, 33.91777, 
    33.94513, 33.97231, 33.99931, 34.02614, 34.0528, 34.07928, 34.10558, 
    34.13171, 34.15766, 34.18343, 34.20903, 34.23445, 34.25969, 34.28476, 
    34.30965, 34.33436, 34.35889, 34.38324, 34.40742, 34.43141, 34.45523, 
    34.47886, 34.50232, 34.5256, 34.54869, 34.57161, 34.59434, 34.6169, 
    34.63927, 34.66146, 34.68347, 34.7053, 34.72694, 34.74841, 34.76969, 
    34.79079, 34.81171, 34.83244, 34.85299, 34.87335, 34.89354, 34.91353, 
    34.93335, 34.95298, 34.97242, 34.99168, 35.01076, 35.02964, 35.04835, 
    35.06687, 35.0852, 35.10335, 35.12131, 35.13908, 35.15667, 35.17408, 
    35.19129, 35.20832, 35.22516, 35.24181, 35.25828, 35.27456, 35.29064, 
    35.30655, 35.32226, 35.33778, 35.35312, 35.36827, 35.38322, 35.39799, 
    35.41257, 35.42697, 35.44117, 35.45518, 35.469, 35.48263, 35.49607, 
    35.50932, 35.52238, 35.53526, 35.54794, 35.56042, 35.57272, 35.58483, 
    35.59674, 35.60847, 35.62, 35.63134, 35.64249, 35.65345, 35.66421, 
    35.67478, 35.68517, 35.69535, 35.70535, 35.71515, 35.72476, 35.73418, 
    35.7434, 35.75244, 35.76128, 35.76992, 35.77837, 35.78663, 35.7947, 
    35.80257, 35.81025, 35.81773, 35.82503, 35.83212, 35.83903, 35.84574, 
    35.85225, 35.85857, 35.8647, 35.87063, 35.87637, 35.88191, 35.88726, 
    35.89241, 35.89738, 35.90214, 35.90671, 35.91109, 35.91527, 35.91925, 
    35.92305, 35.92664, 35.93004, 35.93325, 35.93626, 35.93908, 35.9417, 
    35.94412, 35.94635, 35.94839, 35.95023, 35.95187, 35.95332, 35.95457, 
    35.95564, 35.9565, 35.95717, 35.95764, 35.95792, 35.958, 35.95789, 
    35.95758, 35.95707, 35.95638, 35.95548, 35.95439, 35.95311, 35.95163, 
    35.94995, 35.94808, 35.94601, 35.94375, 35.9413, 35.93864, 35.93579, 
    35.93275, 35.92952, 35.92609, 35.92246, 35.91864, 35.91462, 35.91041, 
    35.906, 35.9014, 35.8966, 35.89161, 35.88643, 35.88105, 35.87547, 
    35.86971, 35.86374, 35.85759, 35.85123, 35.84469, 35.83795, 35.83101, 
    35.82389, 35.81656, 35.80905, 35.80134, 35.79344, 35.78534, 35.77705, 
    35.76857, 35.75989, 35.75102, 35.74196, 35.7327, 35.72326, 35.71362, 
    35.70378, 35.69375, 35.68354, 35.67312, 35.66252, 35.65173, 35.64074, 
    35.62956, 35.61819, 35.60662, 35.59487, 35.58292, 35.57079, 35.55846, 
    35.54594, 35.53323, 35.52033, 35.50724, 35.49396, 35.48049, 35.46683, 
    35.45298, 35.43893, 35.4247, 35.41028, 35.39567, 35.38087, 35.36588, 
    35.3507, 35.33534, 35.31979, 35.30404, 35.28811, 35.27199, 35.25568, 
    35.23919, 35.22251, 35.20564, 35.18858, 35.17133, 35.1539, 35.13629, 
    35.11848, 35.10049, 35.08231, 35.06395, 35.0454, 35.02667, 35.00775, 
    34.98865, 34.96936, 34.94988, 34.93023, 34.91038, 34.89035, 34.87014, 
    34.84975, 34.82917, 34.80841, 34.78746, 34.76633, 34.74503, 34.72353, 
    34.70186, 34.68, 34.65796, 34.63574, 34.61334, 34.59076, 34.56799, 
    34.54505, 34.52193, 34.49862, 34.47514, 34.45147, 34.42763, 34.4036, 
    34.3794, 34.35502, 34.33046, 34.30572, 34.28081, 34.25571, 34.23044, 
    34.20499, 34.17937, 34.15356, 34.12759, 34.10143, 34.0751, 34.04859, 
    34.02191, 33.99505, 33.96802, 33.94081, 33.91343, 33.88587, 33.85814, 
    33.83023, 33.80216, 33.77391, 33.74548, 33.71689, 33.68812, 33.65918, 
    33.63007, 33.60078, 33.57132, 33.5417, 33.5119, 33.48193, 33.4518, 
    33.42149, 33.39101, 33.36036, 33.32955, 33.29856, 33.26741, 33.23609, 
    33.2046, 33.17295,
  29.64491, 29.69086, 29.73666, 29.78232, 29.82785, 29.87323, 29.91848, 
    29.96359, 30.00855, 30.05338, 30.09806, 30.1426, 30.187, 30.23126, 
    30.27538, 30.31935, 30.36318, 30.40687, 30.45041, 30.49381, 30.53707, 
    30.58018, 30.62314, 30.66596, 30.70864, 30.75117, 30.79355, 30.83578, 
    30.87787, 30.91981, 30.96161, 31.00325, 31.04475, 31.0861, 31.1273, 
    31.16835, 31.20925, 31.25, 31.2906, 31.33105, 31.37135, 31.41149, 
    31.45149, 31.49133, 31.53103, 31.57057, 31.60995, 31.64919, 31.68827, 
    31.72719, 31.76597, 31.80458, 31.84305, 31.88136, 31.91951, 31.95751, 
    31.99535, 32.03303, 32.07056, 32.10793, 32.14515, 32.1822, 32.2191, 
    32.25584, 32.29242, 32.32885, 32.36511, 32.40121, 32.43716, 32.47294, 
    32.50856, 32.54403, 32.57933, 32.61447, 32.64945, 32.68427, 32.71893, 
    32.75342, 32.78775, 32.82191, 32.85592, 32.88976, 32.92343, 32.95694, 
    32.99029, 33.02347, 33.05649, 33.08934, 33.12202, 33.15454, 33.1869, 
    33.21908, 33.2511, 33.28296, 33.31464, 33.34615, 33.3775, 33.40868, 
    33.43969, 33.47054, 33.50121, 33.53171, 33.56204, 33.59221, 33.6222, 
    33.65202, 33.68167, 33.71115, 33.74046, 33.76959, 33.79856, 33.82735, 
    33.85597, 33.88441, 33.91269, 33.94078, 33.96871, 33.99646, 34.02404, 
    34.05145, 34.07867, 34.10572, 34.1326, 34.15931, 34.18583, 34.21218, 
    34.23835, 34.26435, 34.29017, 34.31581, 34.34128, 34.36657, 34.39168, 
    34.41661, 34.44136, 34.46594, 34.49034, 34.51455, 34.53859, 34.56245, 
    34.58613, 34.60963, 34.63295, 34.65609, 34.67904, 34.70182, 34.72441, 
    34.74683, 34.76906, 34.79111, 34.81297, 34.83466, 34.85616, 34.87748, 
    34.89862, 34.91957, 34.94034, 34.96093, 34.98133, 35.00155, 35.02159, 
    35.04144, 35.0611, 35.08058, 35.09988, 35.11899, 35.13791, 35.15665, 
    35.1752, 35.19357, 35.21175, 35.22974, 35.24755, 35.26517, 35.28261, 
    35.29985, 35.31691, 35.33378, 35.35047, 35.36696, 35.38327, 35.39939, 
    35.41532, 35.43106, 35.44662, 35.46198, 35.47716, 35.49215, 35.50694, 
    35.52155, 35.53596, 35.55019, 35.56423, 35.57808, 35.59174, 35.6052, 
    35.61848, 35.63157, 35.64446, 35.65716, 35.66967, 35.682, 35.69412, 
    35.70606, 35.71781, 35.72936, 35.74072, 35.75189, 35.76287, 35.77365, 
    35.78425, 35.79465, 35.80486, 35.81487, 35.82469, 35.83432, 35.84376, 
    35.853, 35.86205, 35.8709, 35.87957, 35.88803, 35.89631, 35.90439, 
    35.91228, 35.91997, 35.92747, 35.93477, 35.94188, 35.9488, 35.95552, 
    35.96205, 35.96838, 35.97452, 35.98046, 35.98621, 35.99177, 35.99713, 
    36.00229, 36.00726, 36.01204, 36.01661, 36.021, 36.02519, 36.02918, 
    36.03298, 36.03658, 36.03999, 36.0432, 36.04622, 36.04904, 36.05167, 
    36.0541, 36.05633, 36.05837, 36.06021, 36.06186, 36.06331, 36.06457, 
    36.06563, 36.06649, 36.06717, 36.06764, 36.06792, 36.068, 36.06789, 
    36.06758, 36.06707, 36.06637, 36.06548, 36.06438, 36.0631, 36.06161, 
    36.05993, 36.05806, 36.05599, 36.05372, 36.05126, 36.04861, 36.04575, 
    36.04271, 36.03946, 36.03603, 36.03239, 36.02856, 36.02454, 36.02032, 
    36.0159, 36.01129, 36.00649, 36.00149, 35.99629, 35.9909, 35.98532, 
    35.97954, 35.97356, 35.9674, 35.96103, 35.95447, 35.94772, 35.94077, 
    35.93363, 35.9263, 35.91877, 35.91104, 35.90313, 35.89501, 35.88671, 
    35.87821, 35.86951, 35.86063, 35.85155, 35.84228, 35.83281, 35.82315, 
    35.8133, 35.80325, 35.79301, 35.78259, 35.77196, 35.76115, 35.75014, 
    35.73894, 35.72755, 35.71596, 35.70419, 35.69222, 35.68006, 35.66771, 
    35.65516, 35.64243, 35.62951, 35.61639, 35.60308, 35.58959, 35.5759, 
    35.56202, 35.54795, 35.5337, 35.51925, 35.50461, 35.48979, 35.47477, 
    35.45956, 35.44417, 35.42859, 35.41282, 35.39685, 35.3807, 35.36436, 
    35.34784, 35.33113, 35.31423, 35.29714, 35.27986, 35.2624, 35.24475, 
    35.22691, 35.20889, 35.19068, 35.17228, 35.1537, 35.13493, 35.11598, 
    35.09684, 35.07751, 35.058, 35.03831, 35.01843, 34.99837, 34.97812, 
    34.95769, 34.93707, 34.91627, 34.89529, 34.87412, 34.85277, 34.83124, 
    34.80953, 34.78763, 34.76555, 34.74329, 34.72085, 34.69823, 34.67542, 
    34.65244, 34.62927, 34.60592, 34.5824, 34.55869, 34.5348, 34.51073, 
    34.48649, 34.46207, 34.43746, 34.41268, 34.38772, 34.36258, 34.33727, 
    34.31177, 34.2861, 34.26025, 34.23423, 34.20802, 34.18165, 34.15509, 
    34.12836, 34.10146, 34.07438, 34.04712, 34.01969, 33.99208, 33.96431, 
    33.93635, 33.90823, 33.87992, 33.85145, 33.82281, 33.79399, 33.765, 
    33.73583, 33.7065, 33.67699, 33.64731, 33.61747, 33.58744, 33.55725, 
    33.52689, 33.49636, 33.46567, 33.4348, 33.40376, 33.37255, 33.34118, 
    33.30964, 33.27793,
  29.74409, 29.7901, 29.83597, 29.8817, 29.9273, 29.97275, 30.01806, 
    30.06324, 30.10827, 30.15316, 30.19792, 30.24253, 30.28699, 30.33132, 
    30.3755, 30.41954, 30.46344, 30.50719, 30.55081, 30.59427, 30.63759, 
    30.68077, 30.7238, 30.76669, 30.80943, 30.85202, 30.89447, 30.93677, 
    30.97892, 31.02093, 31.06279, 31.1045, 31.14606, 31.18748, 31.22874, 
    31.26985, 31.31082, 31.35163, 31.3923, 31.43281, 31.47318, 31.51339, 
    31.55345, 31.59336, 31.63311, 31.67271, 31.71216, 31.75146, 31.7906, 
    31.82959, 31.86843, 31.90711, 31.94563, 31.984, 32.02222, 32.06028, 
    32.09818, 32.13593, 32.17351, 32.21095, 32.24822, 32.28534, 32.3223, 
    32.3591, 32.39574, 32.43222, 32.46854, 32.50471, 32.54071, 32.57656, 
    32.61224, 32.64776, 32.68312, 32.71832, 32.75336, 32.78823, 32.82295, 
    32.8575, 32.89189, 32.92611, 32.96017, 32.99407, 33.0278, 33.06137, 
    33.09477, 33.12801, 33.16108, 33.19399, 33.22673, 33.2593, 33.29171, 
    33.32395, 33.35603, 33.38793, 33.41967, 33.45124, 33.48264, 33.51387, 
    33.54494, 33.57583, 33.60656, 33.63711, 33.6675, 33.69771, 33.72776, 
    33.75763, 33.78733, 33.81686, 33.84622, 33.87541, 33.90442, 33.93327, 
    33.96193, 33.99043, 34.01875, 34.0469, 34.07487, 34.10268, 34.1303, 
    34.15775, 34.18503, 34.21213, 34.23906, 34.2658, 34.29238, 34.31878, 
    34.34499, 34.37104, 34.3969, 34.42259, 34.4481, 34.47343, 34.49859, 
    34.52357, 34.54837, 34.57299, 34.59742, 34.62169, 34.64577, 34.66967, 
    34.69339, 34.71693, 34.74029, 34.76347, 34.78647, 34.80928, 34.83192, 
    34.85437, 34.87665, 34.89874, 34.92064, 34.94237, 34.96391, 34.98527, 
    35.00644, 35.02744, 35.04824, 35.06887, 35.08931, 35.10956, 35.12963, 
    35.14952, 35.16922, 35.18874, 35.20807, 35.22721, 35.24617, 35.26495, 
    35.28354, 35.30193, 35.32015, 35.33818, 35.35601, 35.37367, 35.39114, 
    35.40841, 35.4255, 35.44241, 35.45912, 35.47565, 35.49199, 35.50813, 
    35.52409, 35.53987, 35.55545, 35.57084, 35.58604, 35.60106, 35.61588, 
    35.63052, 35.64496, 35.65922, 35.67328, 35.68716, 35.70084, 35.71433, 
    35.72763, 35.74074, 35.75366, 35.76638, 35.77892, 35.79126, 35.80342, 
    35.81538, 35.82714, 35.83872, 35.8501, 35.86129, 35.87229, 35.8831, 
    35.89371, 35.90413, 35.91436, 35.92439, 35.93423, 35.94388, 35.95333, 
    35.96259, 35.97166, 35.98053, 35.98921, 35.99769, 36.00598, 36.01408, 
    36.02198, 36.02969, 36.0372, 36.04452, 36.05164, 36.05857, 36.06531, 
    36.07185, 36.07819, 36.08434, 36.0903, 36.09606, 36.10162, 36.10699, 
    36.11217, 36.11715, 36.12193, 36.12651, 36.13091, 36.13511, 36.13911, 
    36.14291, 36.14652, 36.14994, 36.15315, 36.15618, 36.159, 36.16163, 
    36.16407, 36.16631, 36.16835, 36.1702, 36.17185, 36.17331, 36.17456, 
    36.17562, 36.17649, 36.17716, 36.17764, 36.17792, 36.178, 36.17789, 
    36.17758, 36.17707, 36.17637, 36.17547, 36.17438, 36.17309, 36.1716, 
    36.16992, 36.16804, 36.16597, 36.1637, 36.16123, 36.15857, 36.15571, 
    36.15266, 36.14941, 36.14597, 36.14232, 36.13848, 36.13445, 36.13023, 
    36.1258, 36.12119, 36.11637, 36.11136, 36.10616, 36.10075, 36.09516, 
    36.08937, 36.08339, 36.0772, 36.07083, 36.06426, 36.05749, 36.05053, 
    36.04338, 36.03603, 36.02848, 36.02074, 36.01281, 36.00468, 35.99636, 
    35.98785, 35.97914, 35.97024, 35.96114, 35.95185, 35.94236, 35.93269, 
    35.92282, 35.91275, 35.9025, 35.89204, 35.8814, 35.87056, 35.85954, 
    35.84832, 35.8369, 35.82529, 35.8135, 35.80151, 35.78933, 35.77695, 
    35.76439, 35.75163, 35.73868, 35.72554, 35.71221, 35.69868, 35.68497, 
    35.67107, 35.65697, 35.64269, 35.62822, 35.61355, 35.5987, 35.58365, 
    35.56842, 35.553, 35.53738, 35.52158, 35.50559, 35.48941, 35.47305, 
    35.45649, 35.43974, 35.42281, 35.40569, 35.38839, 35.37089, 35.35321, 
    35.33533, 35.31728, 35.29903, 35.28061, 35.26199, 35.24319, 35.2242, 
    35.20502, 35.18566, 35.16612, 35.14639, 35.12647, 35.10637, 35.08609, 
    35.06562, 35.04496, 35.02413, 35.00311, 34.9819, 34.96051, 34.93894, 
    34.91719, 34.89525, 34.87313, 34.85083, 34.82835, 34.80569, 34.78284, 
    34.75982, 34.73661, 34.71322, 34.68965, 34.6659, 34.64197, 34.61786, 
    34.59357, 34.5691, 34.54446, 34.51963, 34.49463, 34.46944, 34.44408, 
    34.41854, 34.39282, 34.36693, 34.34086, 34.31461, 34.28819, 34.26159, 
    34.23481, 34.20786, 34.18073, 34.15342, 34.12594, 34.09829, 34.07046, 
    34.04246, 34.01429, 33.98594, 33.95741, 33.92871, 33.89985, 33.8708, 
    33.84159, 33.8122, 33.78265, 33.75292, 33.72302, 33.69295, 33.6627, 
    33.63229, 33.60171, 33.57096, 33.54004, 33.50895, 33.47768, 33.44625, 
    33.41466, 33.3829,
  29.84324, 29.88932, 29.93526, 29.98106, 30.02672, 30.07224, 30.11762, 
    30.16287, 30.20797, 30.25293, 30.29775, 30.34243, 30.38696, 30.43135, 
    30.47561, 30.51971, 30.56368, 30.6075, 30.65118, 30.69471, 30.7381, 
    30.78134, 30.82444, 30.86739, 30.9102, 30.95286, 30.99537, 31.03774, 
    31.07996, 31.12203, 31.16395, 31.20573, 31.24735, 31.28883, 31.33016, 
    31.37134, 31.41237, 31.45325, 31.49398, 31.53456, 31.57499, 31.61526, 
    31.65538, 31.69536, 31.73517, 31.77484, 31.81435, 31.85371, 31.89292, 
    31.93197, 31.97087, 32.00961, 32.0482, 32.08663, 32.12491, 32.16303, 
    32.20099, 32.2388, 32.27645, 32.31395, 32.35128, 32.38846, 32.42548, 
    32.46234, 32.49904, 32.53558, 32.57197, 32.60819, 32.64425, 32.68016, 
    32.7159, 32.75148, 32.7869, 32.82216, 32.85725, 32.89219, 32.92696, 
    32.96157, 32.99601, 33.03029, 33.06441, 33.09837, 33.13215, 33.16578, 
    33.19924, 33.23253, 33.26566, 33.29862, 33.33142, 33.36405, 33.39651, 
    33.42881, 33.46093, 33.4929, 33.52469, 33.55631, 33.58777, 33.61905, 
    33.65017, 33.68112, 33.7119, 33.7425, 33.77295, 33.80321, 33.83331, 
    33.86323, 33.89299, 33.92257, 33.95198, 33.98122, 34.01028, 34.03917, 
    34.06789, 34.09644, 34.12481, 34.15301, 34.18103, 34.20888, 34.23655, 
    34.26405, 34.29138, 34.31852, 34.3455, 34.3723, 34.39891, 34.42536, 
    34.45163, 34.47771, 34.50362, 34.52936, 34.55492, 34.5803, 34.6055, 
    34.63052, 34.65536, 34.68002, 34.70451, 34.72881, 34.75293, 34.77688, 
    34.80064, 34.82423, 34.84763, 34.87085, 34.89389, 34.91674, 34.93942, 
    34.96192, 34.98423, 35.00636, 35.02831, 35.05007, 35.07165, 35.09305, 
    35.11426, 35.13529, 35.15614, 35.1768, 35.19728, 35.21757, 35.23768, 
    35.2576, 35.27734, 35.29689, 35.31625, 35.33543, 35.35443, 35.37324, 
    35.39186, 35.41029, 35.42854, 35.4466, 35.46447, 35.48216, 35.49966, 
    35.51697, 35.53409, 35.55103, 35.56777, 35.58433, 35.6007, 35.61687, 
    35.63287, 35.64867, 35.66428, 35.6797, 35.69493, 35.70997, 35.72483, 
    35.73949, 35.75396, 35.76824, 35.78233, 35.79623, 35.80994, 35.82345, 
    35.83678, 35.84991, 35.86286, 35.87561, 35.88816, 35.90053, 35.91271, 
    35.92469, 35.93648, 35.94808, 35.95948, 35.9707, 35.98171, 35.99254, 
    36.00317, 36.01361, 36.02386, 36.03391, 36.04377, 36.05343, 36.0629, 
    36.07218, 36.08126, 36.09016, 36.09885, 36.10735, 36.11566, 36.12377, 
    36.13168, 36.13941, 36.14693, 36.15427, 36.1614, 36.16835, 36.17509, 
    36.18165, 36.188, 36.19416, 36.20013, 36.2059, 36.21148, 36.21686, 
    36.22204, 36.22703, 36.23182, 36.23642, 36.24082, 36.24502, 36.24903, 
    36.25285, 36.25646, 36.25988, 36.26311, 36.26614, 36.26897, 36.2716, 
    36.27404, 36.27629, 36.27833, 36.28018, 36.28184, 36.28329, 36.28456, 
    36.28562, 36.28649, 36.28716, 36.28764, 36.28792, 36.288, 36.28789, 
    36.28757, 36.28707, 36.28637, 36.28547, 36.28437, 36.28308, 36.28159, 
    36.2799, 36.27802, 36.27594, 36.27367, 36.2712, 36.26853, 36.26567, 
    36.26261, 36.25935, 36.2559, 36.25225, 36.24841, 36.24437, 36.24014, 
    36.2357, 36.23108, 36.22625, 36.22123, 36.21602, 36.21061, 36.205, 
    36.1992, 36.1932, 36.18701, 36.18062, 36.17404, 36.16726, 36.16029, 
    36.15312, 36.14576, 36.1382, 36.13045, 36.1225, 36.11436, 36.10602, 
    36.09749, 36.08876, 36.07984, 36.07073, 36.06142, 36.05192, 36.04222, 
    36.03233, 36.02225, 36.01197, 36.0015, 35.99084, 35.97998, 35.96893, 
    35.95769, 35.94625, 35.93463, 35.92281, 35.91079, 35.89859, 35.88619, 
    35.8736, 35.86082, 35.84785, 35.83468, 35.82133, 35.80778, 35.79404, 
    35.78011, 35.76599, 35.75168, 35.73718, 35.72249, 35.70761, 35.69254, 
    35.67727, 35.66182, 35.64618, 35.63035, 35.61433, 35.59812, 35.58172, 
    35.56513, 35.54836, 35.53139, 35.51424, 35.4969, 35.47937, 35.46166, 
    35.44376, 35.42567, 35.40739, 35.38892, 35.37027, 35.35144, 35.33241, 
    35.31321, 35.29381, 35.27423, 35.25446, 35.23451, 35.21437, 35.19405, 
    35.17354, 35.15285, 35.13198, 35.11092, 35.08968, 35.06825, 35.04664, 
    35.02485, 35.00287, 34.98071, 34.95837, 34.93585, 34.91314, 34.89025, 
    34.86719, 34.84394, 34.82051, 34.79689, 34.7731, 34.74913, 34.72498, 
    34.70065, 34.67613, 34.65144, 34.62657, 34.60152, 34.57629, 34.55088, 
    34.5253, 34.49954, 34.4736, 34.44748, 34.42119, 34.39471, 34.36807, 
    34.34124, 34.31424, 34.28707, 34.25972, 34.23219, 34.20449, 34.17661, 
    34.14856, 34.12033, 34.09193, 34.06336, 34.03461, 34.0057, 33.9766, 
    33.94734, 33.9179, 33.88829, 33.85851, 33.82856, 33.79844, 33.76814, 
    33.73767, 33.70704, 33.67624, 33.64526, 33.61412, 33.5828, 33.55132, 
    33.51967, 33.48785,
  29.94237, 29.98851, 30.03452, 30.08039, 30.12612, 30.17171, 30.21716, 
    30.26247, 30.30764, 30.35267, 30.39756, 30.4423, 30.48691, 30.53137, 
    30.57569, 30.61986, 30.66389, 30.70778, 30.75153, 30.79513, 30.83858, 
    30.88189, 30.92505, 30.96807, 31.01095, 31.05367, 31.09625, 31.13868, 
    31.18097, 31.22311, 31.2651, 31.30694, 31.34863, 31.39017, 31.43157, 
    31.47281, 31.51391, 31.55485, 31.59564, 31.63629, 31.67678, 31.71712, 
    31.75731, 31.79734, 31.83722, 31.87695, 31.91653, 31.95595, 31.99522, 
    32.03434, 32.0733, 32.1121, 32.15075, 32.18924, 32.22758, 32.26577, 
    32.30379, 32.34166, 32.37937, 32.41693, 32.45432, 32.49156, 32.52864, 
    32.56556, 32.60233, 32.63893, 32.67537, 32.71165, 32.74778, 32.78374, 
    32.81954, 32.85518, 32.89066, 32.92598, 32.96113, 32.99612, 33.03095, 
    33.06562, 33.10012, 33.13446, 33.16864, 33.20265, 33.2365, 33.27018, 
    33.30369, 33.33704, 33.37022, 33.40324, 33.4361, 33.46878, 33.5013, 
    33.53365, 33.56583, 33.59785, 33.6297, 33.66137, 33.69288, 33.72422, 
    33.75539, 33.7864, 33.81723, 33.84789, 33.87838, 33.9087, 33.93885, 
    33.96882, 33.99863, 34.02826, 34.05772, 34.08701, 34.11613, 34.14507, 
    34.17384, 34.20243, 34.23085, 34.2591, 34.28717, 34.31507, 34.3428, 
    34.37034, 34.39772, 34.42491, 34.45193, 34.47878, 34.50544, 34.53193, 
    34.55825, 34.58438, 34.61034, 34.63612, 34.66172, 34.68715, 34.71239, 
    34.73746, 34.76234, 34.78705, 34.81158, 34.83593, 34.86009, 34.88408, 
    34.90789, 34.93151, 34.95496, 34.97822, 35.0013, 35.0242, 35.04692, 
    35.06945, 35.0918, 35.11398, 35.13596, 35.15776, 35.17939, 35.20082, 
    35.22207, 35.24314, 35.26403, 35.28473, 35.30524, 35.32557, 35.34571, 
    35.36567, 35.38545, 35.40504, 35.42444, 35.44365, 35.46268, 35.48153, 
    35.50018, 35.51865, 35.53693, 35.55502, 35.57293, 35.59065, 35.60818, 
    35.62552, 35.64267, 35.65964, 35.67641, 35.693, 35.7094, 35.72561, 
    35.74163, 35.75746, 35.7731, 35.78855, 35.80381, 35.81888, 35.83376, 
    35.84845, 35.86295, 35.87726, 35.89137, 35.9053, 35.91903, 35.93258, 
    35.94593, 35.95908, 35.97205, 35.98483, 35.99741, 36.0098, 36.022, 
    36.034, 36.04581, 36.05743, 36.06886, 36.08009, 36.09113, 36.10198, 
    36.11263, 36.12309, 36.13335, 36.14343, 36.15331, 36.16299, 36.17248, 
    36.18177, 36.19087, 36.19978, 36.20849, 36.21701, 36.22533, 36.23346, 
    36.24139, 36.24913, 36.25667, 36.26401, 36.27116, 36.27812, 36.28488, 
    36.29144, 36.29781, 36.30399, 36.30996, 36.31575, 36.32133, 36.32672, 
    36.33192, 36.33691, 36.34171, 36.34632, 36.35073, 36.35494, 36.35896, 
    36.36278, 36.3664, 36.36983, 36.37306, 36.37609, 36.37893, 36.38157, 
    36.38401, 36.38626, 36.38831, 36.39017, 36.39183, 36.39329, 36.39455, 
    36.39562, 36.39649, 36.39716, 36.39764, 36.39791, 36.398, 36.39788, 
    36.39758, 36.39707, 36.39636, 36.39546, 36.39436, 36.39307, 36.39157, 
    36.38989, 36.388, 36.38592, 36.38364, 36.38117, 36.37849, 36.37563, 
    36.37256, 36.3693, 36.36584, 36.36219, 36.35834, 36.35429, 36.35004, 
    36.3456, 36.34097, 36.33614, 36.33111, 36.32588, 36.32046, 36.31485, 
    36.30903, 36.30302, 36.29682, 36.29042, 36.28382, 36.27703, 36.27005, 
    36.26286, 36.25549, 36.24791, 36.24015, 36.23218, 36.22403, 36.21567, 
    36.20713, 36.19838, 36.18945, 36.18032, 36.17099, 36.16147, 36.15176, 
    36.14185, 36.13174, 36.12145, 36.11096, 36.10028, 36.0894, 36.07833, 
    36.06707, 36.05561, 36.04396, 36.03212, 36.02008, 36.00785, 35.99543, 
    35.98282, 35.97001, 35.95702, 35.94383, 35.93045, 35.91687, 35.90311, 
    35.88915, 35.87501, 35.86067, 35.84614, 35.83142, 35.81651, 35.80141, 
    35.78612, 35.77064, 35.75497, 35.73911, 35.72306, 35.70682, 35.69039, 
    35.67377, 35.65697, 35.63997, 35.62279, 35.60542, 35.58786, 35.57011, 
    35.55217, 35.53405, 35.51574, 35.49724, 35.47855, 35.45968, 35.44062, 
    35.42138, 35.40195, 35.38233, 35.36253, 35.34254, 35.32237, 35.30201, 
    35.28146, 35.26073, 35.23982, 35.21872, 35.19744, 35.17598, 35.15433, 
    35.1325, 35.11048, 35.08828, 35.0659, 35.04333, 35.02059, 34.99766, 
    34.97455, 34.95126, 34.92779, 34.90413, 34.8803, 34.85628, 34.83208, 
    34.80771, 34.78315, 34.75842, 34.7335, 34.70841, 34.68314, 34.65768, 
    34.63205, 34.60625, 34.58026, 34.5541, 34.52776, 34.50124, 34.47454, 
    34.44767, 34.42062, 34.3934, 34.366, 34.33842, 34.31067, 34.28275, 
    34.25465, 34.22637, 34.19792, 34.1693, 34.1405, 34.11153, 34.08239, 
    34.05307, 34.02359, 33.99392, 33.96409, 33.93409, 33.90391, 33.87357, 
    33.84305, 33.81236, 33.7815, 33.75047, 33.71928, 33.68791, 33.65637, 
    33.62467, 33.5928,
  30.04147, 30.08769, 30.13376, 30.1797, 30.2255, 30.27116, 30.31668, 
    30.36206, 30.4073, 30.45239, 30.49735, 30.54216, 30.58683, 30.63136, 
    30.67575, 30.71999, 30.76409, 30.80804, 30.85185, 30.89552, 30.93904, 
    30.98242, 31.02565, 31.06874, 31.11167, 31.15447, 31.19711, 31.23961, 
    31.28196, 31.32417, 31.36622, 31.40813, 31.44988, 31.49149, 31.53295, 
    31.57426, 31.61542, 31.65643, 31.69729, 31.738, 31.77855, 31.81895, 
    31.85921, 31.89931, 31.93925, 31.97904, 32.01868, 32.05817, 32.0975, 
    32.13668, 32.1757, 32.21457, 32.25328, 32.29184, 32.33024, 32.36848, 
    32.40657, 32.4445, 32.48228, 32.51989, 32.55735, 32.59465, 32.63179, 
    32.66877, 32.7056, 32.74226, 32.77876, 32.81511, 32.85129, 32.88731, 
    32.92317, 32.95887, 32.99441, 33.02979, 33.065, 33.10005, 33.13493, 
    33.16966, 33.20422, 33.23862, 33.27285, 33.30692, 33.34082, 33.37456, 
    33.40813, 33.44154, 33.47478, 33.50785, 33.54076, 33.5735, 33.60608, 
    33.63848, 33.67072, 33.70279, 33.73469, 33.76642, 33.79799, 33.82938, 
    33.8606, 33.89166, 33.92254, 33.95325, 33.9838, 34.01417, 34.04437, 
    34.0744, 34.10426, 34.13394, 34.16346, 34.19279, 34.22196, 34.25095, 
    34.27977, 34.30842, 34.33689, 34.36518, 34.39331, 34.42126, 34.44903, 
    34.47662, 34.50404, 34.53129, 34.55836, 34.58525, 34.61196, 34.6385, 
    34.66486, 34.69104, 34.71704, 34.74287, 34.76852, 34.79399, 34.81928, 
    34.84439, 34.86932, 34.89407, 34.91864, 34.94304, 34.96724, 34.99128, 
    35.01513, 35.03879, 35.06228, 35.08558, 35.10871, 35.13165, 35.15441, 
    35.17698, 35.19938, 35.22158, 35.24361, 35.26545, 35.28711, 35.30859, 
    35.32988, 35.35099, 35.37191, 35.39265, 35.4132, 35.43357, 35.45375, 
    35.47374, 35.49355, 35.51318, 35.53262, 35.55186, 35.57093, 35.58981, 
    35.60849, 35.627, 35.64531, 35.66344, 35.68138, 35.69913, 35.71669, 
    35.73407, 35.75126, 35.76825, 35.78506, 35.80168, 35.8181, 35.83434, 
    35.8504, 35.86625, 35.88192, 35.8974, 35.91269, 35.92779, 35.9427, 
    35.95741, 35.97194, 35.98627, 36.00042, 36.01437, 36.02813, 36.04169, 
    36.05507, 36.06826, 36.08125, 36.09404, 36.10665, 36.11906, 36.13128, 
    36.14331, 36.15515, 36.16679, 36.17823, 36.18949, 36.20055, 36.21142, 
    36.22209, 36.23257, 36.24286, 36.25294, 36.26284, 36.27254, 36.28205, 
    36.29136, 36.30048, 36.3094, 36.31813, 36.32666, 36.335, 36.34314, 
    36.35109, 36.35884, 36.3664, 36.37376, 36.38092, 36.38789, 36.39466, 
    36.40124, 36.40762, 36.41381, 36.4198, 36.42559, 36.43119, 36.43658, 
    36.44179, 36.4468, 36.45161, 36.45622, 36.46064, 36.46486, 36.46888, 
    36.47271, 36.47634, 36.47977, 36.48301, 36.48605, 36.4889, 36.49154, 
    36.49399, 36.49624, 36.49829, 36.50015, 36.50181, 36.50328, 36.50454, 
    36.50561, 36.50648, 36.50716, 36.50764, 36.50792, 36.508, 36.50788, 
    36.50757, 36.50706, 36.50636, 36.50546, 36.50436, 36.50306, 36.50156, 
    36.49987, 36.49798, 36.4959, 36.49361, 36.49113, 36.48846, 36.48558, 
    36.48251, 36.47924, 36.47578, 36.47212, 36.46826, 36.46421, 36.45995, 
    36.45551, 36.45086, 36.44602, 36.44098, 36.43575, 36.43031, 36.42469, 
    36.41886, 36.41284, 36.40663, 36.40022, 36.3936, 36.3868, 36.3798, 
    36.37261, 36.36522, 36.35763, 36.34985, 36.34187, 36.33369, 36.32533, 
    36.31676, 36.308, 36.29905, 36.2899, 36.28056, 36.27102, 36.26129, 
    36.25136, 36.24124, 36.23092, 36.22041, 36.20971, 36.19881, 36.18772, 
    36.17644, 36.16496, 36.15329, 36.14142, 36.12936, 36.11712, 36.10467, 
    36.09203, 36.0792, 36.06618, 36.05297, 36.03956, 36.02596, 36.01217, 
    35.99819, 35.98402, 35.96965, 35.9551, 35.94035, 35.92542, 35.91029, 
    35.89497, 35.87946, 35.86376, 35.84787, 35.83179, 35.81552, 35.79906, 
    35.78241, 35.76558, 35.74855, 35.73133, 35.71393, 35.69633, 35.67855, 
    35.66058, 35.64243, 35.62408, 35.60555, 35.58683, 35.56792, 35.54883, 
    35.52955, 35.51009, 35.49043, 35.47059, 35.45057, 35.43036, 35.40996, 
    35.38938, 35.36861, 35.34766, 35.32653, 35.30521, 35.2837, 35.26201, 
    35.24014, 35.21809, 35.19585, 35.17342, 35.15082, 35.12803, 35.10506, 
    35.08191, 35.05857, 35.03506, 35.01136, 34.98749, 34.96343, 34.93919, 
    34.91477, 34.89017, 34.86539, 34.84043, 34.81529, 34.78997, 34.76447, 
    34.7388, 34.71294, 34.68691, 34.6607, 34.63431, 34.60775, 34.58101, 
    34.55408, 34.52699, 34.49972, 34.47227, 34.44464, 34.41685, 34.38887, 
    34.36072, 34.3324, 34.3039, 34.27523, 34.24638, 34.21736, 34.18816, 
    34.1588, 34.12926, 34.09954, 34.06966, 34.0396, 34.00938, 33.97898, 
    33.94841, 33.91767, 33.88676, 33.85567, 33.82442, 33.793, 33.76141, 
    33.72965, 33.69773,
  30.14055, 30.18684, 30.23298, 30.27899, 30.32486, 30.37059, 30.41617, 
    30.46162, 30.50693, 30.55209, 30.59711, 30.642, 30.68674, 30.73133, 
    30.77578, 30.82009, 30.86426, 30.90828, 30.95216, 30.9959, 31.03948, 
    31.08293, 31.12622, 31.16938, 31.21238, 31.25524, 31.29795, 31.34052, 
    31.38293, 31.4252, 31.46733, 31.5093, 31.55112, 31.59279, 31.63432, 
    31.67569, 31.71692, 31.75799, 31.79891, 31.83969, 31.8803, 31.92077, 
    31.96109, 32.00125, 32.04126, 32.08112, 32.12082, 32.16037, 32.19976, 
    32.23901, 32.27809, 32.31702, 32.3558, 32.39442, 32.43288, 32.47119, 
    32.50933, 32.54733, 32.58516, 32.62284, 32.66036, 32.69772, 32.73492, 
    32.77197, 32.80885, 32.84557, 32.88214, 32.91854, 32.95478, 32.99086, 
    33.02678, 33.06254, 33.09814, 33.13358, 33.16885, 33.20396, 33.2389, 
    33.27369, 33.3083, 33.34276, 33.37705, 33.41117, 33.44513, 33.47893, 
    33.51256, 33.54602, 33.57932, 33.61245, 33.64541, 33.67821, 33.71083, 
    33.7433, 33.77559, 33.80771, 33.83967, 33.87146, 33.90308, 33.93452, 
    33.9658, 33.99691, 34.02785, 34.05861, 34.08921, 34.11963, 34.14989, 
    34.17997, 34.20988, 34.23961, 34.26918, 34.29857, 34.32779, 34.35683, 
    34.3857, 34.41439, 34.44291, 34.47126, 34.49943, 34.52743, 34.55525, 
    34.58289, 34.61036, 34.63766, 34.66477, 34.69171, 34.71847, 34.74506, 
    34.77146, 34.79769, 34.82374, 34.84961, 34.87531, 34.90082, 34.92616, 
    34.95131, 34.97629, 35.00108, 35.0257, 35.05014, 35.07439, 35.09846, 
    35.12236, 35.14606, 35.16959, 35.19294, 35.21611, 35.23909, 35.26189, 
    35.2845, 35.30694, 35.32919, 35.35126, 35.37314, 35.39484, 35.41635, 
    35.43768, 35.45883, 35.47979, 35.50056, 35.52115, 35.54156, 35.56178, 
    35.58181, 35.60165, 35.62131, 35.64079, 35.66007, 35.67917, 35.69808, 
    35.71681, 35.73534, 35.75369, 35.77185, 35.78983, 35.80761, 35.8252, 
    35.84261, 35.85983, 35.87686, 35.8937, 35.91035, 35.9268, 35.94307, 
    35.95915, 35.97504, 35.99074, 36.00625, 36.02157, 36.03669, 36.05163, 
    36.06637, 36.08092, 36.09529, 36.10946, 36.12344, 36.13722, 36.15081, 
    36.16422, 36.17742, 36.19044, 36.20326, 36.21589, 36.22832, 36.24057, 
    36.25262, 36.26448, 36.27614, 36.28761, 36.29889, 36.30997, 36.32085, 
    36.33155, 36.34204, 36.35235, 36.36246, 36.37238, 36.3821, 36.39162, 
    36.40095, 36.41008, 36.41903, 36.42777, 36.43632, 36.44467, 36.45283, 
    36.46079, 36.46856, 36.47613, 36.4835, 36.49068, 36.49766, 36.50445, 
    36.51104, 36.51743, 36.52363, 36.52963, 36.53543, 36.54104, 36.54645, 
    36.55166, 36.55668, 36.5615, 36.56612, 36.57055, 36.57478, 36.57881, 
    36.58265, 36.58628, 36.58972, 36.59296, 36.59601, 36.59886, 36.60151, 
    36.60396, 36.60622, 36.60828, 36.61014, 36.6118, 36.61327, 36.61454, 
    36.61561, 36.61648, 36.61716, 36.61763, 36.61792, 36.618, 36.61789, 
    36.61757, 36.61706, 36.61636, 36.61545, 36.61435, 36.61305, 36.61155, 
    36.60986, 36.60796, 36.60587, 36.60359, 36.6011, 36.59842, 36.59554, 
    36.59246, 36.58919, 36.58572, 36.58205, 36.57819, 36.57412, 36.56986, 
    36.5654, 36.56075, 36.5559, 36.55085, 36.54561, 36.54016, 36.53453, 
    36.52869, 36.52266, 36.51643, 36.51001, 36.50339, 36.49657, 36.48956, 
    36.48235, 36.47494, 36.46734, 36.45955, 36.45155, 36.44336, 36.43498, 
    36.4264, 36.41762, 36.40865, 36.39949, 36.39013, 36.38057, 36.37082, 
    36.36087, 36.35073, 36.3404, 36.32987, 36.31915, 36.30823, 36.29712, 
    36.28581, 36.27431, 36.26262, 36.25073, 36.23865, 36.22637, 36.21391, 
    36.20124, 36.18839, 36.17535, 36.16211, 36.14867, 36.13505, 36.12123, 
    36.10723, 36.09303, 36.07864, 36.06405, 36.04928, 36.03431, 36.01916, 
    36.00381, 35.98827, 35.97254, 35.95662, 35.94051, 35.92421, 35.90772, 
    35.89104, 35.87418, 35.85712, 35.83987, 35.82243, 35.80481, 35.78699, 
    35.76899, 35.7508, 35.73243, 35.71386, 35.6951, 35.67616, 35.65703, 
    35.63772, 35.61821, 35.59853, 35.57865, 35.55859, 35.53834, 35.51791, 
    35.49729, 35.47648, 35.45549, 35.43432, 35.41296, 35.39142, 35.36969, 
    35.34778, 35.32568, 35.3034, 35.28094, 35.25829, 35.23547, 35.21246, 
    35.18926, 35.16589, 35.14233, 35.11859, 35.09467, 35.07056, 35.04628, 
    35.02182, 34.99717, 34.97235, 34.94735, 34.92216, 34.8968, 34.87125, 
    34.84554, 34.81963, 34.79356, 34.7673, 34.74086, 34.71425, 34.68746, 
    34.66049, 34.63335, 34.60603, 34.57853, 34.55086, 34.52301, 34.49499, 
    34.46679, 34.43842, 34.40987, 34.38114, 34.35225, 34.32317, 34.29393, 
    34.26451, 34.23492, 34.20516, 34.17522, 34.14511, 34.11483, 34.08438, 
    34.05376, 34.02296, 33.992, 33.96087, 33.92956, 33.89809, 33.86644, 
    33.83463, 33.80264,
  30.23961, 30.28597, 30.33218, 30.37826, 30.42419, 30.46999, 30.51565, 
    30.56116, 30.60653, 30.65177, 30.69686, 30.74181, 30.78662, 30.83128, 
    30.8758, 30.92018, 30.96441, 31.0085, 31.05245, 31.09625, 31.1399, 
    31.18341, 31.22678, 31.27, 31.31307, 31.356, 31.39877, 31.4414, 31.48389, 
    31.52622, 31.56841, 31.61045, 31.65234, 31.69407, 31.73566, 31.7771, 
    31.81839, 31.85953, 31.90052, 31.94135, 31.98204, 32.02257, 32.06295, 
    32.10318, 32.14325, 32.18317, 32.22294, 32.26255, 32.30201, 32.34132, 
    32.38047, 32.41946, 32.45829, 32.49698, 32.5355, 32.57387, 32.61208, 
    32.65014, 32.68803, 32.72577, 32.76336, 32.80078, 32.83804, 32.87514, 
    32.91209, 32.94887, 32.9855, 33.02196, 33.05826, 33.0944, 33.13038, 
    33.1662, 33.20185, 33.23735, 33.27268, 33.30785, 33.34285, 33.37769, 
    33.41237, 33.44688, 33.48123, 33.51541, 33.54943, 33.58328, 33.61697, 
    33.65049, 33.68384, 33.71703, 33.75005, 33.7829, 33.81559, 33.8481, 
    33.88045, 33.91263, 33.94464, 33.97648, 34.00815, 34.03965, 34.07099, 
    34.10215, 34.13314, 34.16396, 34.19461, 34.22509, 34.25539, 34.28552, 
    34.31548, 34.34527, 34.37489, 34.40433, 34.4336, 34.46269, 34.49161, 
    34.52036, 34.54893, 34.57733, 34.60555, 34.63359, 34.66146, 34.68916, 
    34.71667, 34.74401, 34.77118, 34.79816, 34.82497, 34.8516, 34.87806, 
    34.90434, 34.93043, 34.95635, 34.98209, 35.00765, 35.03303, 35.05823, 
    35.08325, 35.10809, 35.13275, 35.15723, 35.18153, 35.20564, 35.22958, 
    35.25333, 35.2769, 35.30029, 35.3235, 35.34652, 35.36936, 35.39202, 
    35.4145, 35.43679, 35.45889, 35.48082, 35.50256, 35.52411, 35.54548, 
    35.56666, 35.58766, 35.60847, 35.6291, 35.64954, 35.6698, 35.68987, 
    35.70975, 35.72944, 35.74895, 35.76828, 35.78741, 35.80635, 35.82512, 
    35.84369, 35.86207, 35.88026, 35.89827, 35.91608, 35.93371, 35.95115, 
    35.9684, 35.98546, 36.00233, 36.01901, 36.0355, 36.0518, 36.06791, 
    36.08383, 36.09956, 36.11509, 36.13044, 36.1456, 36.16056, 36.17533, 
    36.18991, 36.2043, 36.21849, 36.2325, 36.24631, 36.25993, 36.27335, 
    36.28659, 36.29963, 36.31247, 36.32513, 36.33759, 36.34985, 36.36193, 
    36.37381, 36.38549, 36.39698, 36.40828, 36.41938, 36.43029, 36.441, 
    36.45152, 36.46185, 36.47197, 36.48191, 36.49165, 36.50119, 36.51054, 
    36.51969, 36.52864, 36.53741, 36.54597, 36.55434, 36.56252, 36.57049, 
    36.57827, 36.58586, 36.59325, 36.60044, 36.60743, 36.61423, 36.62083, 
    36.62724, 36.63345, 36.63946, 36.64528, 36.65089, 36.65631, 36.66154, 
    36.66656, 36.67139, 36.67602, 36.68046, 36.6847, 36.68874, 36.69258, 
    36.69622, 36.69967, 36.70292, 36.70597, 36.70882, 36.71148, 36.71394, 
    36.71619, 36.71826, 36.72012, 36.72179, 36.72326, 36.72453, 36.72561, 
    36.72648, 36.72715, 36.72763, 36.72792, 36.728, 36.72789, 36.72757, 
    36.72706, 36.72635, 36.72544, 36.72434, 36.72304, 36.72154, 36.71984, 
    36.71795, 36.71585, 36.71356, 36.71107, 36.70838, 36.7055, 36.70242, 
    36.69913, 36.69566, 36.69198, 36.68811, 36.68404, 36.67977, 36.6753, 
    36.67064, 36.66578, 36.66072, 36.65547, 36.65002, 36.64437, 36.63852, 
    36.63248, 36.62624, 36.6198, 36.61317, 36.60634, 36.59931, 36.59209, 
    36.58467, 36.57705, 36.56924, 36.56123, 36.55303, 36.54463, 36.53603, 
    36.52724, 36.51825, 36.50907, 36.49969, 36.49012, 36.48035, 36.47038, 
    36.46022, 36.44987, 36.43932, 36.42858, 36.41764, 36.40651, 36.39518, 
    36.38366, 36.37194, 36.36003, 36.34793, 36.33563, 36.32314, 36.31046, 
    36.29758, 36.28451, 36.27124, 36.25779, 36.24414, 36.2303, 36.21626, 
    36.20203, 36.18762, 36.17301, 36.1582, 36.14321, 36.12803, 36.11265, 
    36.09708, 36.08133, 36.06538, 36.04924, 36.03291, 36.01638, 35.99968, 
    35.98277, 35.96568, 35.94841, 35.93093, 35.91328, 35.89543, 35.8774, 
    35.85917, 35.84076, 35.82216, 35.80337, 35.78439, 35.76523, 35.74588, 
    35.72634, 35.70662, 35.6867, 35.66661, 35.64632, 35.62585, 35.60519, 
    35.58435, 35.56332, 35.54211, 35.52071, 35.49913, 35.47736, 35.45541, 
    35.43327, 35.41095, 35.38845, 35.36576, 35.34289, 35.31984, 35.2966, 
    35.27319, 35.24959, 35.2258, 35.20184, 35.1777, 35.15337, 35.12886, 
    35.10417, 35.0793, 35.05425, 35.02903, 35.00362, 34.97803, 34.95226, 
    34.92632, 34.90019, 34.87389, 34.8474, 34.82074, 34.79391, 34.76689, 
    34.7397, 34.71233, 34.68479, 34.65707, 34.62917, 34.60109, 34.57285, 
    34.54442, 34.51582, 34.48705, 34.4581, 34.42898, 34.39968, 34.37022, 
    34.34057, 34.31076, 34.28077, 34.25061, 34.22028, 34.18977, 34.1591, 
    34.12825, 34.09723, 34.06604, 34.03468, 34.00315, 33.97145, 33.93959, 
    33.90755,
  30.33865, 30.38507, 30.43136, 30.4775, 30.52351, 30.56937, 30.6151, 
    30.66068, 30.70612, 30.75142, 30.79658, 30.8416, 30.88647, 30.93121, 
    30.97579, 31.02024, 31.06454, 31.1087, 31.15271, 31.19658, 31.2403, 
    31.28388, 31.32731, 31.3706, 31.41373, 31.45673, 31.49957, 31.54227, 
    31.58482, 31.62722, 31.66947, 31.71158, 31.75353, 31.79534, 31.83699, 
    31.8785, 31.91985, 31.96105, 32.00211, 32.04301, 32.08376, 32.12435, 
    32.16479, 32.20509, 32.24523, 32.28521, 32.32504, 32.36472, 32.40424, 
    32.44361, 32.48282, 32.52187, 32.56078, 32.59952, 32.63811, 32.67654, 
    32.71481, 32.75293, 32.79089, 32.82869, 32.86633, 32.90381, 32.94114, 
    32.9783, 33.01531, 33.05215, 33.08884, 33.12536, 33.16172, 33.19793, 
    33.23396, 33.26984, 33.30556, 33.34111, 33.3765, 33.41173, 33.44679, 
    33.48169, 33.51642, 33.55099, 33.5854, 33.61964, 33.65371, 33.68762, 
    33.72137, 33.75494, 33.78835, 33.82159, 33.85467, 33.88758, 33.92032, 
    33.95289, 33.98529, 34.01753, 34.04959, 34.08149, 34.11322, 34.14478, 
    34.17616, 34.20737, 34.23842, 34.26929, 34.3, 34.33052, 34.36088, 
    34.39107, 34.42108, 34.45092, 34.48059, 34.51008, 34.5394, 34.56855, 
    34.59752, 34.62631, 34.65493, 34.68338, 34.71165, 34.73975, 34.76767, 
    34.79541, 34.82297, 34.85036, 34.87757, 34.90461, 34.93147, 34.95815, 
    34.98465, 35.01097, 35.03711, 35.06307, 35.08886, 35.11446, 35.13989, 
    35.16513, 35.1902, 35.21509, 35.23979, 35.26431, 35.28865, 35.31282, 
    35.33679, 35.36059, 35.3842, 35.40763, 35.43089, 35.45395, 35.47683, 
    35.49953, 35.52205, 35.54438, 35.56652, 35.58849, 35.61026, 35.63186, 
    35.65327, 35.67449, 35.69553, 35.71638, 35.73704, 35.75752, 35.77781, 
    35.79792, 35.81784, 35.83757, 35.85711, 35.87647, 35.89564, 35.91462, 
    35.93341, 35.95202, 35.97044, 35.98867, 36.00671, 36.02456, 36.04222, 
    36.05968, 36.07697, 36.09406, 36.11096, 36.12767, 36.14419, 36.16052, 
    36.17666, 36.19261, 36.20837, 36.22393, 36.23931, 36.25449, 36.26949, 
    36.28428, 36.29889, 36.3133, 36.32753, 36.34156, 36.3554, 36.36904, 
    36.38249, 36.39575, 36.40881, 36.42168, 36.43436, 36.44685, 36.45913, 
    36.47123, 36.48313, 36.49484, 36.50635, 36.51767, 36.52879, 36.53972, 
    36.55046, 36.56099, 36.57134, 36.58149, 36.59144, 36.6012, 36.61076, 
    36.62012, 36.62929, 36.63826, 36.64704, 36.65562, 36.66401, 36.6722, 
    36.68019, 36.68798, 36.69559, 36.70299, 36.71019, 36.7172, 36.72401, 
    36.73063, 36.73705, 36.74327, 36.74929, 36.75512, 36.76075, 36.76617, 
    36.77141, 36.77644, 36.78128, 36.78592, 36.79037, 36.79461, 36.79866, 
    36.80251, 36.80616, 36.80961, 36.81287, 36.81593, 36.81879, 36.82145, 
    36.82391, 36.82617, 36.82824, 36.83011, 36.83178, 36.83325, 36.83452, 
    36.8356, 36.83648, 36.83715, 36.83764, 36.83792, 36.838, 36.83788, 
    36.83757, 36.83706, 36.83635, 36.83544, 36.83434, 36.83303, 36.83153, 
    36.82983, 36.82793, 36.82583, 36.82353, 36.82104, 36.81834, 36.81546, 
    36.81237, 36.80908, 36.8056, 36.80191, 36.79803, 36.79395, 36.78968, 
    36.7852, 36.78053, 36.77566, 36.7706, 36.76533, 36.75987, 36.75421, 
    36.74835, 36.7423, 36.73605, 36.7296, 36.72295, 36.71611, 36.70907, 
    36.70183, 36.6944, 36.68677, 36.67894, 36.67092, 36.6627, 36.65428, 
    36.64567, 36.63686, 36.62785, 36.61865, 36.60926, 36.59966, 36.58988, 
    36.57989, 36.56971, 36.55934, 36.54877, 36.53801, 36.52705, 36.51589, 
    36.50454, 36.493, 36.48126, 36.46933, 36.4572, 36.44489, 36.43237, 
    36.41966, 36.40676, 36.39367, 36.38037, 36.36689, 36.35322, 36.33935, 
    36.32529, 36.31104, 36.29659, 36.28196, 36.26712, 36.25211, 36.23689, 
    36.22149, 36.20589, 36.1901, 36.17412, 36.15795, 36.14159, 36.12504, 
    36.1083, 36.09137, 36.07425, 36.05693, 36.03944, 36.02174, 36.00386, 
    35.98579, 35.96754, 35.94909, 35.93045, 35.91163, 35.89262, 35.87342, 
    35.85403, 35.83446, 35.8147, 35.79475, 35.77462, 35.7543, 35.73378, 
    35.71309, 35.69221, 35.67114, 35.64989, 35.62846, 35.60683, 35.58503, 
    35.56303, 35.54086, 35.5185, 35.49595, 35.47322, 35.45031, 35.42722, 
    35.40394, 35.38048, 35.35684, 35.33301, 35.30901, 35.28482, 35.26044, 
    35.23589, 35.21116, 35.18625, 35.16116, 35.13588, 35.11043, 35.08479, 
    35.05898, 35.03299, 35.00681, 34.98046, 34.95393, 34.92723, 34.90034, 
    34.87328, 34.84604, 34.81862, 34.79103, 34.76326, 34.73531, 34.70719, 
    34.67889, 34.65042, 34.62177, 34.59295, 34.56395, 34.53477, 34.50543, 
    34.47591, 34.44621, 34.41634, 34.38631, 34.35609, 34.32571, 34.29515, 
    34.26442, 34.23352, 34.20245, 34.17121, 34.13979, 34.10821, 34.07646, 
    34.04453, 34.01244,
  30.43766, 30.48415, 30.53051, 30.57672, 30.6228, 30.66873, 30.71452, 
    30.76017, 30.80569, 30.85105, 30.89628, 30.94137, 30.98631, 31.03111, 
    31.07577, 31.12028, 31.16465, 31.20887, 31.25295, 31.29689, 31.34068, 
    31.38432, 31.42782, 31.47117, 31.51438, 31.55744, 31.60035, 31.64311, 
    31.68573, 31.7282, 31.77052, 31.81269, 31.85471, 31.89658, 31.9383, 
    31.97987, 32.02129, 32.06256, 32.10367, 32.14464, 32.18545, 32.22611, 
    32.26662, 32.30698, 32.34718, 32.38723, 32.42712, 32.46687, 32.50645, 
    32.54588, 32.58516, 32.62428, 32.66324, 32.70205, 32.7407, 32.77919, 
    32.81752, 32.85571, 32.89373, 32.93159, 32.96929, 33.00684, 33.04422, 
    33.08145, 33.11851, 33.15542, 33.19216, 33.22875, 33.26517, 33.30143, 
    33.33753, 33.37347, 33.40924, 33.44485, 33.4803, 33.51559, 33.55071, 
    33.58567, 33.62046, 33.65509, 33.68955, 33.72385, 33.75798, 33.79195, 
    33.82575, 33.85938, 33.89285, 33.92615, 33.95928, 33.99224, 34.02504, 
    34.05767, 34.09013, 34.12242, 34.15454, 34.18649, 34.21827, 34.24988, 
    34.28132, 34.31259, 34.34369, 34.37461, 34.40537, 34.43595, 34.46636, 
    34.4966, 34.52667, 34.55656, 34.58628, 34.61582, 34.64519, 34.67439, 
    34.70341, 34.73226, 34.76093, 34.78942, 34.81775, 34.84589, 34.87386, 
    34.90165, 34.92926, 34.9567, 34.98396, 35.01104, 35.03795, 35.06467, 
    35.09122, 35.11759, 35.14378, 35.16979, 35.19562, 35.22127, 35.24675, 
    35.27203, 35.29715, 35.32207, 35.34682, 35.37139, 35.39577, 35.41998, 
    35.444, 35.46784, 35.4915, 35.51497, 35.53826, 35.56137, 35.58429, 
    35.60703, 35.62959, 35.65196, 35.67415, 35.69615, 35.71797, 35.7396, 
    35.76105, 35.78231, 35.80339, 35.82428, 35.84498, 35.86549, 35.88582, 
    35.90597, 35.92592, 35.94569, 35.96527, 35.98466, 36.00387, 36.02288, 
    36.04171, 36.06035, 36.0788, 36.09706, 36.11514, 36.13302, 36.15071, 
    36.16822, 36.18553, 36.20266, 36.21959, 36.23633, 36.25288, 36.26924, 
    36.28541, 36.30139, 36.31718, 36.33277, 36.34818, 36.36339, 36.37841, 
    36.39323, 36.40787, 36.42231, 36.43656, 36.45061, 36.46448, 36.47815, 
    36.49163, 36.50491, 36.518, 36.53089, 36.54359, 36.5561, 36.56841, 
    36.58053, 36.59246, 36.60419, 36.61572, 36.62706, 36.6382, 36.64915, 
    36.65991, 36.67047, 36.68083, 36.69099, 36.70097, 36.71074, 36.72032, 
    36.72971, 36.73889, 36.74788, 36.75668, 36.76527, 36.77368, 36.78188, 
    36.78989, 36.7977, 36.80531, 36.81273, 36.81995, 36.82697, 36.8338, 
    36.84042, 36.84686, 36.85308, 36.85912, 36.86496, 36.8706, 36.87604, 
    36.88128, 36.88633, 36.89117, 36.89582, 36.90028, 36.90453, 36.90858, 
    36.91244, 36.9161, 36.91956, 36.92282, 36.92588, 36.92875, 36.93142, 
    36.93388, 36.93615, 36.93822, 36.94009, 36.94176, 36.94324, 36.94452, 
    36.94559, 36.94647, 36.94715, 36.94763, 36.94791, 36.948, 36.94788, 
    36.94757, 36.94706, 36.94635, 36.94544, 36.94433, 36.94302, 36.94151, 
    36.93981, 36.93791, 36.93581, 36.93351, 36.93101, 36.92831, 36.92541, 
    36.92232, 36.91903, 36.91553, 36.91184, 36.90796, 36.90387, 36.89959, 
    36.8951, 36.89042, 36.88554, 36.88047, 36.87519, 36.86972, 36.86405, 
    36.85818, 36.85211, 36.84585, 36.83939, 36.83273, 36.82587, 36.81882, 
    36.81157, 36.80412, 36.79648, 36.78864, 36.7806, 36.77236, 36.76393, 
    36.7553, 36.74648, 36.73745, 36.72823, 36.71882, 36.70921, 36.6994, 
    36.6894, 36.6792, 36.66881, 36.65822, 36.64743, 36.63646, 36.62528, 
    36.61391, 36.60234, 36.59058, 36.57863, 36.56648, 36.55413, 36.5416, 
    36.52887, 36.51594, 36.50282, 36.48951, 36.476, 36.4623, 36.44841, 
    36.43432, 36.42004, 36.40557, 36.3909, 36.37605, 36.361, 36.34575, 
    36.33032, 36.31469, 36.29888, 36.28287, 36.26667, 36.25028, 36.2337, 
    36.21692, 36.19996, 36.1828, 36.16546, 36.14793, 36.1302, 36.11229, 
    36.09419, 36.0759, 36.05742, 36.03875, 36.01989, 36.00084, 35.98161, 
    35.96218, 35.94258, 35.92278, 35.90279, 35.88262, 35.86226, 35.84172, 
    35.82098, 35.80006, 35.77896, 35.75767, 35.73619, 35.71453, 35.69268, 
    35.67065, 35.64843, 35.62603, 35.60345, 35.58068, 35.55773, 35.53459, 
    35.51127, 35.48777, 35.46408, 35.44021, 35.41616, 35.39193, 35.36752, 
    35.34292, 35.31815, 35.29319, 35.26805, 35.24273, 35.21723, 35.19155, 
    35.16569, 35.13965, 35.11343, 35.08703, 35.06046, 35.0337, 35.00677, 
    34.97966, 34.95237, 34.92491, 34.89726, 34.86945, 34.84145, 34.81328, 
    34.78493, 34.7564, 34.72771, 34.69883, 34.66978, 34.64056, 34.61116, 
    34.58159, 34.55184, 34.52192, 34.49183, 34.46156, 34.43113, 34.40052, 
    34.36974, 34.33878, 34.30766, 34.27636, 34.24489, 34.21325, 34.18145, 
    34.14947, 34.11732,
  30.53665, 30.58321, 30.62963, 30.67592, 30.72206, 30.76806, 30.81392, 
    30.85965, 30.90522, 30.95066, 30.99596, 31.04111, 31.08612, 31.13099, 
    31.17572, 31.2203, 31.26473, 31.30903, 31.35317, 31.39718, 31.44103, 
    31.48475, 31.52831, 31.57173, 31.615, 31.65813, 31.70111, 31.74394, 
    31.78662, 31.82915, 31.87154, 31.91377, 31.95586, 31.9978, 32.03959, 
    32.08122, 32.1227, 32.16404, 32.20522, 32.24625, 32.28713, 32.32786, 
    32.36843, 32.40885, 32.44912, 32.48923, 32.52919, 32.56899, 32.60864, 
    32.64814, 32.68747, 32.72665, 32.76568, 32.80455, 32.84327, 32.88182, 
    32.92022, 32.95846, 32.99654, 33.03447, 33.07224, 33.10984, 33.14729, 
    33.18457, 33.2217, 33.25867, 33.29547, 33.33212, 33.3686, 33.40492, 
    33.44108, 33.47708, 33.51291, 33.54858, 33.58409, 33.61944, 33.65462, 
    33.68963, 33.72448, 33.75917, 33.79369, 33.82805, 33.86224, 33.89626, 
    33.93012, 33.96381, 33.99733, 34.03069, 34.06388, 34.0969, 34.12975, 
    34.16243, 34.19495, 34.22729, 34.25947, 34.29147, 34.32331, 34.35498, 
    34.38647, 34.41779, 34.44894, 34.47993, 34.51073, 34.54137, 34.57183, 
    34.60212, 34.63224, 34.66219, 34.69196, 34.72155, 34.75097, 34.78022, 
    34.80929, 34.83819, 34.86691, 34.89546, 34.92383, 34.95202, 34.98004, 
    35.00788, 35.03555, 35.06303, 35.09034, 35.11747, 35.14442, 35.1712, 
    35.19779, 35.22421, 35.25044, 35.2765, 35.30238, 35.32807, 35.35359, 
    35.37893, 35.40408, 35.42906, 35.45385, 35.47846, 35.50289, 35.52714, 
    35.5512, 35.57508, 35.59879, 35.6223, 35.64563, 35.66878, 35.69175, 
    35.71453, 35.73713, 35.75954, 35.78176, 35.80381, 35.82567, 35.84734, 
    35.86882, 35.89013, 35.91124, 35.93217, 35.95291, 35.97346, 35.99383, 
    36.01401, 36.034, 36.05381, 36.07342, 36.09285, 36.11209, 36.13115, 
    36.15001, 36.16868, 36.18716, 36.20546, 36.22357, 36.24148, 36.25921, 
    36.27674, 36.29409, 36.31124, 36.32821, 36.34499, 36.36157, 36.37796, 
    36.39416, 36.41017, 36.42598, 36.44161, 36.45704, 36.47228, 36.48733, 
    36.50218, 36.51685, 36.53131, 36.54559, 36.55967, 36.57356, 36.58726, 
    36.60076, 36.61407, 36.62718, 36.6401, 36.65282, 36.66536, 36.67769, 
    36.68983, 36.70178, 36.71353, 36.72509, 36.73645, 36.74761, 36.75858, 
    36.76936, 36.77994, 36.79032, 36.80051, 36.8105, 36.82029, 36.82989, 
    36.83929, 36.84849, 36.8575, 36.86631, 36.87493, 36.88334, 36.89156, 
    36.89959, 36.90741, 36.91504, 36.92247, 36.9297, 36.93674, 36.94358, 
    36.95022, 36.95666, 36.96291, 36.96895, 36.9748, 36.98045, 36.9859, 
    36.99115, 36.99621, 37.00106, 37.00573, 37.01019, 37.01445, 37.01851, 
    37.02237, 37.02604, 37.0295, 37.03277, 37.03584, 37.03871, 37.04138, 
    37.04385, 37.04613, 37.0482, 37.05008, 37.05175, 37.05323, 37.05451, 
    37.05559, 37.05647, 37.05715, 37.05763, 37.05791, 37.058, 37.05788, 
    37.05757, 37.05706, 37.05634, 37.05543, 37.05432, 37.05301, 37.0515, 
    37.04979, 37.04789, 37.04578, 37.04348, 37.04097, 37.03827, 37.03537, 
    37.03227, 37.02897, 37.02547, 37.02177, 37.01788, 37.01379, 37.00949, 
    37.005, 37.00031, 36.99542, 36.99034, 36.98505, 36.97957, 36.97389, 
    36.96801, 36.96193, 36.95565, 36.94918, 36.94251, 36.93564, 36.92857, 
    36.92131, 36.91385, 36.90619, 36.89833, 36.89028, 36.88203, 36.87358, 
    36.86493, 36.85609, 36.84705, 36.83781, 36.82838, 36.81875, 36.80893, 
    36.79891, 36.78869, 36.77827, 36.76767, 36.75686, 36.74586, 36.73466, 
    36.72327, 36.71169, 36.6999, 36.68793, 36.67575, 36.66339, 36.65083, 
    36.63807, 36.62512, 36.61197, 36.59864, 36.5851, 36.57138, 36.55746, 
    36.54334, 36.52904, 36.51454, 36.49984, 36.48496, 36.46988, 36.45461, 
    36.43915, 36.42349, 36.40765, 36.39161, 36.37538, 36.35896, 36.34234, 
    36.32554, 36.30854, 36.29136, 36.27398, 36.25642, 36.23866, 36.22071, 
    36.20258, 36.18425, 36.16574, 36.14703, 36.12814, 36.10906, 36.08979, 
    36.07033, 36.05069, 36.03085, 36.01083, 35.99062, 35.97022, 35.94964, 
    35.92887, 35.90791, 35.88677, 35.86544, 35.84392, 35.82222, 35.80033, 
    35.77826, 35.756, 35.73357, 35.71094, 35.68813, 35.66513, 35.64196, 
    35.61859, 35.59505, 35.57132, 35.54741, 35.52332, 35.49904, 35.47458, 
    35.44994, 35.42512, 35.40012, 35.37493, 35.34957, 35.32402, 35.29829, 
    35.27239, 35.2463, 35.22004, 35.1936, 35.16697, 35.14017, 35.11319, 
    35.08603, 35.05869, 35.03118, 35.00349, 34.97562, 34.94757, 34.91935, 
    34.89095, 34.86238, 34.83363, 34.80471, 34.7756, 34.74633, 34.71688, 
    34.68726, 34.65746, 34.62749, 34.59734, 34.56702, 34.53653, 34.50587, 
    34.47504, 34.44403, 34.41285, 34.3815, 34.34998, 34.31829, 34.28642, 
    34.25439, 34.22219,
  30.63562, 30.68225, 30.72874, 30.77509, 30.8213, 30.86737, 30.9133, 
    30.95909, 31.00474, 31.05025, 31.09561, 31.14083, 31.18591, 31.23085, 
    31.27564, 31.32029, 31.3648, 31.40916, 31.45337, 31.49744, 31.54137, 
    31.58515, 31.62878, 31.67227, 31.71561, 31.7588, 31.80184, 31.84474, 
    31.88749, 31.93009, 31.97254, 32.01484, 32.057, 32.099, 32.14085, 
    32.18255, 32.2241, 32.2655, 32.30675, 32.34785, 32.38879, 32.42958, 
    32.47022, 32.5107, 32.55103, 32.59121, 32.63123, 32.6711, 32.71081, 
    32.75037, 32.78977, 32.82902, 32.86811, 32.90704, 32.94582, 32.98444, 
    33.0229, 33.0612, 33.09935, 33.13733, 33.17516, 33.21283, 33.25034, 
    33.28769, 33.32487, 33.3619, 33.39877, 33.43547, 33.47202, 33.5084, 
    33.54462, 33.58067, 33.61657, 33.6523, 33.68787, 33.72327, 33.75851, 
    33.79358, 33.8285, 33.86324, 33.89782, 33.93223, 33.96648, 34.00056, 
    34.03448, 34.06823, 34.1018, 34.13522, 34.16846, 34.20154, 34.23445, 
    34.26719, 34.29976, 34.33216, 34.36439, 34.39645, 34.42834, 34.46006, 
    34.49161, 34.52298, 34.55419, 34.58522, 34.61609, 34.64677, 34.67729, 
    34.70763, 34.7378, 34.7678, 34.79762, 34.82727, 34.85674, 34.88604, 
    34.91516, 34.94411, 34.97289, 35.00148, 35.0299, 35.05814, 35.08621, 
    35.1141, 35.14182, 35.16935, 35.1967, 35.22388, 35.25089, 35.27771, 
    35.30435, 35.33081, 35.35709, 35.3832, 35.40912, 35.43486, 35.46043, 
    35.48581, 35.51101, 35.53603, 35.56087, 35.58552, 35.61, 35.63428, 
    35.65839, 35.68232, 35.70606, 35.72962, 35.753, 35.77619, 35.79919, 
    35.82202, 35.84466, 35.86711, 35.88938, 35.91146, 35.93336, 35.95507, 
    35.9766, 35.99794, 36.01909, 36.04005, 36.06083, 36.08142, 36.10183, 
    36.12205, 36.14207, 36.16192, 36.18157, 36.20103, 36.22031, 36.2394, 
    36.25829, 36.277, 36.29552, 36.31385, 36.33199, 36.34994, 36.3677, 
    36.38527, 36.40265, 36.41983, 36.43683, 36.45364, 36.47025, 36.48667, 
    36.5029, 36.51894, 36.53479, 36.55044, 36.5659, 36.58117, 36.59624, 
    36.61113, 36.62582, 36.64031, 36.65461, 36.66872, 36.68264, 36.69636, 
    36.70989, 36.72322, 36.73636, 36.74931, 36.76205, 36.77461, 36.78697, 
    36.79913, 36.8111, 36.82288, 36.83445, 36.84584, 36.85702, 36.86801, 
    36.87881, 36.8894, 36.89981, 36.91002, 36.92002, 36.92984, 36.93945, 
    36.94887, 36.95809, 36.96712, 36.97594, 36.98458, 36.99301, 37.00124, 
    37.00928, 37.01712, 37.02477, 37.03221, 37.03946, 37.04651, 37.05336, 
    37.06001, 37.06647, 37.07272, 37.07878, 37.08464, 37.0903, 37.09576, 
    37.10102, 37.10609, 37.11096, 37.11562, 37.12009, 37.12436, 37.12843, 
    37.13231, 37.13597, 37.13945, 37.14272, 37.1458, 37.14867, 37.15135, 
    37.15383, 37.15611, 37.15818, 37.16006, 37.16174, 37.16322, 37.16451, 
    37.16558, 37.16647, 37.16715, 37.16763, 37.16792, 37.168, 37.16788, 
    37.16757, 37.16705, 37.16634, 37.16543, 37.16431, 37.163, 37.16149, 
    37.15978, 37.15787, 37.15576, 37.15345, 37.15094, 37.14823, 37.14532, 
    37.14222, 37.13891, 37.13541, 37.13171, 37.1278, 37.1237, 37.1194, 
    37.1149, 37.1102, 37.1053, 37.1002, 37.09491, 37.08942, 37.08372, 
    37.07784, 37.07175, 37.06546, 37.05897, 37.05229, 37.04541, 37.03833, 
    37.03105, 37.02357, 37.0159, 37.00803, 36.99995, 36.99169, 36.98322, 
    36.97456, 36.9657, 36.95665, 36.9474, 36.93794, 36.9283, 36.91845, 
    36.90841, 36.89817, 36.88774, 36.87711, 36.86629, 36.85527, 36.84405, 
    36.83263, 36.82103, 36.80922, 36.79722, 36.78503, 36.77264, 36.76005, 
    36.74727, 36.73429, 36.72113, 36.70776, 36.6942, 36.68045, 36.6665, 
    36.65237, 36.63803, 36.6235, 36.60878, 36.59387, 36.57877, 36.56347, 
    36.54797, 36.53229, 36.51641, 36.50035, 36.48409, 36.46763, 36.45099, 
    36.43415, 36.41713, 36.39991, 36.3825, 36.3649, 36.34711, 36.32914, 
    36.31097, 36.29261, 36.27406, 36.25532, 36.23639, 36.21727, 36.19797, 
    36.17847, 36.15879, 36.13892, 36.11886, 36.09861, 36.07818, 36.05756, 
    36.03675, 36.01575, 35.99457, 35.9732, 35.95165, 35.92991, 35.90798, 
    35.88587, 35.86357, 35.84109, 35.81842, 35.79557, 35.77253, 35.74931, 
    35.72591, 35.70232, 35.67855, 35.65459, 35.63046, 35.60614, 35.58163, 
    35.55695, 35.53209, 35.50703, 35.48181, 35.45639, 35.43081, 35.40503, 
    35.37908, 35.35295, 35.32664, 35.30014, 35.27348, 35.24662, 35.2196, 
    35.19239, 35.165, 35.13744, 35.1097, 35.08178, 35.05369, 35.02542, 
    34.99697, 34.96835, 34.93954, 34.91057, 34.88142, 34.85209, 34.82259, 
    34.79292, 34.76307, 34.73304, 34.70285, 34.67247, 34.64193, 34.61121, 
    34.58033, 34.54926, 34.51803, 34.48663, 34.45505, 34.42331, 34.39139, 
    34.3593, 34.32704,
  30.73456, 30.78126, 30.82782, 30.87424, 30.92052, 30.96666, 31.01266, 
    31.05852, 31.10424, 31.14981, 31.19525, 31.24054, 31.28568, 31.33069, 
    31.37555, 31.42027, 31.46484, 31.50927, 31.55355, 31.59769, 31.64168, 
    31.68553, 31.72923, 31.77278, 31.81619, 31.85945, 31.90256, 31.94552, 
    31.98834, 32.03101, 32.07352, 32.11589, 32.15811, 32.20018, 32.2421, 
    32.28386, 32.32548, 32.36694, 32.40826, 32.44942, 32.49043, 32.53128, 
    32.57199, 32.61253, 32.65293, 32.69317, 32.73326, 32.77319, 32.81297, 
    32.85259, 32.89206, 32.93136, 32.97052, 33.00951, 33.04835, 33.08703, 
    33.12556, 33.16392, 33.20213, 33.24018, 33.27807, 33.3158, 33.35337, 
    33.39078, 33.42803, 33.46511, 33.50204, 33.53881, 33.57541, 33.61185, 
    33.64814, 33.68425, 33.72021, 33.756, 33.79162, 33.82709, 33.86238, 
    33.89752, 33.93249, 33.96729, 34.00193, 34.0364, 34.07071, 34.10485, 
    34.13882, 34.17262, 34.20626, 34.23973, 34.27303, 34.30616, 34.33913, 
    34.37193, 34.40455, 34.437, 34.46929, 34.50141, 34.53335, 34.56513, 
    34.59673, 34.62816, 34.65942, 34.69051, 34.72142, 34.75217, 34.78273, 
    34.81313, 34.84335, 34.8734, 34.90328, 34.93298, 34.9625, 34.99185, 
    35.02103, 35.05003, 35.07885, 35.10749, 35.13596, 35.16426, 35.19238, 
    35.22031, 35.24807, 35.27566, 35.30306, 35.33029, 35.35734, 35.38421, 
    35.4109, 35.43741, 35.46374, 35.48989, 35.51586, 35.54165, 35.56726, 
    35.59268, 35.61793, 35.64299, 35.66788, 35.69258, 35.71709, 35.74143, 
    35.76558, 35.78955, 35.81334, 35.83694, 35.86036, 35.88359, 35.90664, 
    35.9295, 35.95218, 35.97467, 35.99698, 36.01911, 36.04104, 36.06279, 
    36.08436, 36.10574, 36.12693, 36.14793, 36.16875, 36.18938, 36.20982, 
    36.23008, 36.25014, 36.27002, 36.28971, 36.30921, 36.32852, 36.34764, 
    36.36658, 36.38532, 36.40387, 36.42224, 36.44041, 36.45839, 36.47618, 
    36.49379, 36.5112, 36.52842, 36.54544, 36.56228, 36.57893, 36.59538, 
    36.61164, 36.62771, 36.64358, 36.65927, 36.67476, 36.69005, 36.70516, 
    36.72007, 36.73479, 36.74931, 36.76364, 36.77777, 36.79172, 36.80546, 
    36.81902, 36.83237, 36.84554, 36.85851, 36.87128, 36.88386, 36.89624, 
    36.90843, 36.92042, 36.93222, 36.94382, 36.95522, 36.96643, 36.97744, 
    36.98825, 36.99887, 37.0093, 37.01952, 37.02955, 37.03938, 37.04902, 
    37.05845, 37.06769, 37.07673, 37.08558, 37.09423, 37.10267, 37.11093, 
    37.11898, 37.12683, 37.13449, 37.14195, 37.14921, 37.15627, 37.16314, 
    37.1698, 37.17627, 37.18254, 37.18861, 37.19448, 37.20015, 37.20562, 
    37.2109, 37.21597, 37.22085, 37.22552, 37.23, 37.23428, 37.23836, 
    37.24223, 37.24591, 37.24939, 37.25267, 37.25576, 37.25864, 37.26132, 
    37.2638, 37.26608, 37.26817, 37.27005, 37.27173, 37.27321, 37.2745, 
    37.27558, 37.27646, 37.27715, 37.27763, 37.27792, 37.278, 37.27789, 
    37.27757, 37.27705, 37.27634, 37.27542, 37.27431, 37.27299, 37.27148, 
    37.26976, 37.26785, 37.26574, 37.26342, 37.26091, 37.25819, 37.25528, 
    37.25217, 37.24886, 37.24535, 37.24163, 37.23772, 37.23362, 37.22931, 
    37.2248, 37.22009, 37.21518, 37.21008, 37.20477, 37.19927, 37.19357, 
    37.18766, 37.18156, 37.17526, 37.16876, 37.16207, 37.15517, 37.14808, 
    37.14079, 37.13329, 37.12561, 37.11772, 37.10963, 37.10135, 37.09287, 
    37.08419, 37.07532, 37.06624, 37.05697, 37.0475, 37.03784, 37.02798, 
    37.01792, 37.00766, 36.99721, 36.98656, 36.97571, 36.96467, 36.95343, 
    36.94199, 36.93036, 36.91854, 36.90651, 36.89429, 36.88188, 36.86927, 
    36.85647, 36.84347, 36.83027, 36.81689, 36.8033, 36.78952, 36.77555, 
    36.76138, 36.74702, 36.73247, 36.71772, 36.70278, 36.68764, 36.67232, 
    36.6568, 36.64108, 36.62518, 36.60908, 36.59279, 36.57631, 36.55963, 
    36.54277, 36.52571, 36.50846, 36.49102, 36.47338, 36.45556, 36.43755, 
    36.41935, 36.40095, 36.38237, 36.3636, 36.34464, 36.32548, 36.30614, 
    36.28661, 36.26689, 36.24698, 36.22689, 36.2066, 36.18613, 36.16547, 
    36.14462, 36.12359, 36.10237, 36.08096, 36.05937, 36.03759, 36.01562, 
    35.99347, 35.97113, 35.9486, 35.9259, 35.903, 35.87992, 35.85666, 
    35.83321, 35.80959, 35.78577, 35.76177, 35.73759, 35.71323, 35.68868, 
    35.66395, 35.63904, 35.61395, 35.58867, 35.56322, 35.53758, 35.51176, 
    35.48576, 35.45959, 35.43323, 35.40669, 35.37997, 35.35307, 35.326, 
    35.29874, 35.27131, 35.24369, 35.2159, 35.18794, 35.15979, 35.13147, 
    35.10297, 35.0743, 35.04545, 35.01642, 34.98722, 34.95784, 34.92829, 
    34.89856, 34.86866, 34.83858, 34.80833, 34.77791, 34.74731, 34.71655, 
    34.6856, 34.65449, 34.6232, 34.59174, 34.56011, 34.52831, 34.49634, 
    34.4642, 34.43188,
  30.83348, 30.88024, 30.92687, 30.97337, 31.01972, 31.06593, 31.11199, 
    31.15792, 31.20371, 31.24935, 31.29485, 31.34021, 31.38543, 31.4305, 
    31.47543, 31.52022, 31.56486, 31.60935, 31.65371, 31.69791, 31.74197, 
    31.78589, 31.82965, 31.87328, 31.91675, 31.96008, 32.00325, 32.04628, 
    32.08916, 32.1319, 32.17448, 32.21692, 32.2592, 32.30134, 32.34332, 
    32.38515, 32.42684, 32.46837, 32.50975, 32.55097, 32.59204, 32.63297, 
    32.67373, 32.71435, 32.75481, 32.79511, 32.83527, 32.87526, 32.9151, 
    32.95479, 32.99432, 33.03369, 33.07291, 33.11197, 33.15087, 33.18961, 
    33.2282, 33.26663, 33.3049, 33.34301, 33.38096, 33.41875, 33.45638, 
    33.49385, 33.53117, 33.56831, 33.6053, 33.64213, 33.67879, 33.7153, 
    33.75164, 33.78782, 33.82383, 33.85968, 33.89537, 33.93089, 33.96624, 
    34.00144, 34.03646, 34.07133, 34.10603, 34.14056, 34.17492, 34.20911, 
    34.24314, 34.27701, 34.3107, 34.34423, 34.37759, 34.41078, 34.4438, 
    34.47665, 34.50933, 34.54184, 34.57418, 34.60635, 34.63836, 34.67019, 
    34.70184, 34.73333, 34.76464, 34.79578, 34.82675, 34.85755, 34.88817, 
    34.91862, 34.94889, 34.97899, 35.00892, 35.03867, 35.06825, 35.09765, 
    35.12688, 35.15593, 35.1848, 35.2135, 35.24202, 35.27036, 35.29853, 
    35.32652, 35.35432, 35.38196, 35.40941, 35.43669, 35.46378, 35.4907, 
    35.51744, 35.54399, 35.57037, 35.59657, 35.62259, 35.64842, 35.67408, 
    35.69955, 35.72484, 35.74995, 35.77488, 35.79962, 35.82418, 35.84856, 
    35.87276, 35.89677, 35.9206, 35.94424, 35.9677, 35.99098, 36.01407, 
    36.03698, 36.0597, 36.08223, 36.10458, 36.12675, 36.14872, 36.17051, 
    36.19212, 36.21354, 36.23477, 36.25581, 36.27666, 36.29733, 36.31781, 
    36.3381, 36.35821, 36.37812, 36.39785, 36.41739, 36.43673, 36.45589, 
    36.47486, 36.49363, 36.51222, 36.53062, 36.54883, 36.56684, 36.58467, 
    36.6023, 36.61975, 36.637, 36.65406, 36.67093, 36.6876, 36.70408, 
    36.72038, 36.73647, 36.75238, 36.76809, 36.78361, 36.79893, 36.81407, 
    36.82901, 36.84375, 36.8583, 36.87266, 36.88682, 36.90079, 36.91456, 
    36.92814, 36.94152, 36.95471, 36.9677, 36.9805, 36.99311, 37.00551, 
    37.01772, 37.02974, 37.04155, 37.05318, 37.0646, 37.07583, 37.08686, 
    37.0977, 37.10834, 37.11878, 37.12902, 37.13907, 37.14892, 37.15858, 
    37.16803, 37.17729, 37.18635, 37.19521, 37.20387, 37.21234, 37.2206, 
    37.22868, 37.23655, 37.24422, 37.25169, 37.25896, 37.26604, 37.27292, 
    37.2796, 37.28608, 37.29235, 37.29844, 37.30432, 37.31, 37.31548, 
    37.32077, 37.32585, 37.33074, 37.33542, 37.33991, 37.34419, 37.34828, 
    37.35217, 37.35585, 37.35934, 37.36263, 37.36571, 37.3686, 37.37128, 
    37.37377, 37.37606, 37.37815, 37.38003, 37.38172, 37.38321, 37.38449, 
    37.38557, 37.38646, 37.38715, 37.38763, 37.38792, 37.388, 37.38788, 
    37.38757, 37.38705, 37.38633, 37.38542, 37.3843, 37.38298, 37.38147, 
    37.37975, 37.37783, 37.37571, 37.37339, 37.37088, 37.36816, 37.36524, 
    37.36212, 37.3588, 37.35528, 37.35157, 37.34765, 37.34353, 37.33921, 
    37.33469, 37.32998, 37.32506, 37.31995, 37.31463, 37.30912, 37.3034, 
    37.29749, 37.29137, 37.28506, 37.27855, 37.27184, 37.26493, 37.25783, 
    37.25052, 37.24302, 37.23531, 37.22741, 37.21931, 37.21101, 37.20251, 
    37.19382, 37.18493, 37.17584, 37.16655, 37.15706, 37.14738, 37.1375, 
    37.12742, 37.11714, 37.10667, 37.096, 37.08513, 37.07407, 37.06281, 
    37.05135, 37.0397, 37.02785, 37.0158, 37.00356, 36.99112, 36.97849, 
    36.96566, 36.95264, 36.93942, 36.92601, 36.9124, 36.89859, 36.88459, 
    36.8704, 36.85601, 36.84143, 36.82666, 36.81169, 36.79652, 36.78117, 
    36.76562, 36.74987, 36.73394, 36.71781, 36.70149, 36.68497, 36.66827, 
    36.65137, 36.63428, 36.617, 36.59953, 36.58186, 36.56401, 36.54596, 
    36.52772, 36.5093, 36.49068, 36.47187, 36.45287, 36.43368, 36.41431, 
    36.39474, 36.37498, 36.35504, 36.33491, 36.31459, 36.29408, 36.27338, 
    36.25249, 36.23142, 36.21016, 36.18871, 36.16708, 36.14526, 36.12325, 
    36.10106, 36.07868, 36.05611, 36.03336, 36.01043, 35.98731, 35.964, 
    35.94051, 35.91684, 35.89298, 35.86894, 35.84472, 35.82031, 35.79572, 
    35.77095, 35.74599, 35.72085, 35.69553, 35.67003, 35.64435, 35.61848, 
    35.59244, 35.56621, 35.53981, 35.51322, 35.48645, 35.45951, 35.43238, 
    35.40508, 35.3776, 35.34994, 35.3221, 35.29408, 35.26589, 35.23752, 
    35.20897, 35.18024, 35.15134, 35.12226, 35.09301, 35.06358, 35.03398, 
    35.0042, 34.97424, 34.94411, 34.91381, 34.88334, 34.85269, 34.82187, 
    34.79087, 34.7597, 34.72836, 34.69685, 34.66516, 34.6333, 34.60128, 
    34.56908, 34.53671,
  30.93237, 30.97921, 31.02591, 31.07247, 31.11889, 31.16516, 31.2113, 
    31.2573, 31.30316, 31.34887, 31.39444, 31.43987, 31.48515, 31.53029, 
    31.57529, 31.62015, 31.66485, 31.70942, 31.75384, 31.79811, 31.84224, 
    31.88622, 31.93006, 31.97375, 32.01729, 32.06068, 32.10393, 32.14703, 
    32.18997, 32.23277, 32.27542, 32.31792, 32.36028, 32.40248, 32.44453, 
    32.48643, 32.52818, 32.56977, 32.61121, 32.65251, 32.69365, 32.73463, 
    32.77546, 32.81614, 32.85667, 32.89704, 32.93725, 32.97731, 33.01722, 
    33.05697, 33.09656, 33.136, 33.17528, 33.2144, 33.25336, 33.29218, 
    33.33082, 33.36931, 33.40765, 33.44582, 33.48383, 33.52169, 33.55938, 
    33.59691, 33.63428, 33.6715, 33.70855, 33.74543, 33.78216, 33.81872, 
    33.85513, 33.89136, 33.92744, 33.96334, 33.99909, 34.03467, 34.07009, 
    34.10534, 34.14043, 34.17535, 34.21011, 34.24469, 34.27911, 34.31337, 
    34.34746, 34.38138, 34.41513, 34.44871, 34.48213, 34.51537, 34.54845, 
    34.58136, 34.6141, 34.64666, 34.67906, 34.71129, 34.74334, 34.77523, 
    34.80694, 34.83848, 34.86985, 34.90104, 34.93206, 34.96291, 34.99359, 
    35.02409, 35.05442, 35.08457, 35.11455, 35.14436, 35.17398, 35.20344, 
    35.23272, 35.26182, 35.29074, 35.31949, 35.34806, 35.37645, 35.40467, 
    35.4327, 35.46057, 35.48825, 35.51575, 35.54308, 35.57022, 35.59718, 
    35.62397, 35.65057, 35.677, 35.70324, 35.72931, 35.75519, 35.78089, 
    35.80641, 35.83175, 35.8569, 35.88187, 35.90666, 35.93127, 35.95569, 
    35.97993, 36.00398, 36.02785, 36.05154, 36.07505, 36.09836, 36.1215, 
    36.14444, 36.16721, 36.18978, 36.21217, 36.23438, 36.2564, 36.27822, 
    36.29987, 36.32133, 36.3426, 36.36368, 36.38457, 36.40528, 36.4258, 
    36.44613, 36.46627, 36.48622, 36.50598, 36.52555, 36.54493, 36.56413, 
    36.58313, 36.60194, 36.62057, 36.639, 36.65724, 36.67529, 36.69315, 
    36.71082, 36.72829, 36.74557, 36.76266, 36.77956, 36.79627, 36.81279, 
    36.82911, 36.84523, 36.86117, 36.87691, 36.89246, 36.90781, 36.92298, 
    36.93794, 36.95272, 36.96729, 36.98168, 36.99586, 37.00986, 37.02366, 
    37.03726, 37.05067, 37.06388, 37.0769, 37.08973, 37.10235, 37.11478, 
    37.12701, 37.13905, 37.15089, 37.16254, 37.17398, 37.18523, 37.19629, 
    37.20715, 37.2178, 37.22826, 37.23853, 37.2486, 37.25846, 37.26814, 
    37.27761, 37.28688, 37.29596, 37.30484, 37.31352, 37.322, 37.33028, 
    37.33837, 37.34625, 37.35394, 37.36143, 37.36872, 37.3758, 37.3827, 
    37.38939, 37.39588, 37.40217, 37.40826, 37.41416, 37.41985, 37.42535, 
    37.43064, 37.43573, 37.44063, 37.44532, 37.44981, 37.45411, 37.4582, 
    37.4621, 37.46579, 37.46928, 37.47258, 37.47567, 37.47856, 37.48125, 
    37.48375, 37.48604, 37.48813, 37.49002, 37.49171, 37.49319, 37.49448, 
    37.49557, 37.49646, 37.49714, 37.49763, 37.49791, 37.498, 37.49788, 
    37.49757, 37.49705, 37.49633, 37.49541, 37.49429, 37.49297, 37.49145, 
    37.48973, 37.48781, 37.48569, 37.48336, 37.48084, 37.47812, 37.47519, 
    37.47207, 37.46875, 37.46522, 37.46149, 37.45757, 37.45345, 37.44912, 
    37.44459, 37.43987, 37.43494, 37.42981, 37.42449, 37.41896, 37.41324, 
    37.40731, 37.40119, 37.39487, 37.38834, 37.38162, 37.3747, 37.36758, 
    37.36026, 37.35274, 37.34502, 37.3371, 37.32899, 37.32067, 37.31216, 
    37.30345, 37.29454, 37.28543, 37.27612, 37.26662, 37.25692, 37.24702, 
    37.23692, 37.22662, 37.21613, 37.20544, 37.19455, 37.18347, 37.17219, 
    37.16071, 37.14903, 37.13716, 37.12509, 37.11283, 37.10036, 37.08771, 
    37.07486, 37.06181, 37.04856, 37.03513, 37.02149, 37.00766, 36.99363, 
    36.97942, 36.965, 36.95039, 36.93559, 36.92059, 36.9054, 36.89001, 
    36.87444, 36.85866, 36.8427, 36.82654, 36.81018, 36.79364, 36.7769, 
    36.75997, 36.74285, 36.72554, 36.70803, 36.69033, 36.67245, 36.65437, 
    36.63609, 36.61763, 36.59898, 36.58014, 36.5611, 36.54188, 36.52247, 
    36.50286, 36.48307, 36.46309, 36.44292, 36.42256, 36.40202, 36.38128, 
    36.36036, 36.33924, 36.31795, 36.29646, 36.27478, 36.25293, 36.23088, 
    36.20864, 36.18623, 36.16362, 36.14083, 36.11785, 36.09469, 36.07134, 
    36.04781, 36.02409, 36.00019, 35.9761, 35.95184, 35.92739, 35.90275, 
    35.87793, 35.85293, 35.82775, 35.80238, 35.77684, 35.75111, 35.7252, 
    35.6991, 35.67283, 35.64638, 35.61974, 35.59293, 35.56594, 35.53876, 
    35.51141, 35.48388, 35.45617, 35.42828, 35.40022, 35.37197, 35.34355, 
    35.31495, 35.28618, 35.25723, 35.2281, 35.19879, 35.16931, 35.13965, 
    35.10982, 35.07981, 35.04963, 35.01928, 34.98875, 34.95805, 34.92717, 
    34.89612, 34.8649, 34.8335, 34.80193, 34.7702, 34.73829, 34.7062, 
    34.67395, 34.64153,
  31.03124, 31.07815, 31.12492, 31.17155, 31.21803, 31.26438, 31.31059, 
    31.35666, 31.40258, 31.44836, 31.494, 31.5395, 31.58485, 31.63006, 
    31.67513, 31.72005, 31.76483, 31.80946, 31.85395, 31.89829, 31.94249, 
    31.98654, 32.03044, 32.0742, 32.11781, 32.16127, 32.20458, 32.24774, 
    32.29076, 32.33363, 32.37634, 32.41891, 32.46133, 32.50359, 32.54571, 
    32.58768, 32.62949, 32.67115, 32.71266, 32.75402, 32.79522, 32.83628, 
    32.87717, 32.91792, 32.95851, 32.99894, 33.03922, 33.07935, 33.11932, 
    33.15913, 33.19879, 33.23829, 33.27763, 33.31682, 33.35585, 33.39472, 
    33.43343, 33.47198, 33.51038, 33.54861, 33.58669, 33.6246, 33.66236, 
    33.69995, 33.73739, 33.77466, 33.81177, 33.84872, 33.88551, 33.92213, 
    33.9586, 33.99489, 34.03102, 34.067, 34.1028, 34.13844, 34.17392, 
    34.20923, 34.24438, 34.27936, 34.31417, 34.34882, 34.3833, 34.41761, 
    34.45176, 34.48573, 34.51954, 34.55318, 34.58665, 34.61996, 34.65309, 
    34.68605, 34.71885, 34.75147, 34.78393, 34.81621, 34.84832, 34.88026, 
    34.91203, 34.94362, 34.97504, 35.00629, 35.03737, 35.06827, 35.099, 
    35.12955, 35.15993, 35.19014, 35.22017, 35.25003, 35.27971, 35.30922, 
    35.33854, 35.36769, 35.39667, 35.42547, 35.45409, 35.48253, 35.5108, 
    35.53889, 35.5668, 35.59453, 35.62208, 35.64945, 35.67664, 35.70366, 
    35.73049, 35.75714, 35.78362, 35.80991, 35.83602, 35.86194, 35.88769, 
    35.91325, 35.93864, 35.96384, 35.98885, 36.01369, 36.03834, 36.06281, 
    36.08709, 36.11119, 36.13511, 36.15884, 36.18238, 36.20574, 36.22892, 
    36.25191, 36.27471, 36.29733, 36.31976, 36.342, 36.36406, 36.38593, 
    36.40762, 36.42911, 36.45042, 36.47154, 36.49247, 36.51322, 36.53377, 
    36.55414, 36.57432, 36.59431, 36.61411, 36.63371, 36.65313, 36.67236, 
    36.6914, 36.71025, 36.7289, 36.74737, 36.76564, 36.78373, 36.80162, 
    36.81932, 36.83683, 36.85415, 36.87127, 36.8882, 36.90494, 36.92148, 
    36.93783, 36.95399, 36.96996, 36.98573, 37.00131, 37.01669, 37.03188, 
    37.04688, 37.06168, 37.07628, 37.09069, 37.10491, 37.11893, 37.13276, 
    37.14639, 37.15982, 37.17306, 37.1861, 37.19894, 37.21159, 37.22405, 
    37.23631, 37.24836, 37.26023, 37.27189, 37.28336, 37.29464, 37.30571, 
    37.31659, 37.32727, 37.33775, 37.34803, 37.35812, 37.368, 37.37769, 
    37.38718, 37.39648, 37.40557, 37.41447, 37.42316, 37.43166, 37.43996, 
    37.44806, 37.45596, 37.46367, 37.47116, 37.47847, 37.48557, 37.49247, 
    37.49918, 37.50568, 37.51199, 37.51809, 37.524, 37.5297, 37.53521, 
    37.54051, 37.54561, 37.55052, 37.55522, 37.55972, 37.56403, 37.56813, 
    37.57203, 37.57573, 37.57923, 37.58253, 37.58563, 37.58852, 37.59122, 
    37.59372, 37.59601, 37.59811, 37.6, 37.60169, 37.60319, 37.60448, 
    37.60557, 37.60645, 37.60714, 37.60763, 37.60791, 37.608, 37.60788, 
    37.60757, 37.60705, 37.60633, 37.60541, 37.60429, 37.60296, 37.60144, 
    37.59972, 37.59779, 37.59566, 37.59334, 37.59081, 37.58808, 37.58515, 
    37.58202, 37.57869, 37.57516, 37.57143, 37.56749, 37.56336, 37.55902, 
    37.55449, 37.54976, 37.54482, 37.53968, 37.53435, 37.52881, 37.52308, 
    37.51714, 37.51101, 37.50467, 37.49813, 37.4914, 37.48446, 37.47733, 
    37.46999, 37.46246, 37.45473, 37.44679, 37.43866, 37.43033, 37.4218, 
    37.41307, 37.40415, 37.39502, 37.3857, 37.37617, 37.36646, 37.35654, 
    37.34642, 37.3361, 37.32559, 37.31488, 37.30397, 37.29287, 37.28156, 
    37.27006, 37.25837, 37.24647, 37.23438, 37.22209, 37.20961, 37.19693, 
    37.18405, 37.17097, 37.15771, 37.14424, 37.13058, 37.11672, 37.10267, 
    37.08842, 37.07398, 37.05935, 37.04452, 37.02949, 37.01427, 36.99886, 
    36.98325, 36.96745, 36.95145, 36.93526, 36.91888, 36.9023, 36.88553, 
    36.86857, 36.85142, 36.83407, 36.81653, 36.7988, 36.78088, 36.76277, 
    36.74446, 36.72597, 36.70728, 36.6884, 36.66933, 36.65007, 36.63062, 
    36.61098, 36.59116, 36.57114, 36.55093, 36.53053, 36.50995, 36.48917, 
    36.46821, 36.44706, 36.42572, 36.4042, 36.38248, 36.36058, 36.3385, 
    36.31622, 36.29376, 36.27111, 36.24828, 36.22526, 36.20206, 36.17867, 
    36.15509, 36.13133, 36.10739, 36.08326, 36.05895, 36.03445, 36.00977, 
    35.98491, 35.95987, 35.93464, 35.90923, 35.88363, 35.85786, 35.8319, 
    35.80576, 35.77944, 35.75294, 35.72626, 35.6994, 35.67236, 35.64513, 
    35.61773, 35.59015, 35.56239, 35.53446, 35.50634, 35.47805, 35.44957, 
    35.42093, 35.3921, 35.36309, 35.33392, 35.30456, 35.27503, 35.24532, 
    35.21544, 35.18538, 35.15514, 35.12473, 35.09415, 35.06339, 35.03246, 
    35.00136, 34.97008, 34.93863, 34.90701, 34.87522, 34.84325, 34.81111, 
    34.7788, 34.74632,
  31.13008, 31.17706, 31.2239, 31.2706, 31.31716, 31.36357, 31.40985, 
    31.45599, 31.50198, 31.54783, 31.59354, 31.63911, 31.68453, 31.72981, 
    31.77494, 31.81993, 31.86478, 31.90948, 31.95404, 31.99845, 32.04271, 
    32.08683, 32.1308, 32.17462, 32.2183, 32.26183, 32.30521, 32.34844, 
    32.39152, 32.43446, 32.47724, 32.51987, 32.56236, 32.60469, 32.64688, 
    32.68891, 32.73079, 32.77251, 32.81409, 32.85551, 32.89678, 32.9379, 
    32.97886, 33.01967, 33.06033, 33.10083, 33.14117, 33.18136, 33.22139, 
    33.26127, 33.30099, 33.34056, 33.37997, 33.41922, 33.45831, 33.49724, 
    33.53602, 33.57463, 33.61309, 33.65139, 33.68953, 33.7275, 33.76532, 
    33.80298, 33.84048, 33.87781, 33.91498, 33.95199, 33.98884, 34.02553, 
    34.06205, 34.09841, 34.1346, 34.17063, 34.2065, 34.2422, 34.27773, 
    34.31311, 34.34831, 34.38335, 34.41822, 34.45293, 34.48746, 34.52184, 
    34.55604, 34.59007, 34.62394, 34.65764, 34.69117, 34.72453, 34.75772, 
    34.79074, 34.82359, 34.85627, 34.88878, 34.92112, 34.95328, 34.98528, 
    35.0171, 35.04875, 35.08022, 35.11153, 35.14266, 35.17361, 35.2044, 
    35.235, 35.26544, 35.2957, 35.32578, 35.35569, 35.38542, 35.41498, 
    35.44436, 35.47356, 35.50259, 35.53144, 35.56011, 35.5886, 35.61692, 
    35.64506, 35.67302, 35.7008, 35.7284, 35.75582, 35.78306, 35.81012, 
    35.837, 35.8637, 35.89022, 35.91656, 35.94272, 35.96869, 35.99448, 
    36.0201, 36.04552, 36.07077, 36.09583, 36.12071, 36.1454, 36.16992, 
    36.19424, 36.21839, 36.24235, 36.26612, 36.28971, 36.31311, 36.33633, 
    36.35936, 36.38221, 36.40487, 36.42734, 36.44962, 36.47172, 36.49363, 
    36.51535, 36.53689, 36.55824, 36.5794, 36.60037, 36.62115, 36.64175, 
    36.66215, 36.68237, 36.70239, 36.72223, 36.74187, 36.76133, 36.78059, 
    36.79966, 36.81855, 36.83724, 36.85574, 36.87405, 36.89216, 36.91009, 
    36.92782, 36.94536, 36.96271, 36.97987, 36.99683, 37.0136, 37.03017, 
    37.04656, 37.06275, 37.07874, 37.09454, 37.11015, 37.12556, 37.14078, 
    37.1558, 37.17063, 37.18526, 37.1997, 37.21395, 37.22799, 37.24184, 
    37.2555, 37.26896, 37.28222, 37.29529, 37.30816, 37.32084, 37.33331, 
    37.34559, 37.35767, 37.36956, 37.38125, 37.39274, 37.40403, 37.41513, 
    37.42603, 37.43673, 37.44723, 37.45753, 37.46764, 37.47754, 37.48725, 
    37.49676, 37.50607, 37.51518, 37.5241, 37.53281, 37.54132, 37.54964, 
    37.55775, 37.56567, 37.57339, 37.5809, 37.58822, 37.59534, 37.60225, 
    37.60897, 37.61549, 37.6218, 37.62792, 37.63383, 37.63955, 37.64507, 
    37.65038, 37.65549, 37.6604, 37.66512, 37.66963, 37.67394, 37.67805, 
    37.68196, 37.68567, 37.68917, 37.69248, 37.69558, 37.69849, 37.70119, 
    37.70369, 37.70599, 37.70809, 37.70999, 37.71168, 37.71318, 37.71447, 
    37.71556, 37.71645, 37.71714, 37.71763, 37.71791, 37.718, 37.71788, 
    37.71756, 37.71704, 37.71632, 37.7154, 37.71428, 37.71295, 37.71143, 
    37.7097, 37.70777, 37.70564, 37.70331, 37.70078, 37.69804, 37.69511, 
    37.69197, 37.68863, 37.68509, 37.68135, 37.67741, 37.67327, 37.66893, 
    37.66439, 37.65964, 37.6547, 37.64955, 37.64421, 37.63866, 37.63291, 
    37.62696, 37.62082, 37.61447, 37.60792, 37.60117, 37.59422, 37.58707, 
    37.57973, 37.57218, 37.56443, 37.55648, 37.54834, 37.53999, 37.53144, 
    37.5227, 37.51376, 37.50461, 37.49527, 37.48573, 37.47599, 37.46605, 
    37.45592, 37.44558, 37.43505, 37.42432, 37.41339, 37.40226, 37.39094, 
    37.37941, 37.36769, 37.35578, 37.34366, 37.33135, 37.31884, 37.30614, 
    37.29324, 37.28014, 37.26685, 37.25335, 37.23967, 37.22578, 37.21171, 
    37.19743, 37.18296, 37.1683, 37.15344, 37.13839, 37.12314, 37.10769, 
    37.09206, 37.07623, 37.0602, 37.04398, 37.02757, 37.01096, 36.99416, 
    36.97717, 36.95998, 36.9426, 36.92503, 36.90727, 36.88931, 36.87116, 
    36.85283, 36.83429, 36.81557, 36.79666, 36.77755, 36.75826, 36.73877, 
    36.7191, 36.69923, 36.67918, 36.65894, 36.6385, 36.61788, 36.59706, 
    36.57607, 36.55487, 36.5335, 36.51193, 36.49018, 36.46824, 36.44611, 
    36.42379, 36.40129, 36.3786, 36.35573, 36.33267, 36.30942, 36.28599, 
    36.26237, 36.23857, 36.21458, 36.19041, 36.16605, 36.14151, 36.11679, 
    36.09188, 36.06679, 36.04152, 36.01606, 35.99042, 35.9646, 35.93859, 
    35.91241, 35.88604, 35.85949, 35.83276, 35.80585, 35.77876, 35.7515, 
    35.72404, 35.69641, 35.66861, 35.64062, 35.61245, 35.58411, 35.55559, 
    35.52689, 35.49801, 35.46896, 35.43972, 35.41032, 35.38073, 35.35097, 
    35.32103, 35.29092, 35.26064, 35.23018, 35.19954, 35.16873, 35.13774, 
    35.10659, 35.07526, 35.04375, 35.01207, 34.98022, 34.9482, 34.91601, 
    34.88365, 34.85111,
  31.2289, 31.27595, 31.32286, 31.36963, 31.41626, 31.46274, 31.50909, 
    31.5553, 31.60136, 31.64728, 31.69306, 31.73869, 31.78418, 31.82953, 
    31.87473, 31.91979, 31.96471, 32.00948, 32.0541, 32.09858, 32.14291, 
    32.1871, 32.23114, 32.27503, 32.31877, 32.36237, 32.40582, 32.44912, 
    32.49226, 32.53527, 32.57812, 32.62082, 32.66337, 32.70577, 32.74802, 
    32.79012, 32.83206, 32.87386, 32.9155, 32.95699, 32.99832, 33.03951, 
    33.08053, 33.12141, 33.16213, 33.20269, 33.2431, 33.28336, 33.32345, 
    33.3634, 33.40318, 33.44281, 33.48228, 33.5216, 33.56075, 33.59975, 
    33.63859, 33.67727, 33.71579, 33.75415, 33.79235, 33.83039, 33.86827, 
    33.90599, 33.94355, 33.98094, 34.01818, 34.05525, 34.09216, 34.1289, 
    34.16549, 34.2019, 34.23816, 34.27425, 34.31018, 34.34594, 34.38153, 
    34.41696, 34.45223, 34.48732, 34.52225, 34.55702, 34.59162, 34.62605, 
    34.66031, 34.6944, 34.72832, 34.76208, 34.79567, 34.82909, 34.86233, 
    34.89541, 34.92831, 34.96105, 34.99361, 35.02601, 35.05823, 35.09028, 
    35.12216, 35.15386, 35.18539, 35.21675, 35.24794, 35.27895, 35.30978, 
    35.34044, 35.37093, 35.40124, 35.43138, 35.46134, 35.49112, 35.52073, 
    35.55017, 35.57942, 35.6085, 35.6374, 35.66612, 35.69466, 35.72303, 
    35.75122, 35.77923, 35.80706, 35.83471, 35.86217, 35.88947, 35.91658, 
    35.9435, 35.97025, 35.99682, 36.0232, 36.04941, 36.07543, 36.10127, 
    36.12693, 36.1524, 36.17769, 36.2028, 36.22772, 36.25246, 36.27702, 
    36.30139, 36.32558, 36.34958, 36.3734, 36.39703, 36.42048, 36.44373, 
    36.46681, 36.48969, 36.51239, 36.53491, 36.55724, 36.57937, 36.60133, 
    36.62309, 36.64466, 36.66605, 36.68725, 36.70826, 36.72908, 36.74971, 
    36.77015, 36.79041, 36.81047, 36.83034, 36.85002, 36.86951, 36.88881, 
    36.90792, 36.92684, 36.94557, 36.9641, 36.98244, 37.0006, 37.01855, 
    37.03632, 37.05389, 37.07127, 37.08846, 37.10546, 37.12226, 37.13887, 
    37.15528, 37.1715, 37.18752, 37.20335, 37.21899, 37.23443, 37.24968, 
    37.26473, 37.27959, 37.29425, 37.30871, 37.32298, 37.33706, 37.35093, 
    37.36462, 37.3781, 37.39139, 37.40448, 37.41738, 37.43007, 37.44257, 
    37.45488, 37.46698, 37.47889, 37.4906, 37.50212, 37.51343, 37.52455, 
    37.53547, 37.54619, 37.55671, 37.56703, 37.57716, 37.58708, 37.59681, 
    37.60633, 37.61567, 37.62479, 37.63372, 37.64245, 37.65098, 37.65931, 
    37.66745, 37.67538, 37.68311, 37.69064, 37.69797, 37.7051, 37.71203, 
    37.71876, 37.72529, 37.73162, 37.73774, 37.74367, 37.7494, 37.75492, 
    37.76025, 37.76537, 37.77029, 37.77502, 37.77954, 37.78386, 37.78797, 
    37.79189, 37.7956, 37.79912, 37.80243, 37.80554, 37.80845, 37.81116, 
    37.81366, 37.81597, 37.81807, 37.81997, 37.82167, 37.82317, 37.82446, 
    37.82556, 37.82645, 37.82714, 37.82763, 37.82792, 37.828, 37.82788, 
    37.82756, 37.82704, 37.82632, 37.8254, 37.82427, 37.82294, 37.82141, 
    37.81968, 37.81775, 37.81562, 37.81328, 37.81074, 37.808, 37.80506, 
    37.80192, 37.79858, 37.79503, 37.79128, 37.78733, 37.78318, 37.77884, 
    37.77428, 37.76953, 37.76458, 37.75942, 37.75406, 37.7485, 37.74275, 
    37.73679, 37.73063, 37.72427, 37.71771, 37.71095, 37.70398, 37.69682, 
    37.68946, 37.6819, 37.67413, 37.66617, 37.65801, 37.64965, 37.64109, 
    37.63232, 37.62336, 37.6142, 37.60484, 37.59528, 37.58553, 37.57557, 
    37.56541, 37.55506, 37.54451, 37.53375, 37.5228, 37.51165, 37.50031, 
    37.48877, 37.47702, 37.46508, 37.45295, 37.44061, 37.42808, 37.41535, 
    37.40242, 37.3893, 37.37598, 37.36246, 37.34875, 37.33484, 37.32074, 
    37.30644, 37.29194, 37.27725, 37.26236, 37.24728, 37.232, 37.21653, 
    37.20086, 37.185, 37.16895, 37.15269, 37.13625, 37.11961, 37.10278, 
    37.08576, 37.06854, 37.05113, 37.03352, 37.01573, 36.99774, 36.97956, 
    36.96118, 36.94262, 36.92386, 36.90491, 36.88577, 36.86644, 36.84692, 
    36.82721, 36.80731, 36.78722, 36.76693, 36.74646, 36.7258, 36.70495, 
    36.68391, 36.66268, 36.64126, 36.61966, 36.59787, 36.57589, 36.55371, 
    36.53136, 36.50882, 36.48609, 36.46317, 36.44007, 36.41678, 36.3933, 
    36.36964, 36.34579, 36.32177, 36.29755, 36.27315, 36.24856, 36.22379, 
    36.19884, 36.1737, 36.14838, 36.12288, 36.09719, 36.07133, 36.04528, 
    36.01904, 35.99263, 35.96603, 35.93926, 35.9123, 35.88516, 35.85785, 
    35.83035, 35.80267, 35.77481, 35.74677, 35.71856, 35.69016, 35.66159, 
    35.63284, 35.60391, 35.57481, 35.54552, 35.51606, 35.48643, 35.45661, 
    35.42662, 35.39646, 35.36612, 35.33561, 35.30492, 35.27405, 35.24302, 
    35.2118, 35.18042, 35.14886, 35.11713, 35.08522, 35.05315, 35.0209, 
    34.98848, 34.95588,
  31.3277, 31.37481, 31.42179, 31.46863, 31.51533, 31.56189, 31.6083, 
    31.65458, 31.70071, 31.7467, 31.79255, 31.83825, 31.88381, 31.92923, 
    31.9745, 32.01963, 32.06461, 32.10945, 32.15414, 32.19869, 32.24309, 
    32.28734, 32.33145, 32.37541, 32.41922, 32.46289, 32.5064, 32.54977, 
    32.59298, 32.63605, 32.67897, 32.72174, 32.76436, 32.80682, 32.84914, 
    32.8913, 32.93332, 32.97518, 33.01688, 33.05844, 33.09984, 33.14109, 
    33.18218, 33.22312, 33.26391, 33.30453, 33.34501, 33.38533, 33.42549, 
    33.4655, 33.50535, 33.54504, 33.58458, 33.62395, 33.66317, 33.70224, 
    33.74114, 33.77988, 33.81846, 33.85689, 33.89515, 33.93325, 33.9712, 
    34.00898, 34.0466, 34.08406, 34.12135, 34.15849, 34.19545, 34.23226, 
    34.26891, 34.30539, 34.3417, 34.37785, 34.41384, 34.44966, 34.48531, 
    34.52081, 34.55613, 34.59129, 34.62627, 34.6611, 34.69576, 34.73024, 
    34.76456, 34.79871, 34.8327, 34.86651, 34.90015, 34.93363, 34.96693, 
    35.00006, 35.03303, 35.06582, 35.09844, 35.13089, 35.16317, 35.19527, 
    35.2272, 35.25896, 35.29055, 35.32196, 35.3532, 35.38427, 35.41515, 
    35.44587, 35.47641, 35.50677, 35.53696, 35.56698, 35.59682, 35.62648, 
    35.65596, 35.68526, 35.71439, 35.74335, 35.77212, 35.80072, 35.82913, 
    35.85737, 35.88543, 35.91331, 35.94101, 35.96852, 35.99586, 36.02302, 
    36.05, 36.07679, 36.10341, 36.12984, 36.15609, 36.18216, 36.20805, 
    36.23375, 36.25927, 36.28461, 36.30976, 36.33473, 36.35951, 36.38411, 
    36.40853, 36.43276, 36.45681, 36.48067, 36.50434, 36.52783, 36.55113, 
    36.57425, 36.59718, 36.61992, 36.64247, 36.66484, 36.68702, 36.70901, 
    36.73082, 36.75243, 36.77386, 36.79509, 36.81614, 36.837, 36.85767, 
    36.87815, 36.89844, 36.91854, 36.93845, 36.95817, 36.9777, 36.99703, 
    37.01617, 37.03513, 37.05389, 37.07246, 37.09084, 37.10902, 37.12701, 
    37.14481, 37.16242, 37.17983, 37.19705, 37.21408, 37.23091, 37.24755, 
    37.264, 37.28025, 37.2963, 37.31216, 37.32783, 37.3433, 37.35857, 
    37.37365, 37.38854, 37.40323, 37.41772, 37.43202, 37.44612, 37.46002, 
    37.47373, 37.48724, 37.50055, 37.51367, 37.52659, 37.53931, 37.55183, 
    37.56416, 37.57629, 37.58822, 37.59996, 37.61149, 37.62283, 37.63396, 
    37.64491, 37.65565, 37.66619, 37.67653, 37.68667, 37.69662, 37.70636, 
    37.71591, 37.72525, 37.7344, 37.74335, 37.75209, 37.76064, 37.76899, 
    37.77714, 37.78508, 37.79283, 37.80037, 37.80772, 37.81486, 37.8218, 
    37.82855, 37.83509, 37.84143, 37.84757, 37.85351, 37.85925, 37.86478, 
    37.87012, 37.87525, 37.88018, 37.88491, 37.88944, 37.89377, 37.8979, 
    37.90182, 37.90554, 37.90906, 37.91238, 37.9155, 37.91841, 37.92112, 
    37.92363, 37.92595, 37.92805, 37.92995, 37.93166, 37.93316, 37.93446, 
    37.93555, 37.93645, 37.93714, 37.93763, 37.93792, 37.938, 37.93788, 
    37.93756, 37.93704, 37.93632, 37.93539, 37.93427, 37.93293, 37.9314, 
    37.92967, 37.92773, 37.92559, 37.92325, 37.92071, 37.91796, 37.91502, 
    37.91187, 37.90852, 37.90496, 37.90121, 37.89725, 37.8931, 37.88874, 
    37.88418, 37.87942, 37.87445, 37.86929, 37.86392, 37.85835, 37.85258, 
    37.84661, 37.84044, 37.83407, 37.8275, 37.82072, 37.81375, 37.80657, 
    37.79919, 37.79161, 37.78384, 37.77586, 37.76768, 37.7593, 37.75072, 
    37.74195, 37.73297, 37.72379, 37.71441, 37.70483, 37.69506, 37.68508, 
    37.67491, 37.66453, 37.65396, 37.64319, 37.63222, 37.62105, 37.60968, 
    37.59811, 37.58635, 37.57439, 37.56223, 37.54987, 37.53731, 37.52456, 
    37.51161, 37.49846, 37.48512, 37.47157, 37.45784, 37.4439, 37.42977, 
    37.41544, 37.40092, 37.3862, 37.37128, 37.35617, 37.34086, 37.32536, 
    37.30967, 37.29377, 37.27769, 37.26141, 37.24493, 37.22826, 37.2114, 
    37.19434, 37.17709, 37.15965, 37.14201, 37.12418, 37.10616, 37.08794, 
    37.06953, 37.05093, 37.03214, 37.01316, 36.99398, 36.97462, 36.95506, 
    36.93531, 36.91537, 36.89524, 36.87492, 36.85442, 36.83371, 36.81282, 
    36.79175, 36.77048, 36.74902, 36.72738, 36.70554, 36.68353, 36.66132, 
    36.63892, 36.61633, 36.59356, 36.5706, 36.54746, 36.52412, 36.50061, 
    36.4769, 36.45301, 36.42894, 36.40468, 36.38023, 36.35561, 36.33079, 
    36.30579, 36.28061, 36.25525, 36.22969, 36.20396, 36.17805, 36.15195, 
    36.12567, 36.09921, 36.07257, 36.04574, 36.01874, 35.99155, 35.96418, 
    35.93663, 35.90891, 35.881, 35.85291, 35.82465, 35.7962, 35.76758, 
    35.73878, 35.7098, 35.68064, 35.65131, 35.6218, 35.59211, 35.56224, 
    35.5322, 35.50198, 35.47159, 35.44102, 35.41028, 35.37936, 35.34827, 
    35.31701, 35.28556, 35.25395, 35.22216, 35.1902, 35.15807, 35.12577, 
    35.09329, 35.06064,
  31.42647, 31.47366, 31.5207, 31.56761, 31.61438, 31.66101, 31.70749, 
    31.75384, 31.80004, 31.8461, 31.89202, 31.93779, 31.98342, 32.0289, 
    32.07425, 32.11944, 32.16449, 32.2094, 32.25416, 32.29878, 32.34325, 
    32.38757, 32.43174, 32.47577, 32.51965, 32.56338, 32.60696, 32.6504, 
    32.69368, 32.73682, 32.7798, 32.82264, 32.86533, 32.90786, 32.95024, 
    32.99247, 33.03455, 33.07648, 33.11825, 33.15987, 33.20134, 33.24265, 
    33.28381, 33.32482, 33.36567, 33.40636, 33.4469, 33.48729, 33.52751, 
    33.56758, 33.6075, 33.64725, 33.68686, 33.7263, 33.76558, 33.8047, 
    33.84367, 33.88248, 33.92112, 33.95961, 33.99794, 34.0361, 34.07411, 
    34.11195, 34.14963, 34.18715, 34.22451, 34.2617, 34.29874, 34.33561, 
    34.37231, 34.40885, 34.44523, 34.48144, 34.51749, 34.55337, 34.58908, 
    34.62463, 34.66002, 34.69523, 34.73028, 34.76516, 34.79988, 34.83442, 
    34.8688, 34.90301, 34.93705, 34.97092, 35.00462, 35.03815, 35.07151, 
    35.10471, 35.13773, 35.17057, 35.20325, 35.23576, 35.26809, 35.30025, 
    35.33224, 35.36405, 35.39569, 35.42716, 35.45845, 35.48957, 35.52052, 
    35.55128, 35.58188, 35.6123, 35.64254, 35.6726, 35.7025, 35.73221, 
    35.76174, 35.7911, 35.82028, 35.84929, 35.87811, 35.90675, 35.93522, 
    35.96351, 35.99162, 36.01955, 36.04729, 36.07486, 36.10225, 36.12946, 
    36.15648, 36.18333, 36.20999, 36.23647, 36.26276, 36.28888, 36.31482, 
    36.34056, 36.36613, 36.39151, 36.41671, 36.44172, 36.46655, 36.4912, 
    36.51566, 36.53994, 36.56402, 36.58793, 36.61164, 36.63518, 36.65852, 
    36.68168, 36.70465, 36.72744, 36.75003, 36.77244, 36.79466, 36.81669, 
    36.83854, 36.86019, 36.88166, 36.90293, 36.92402, 36.94492, 36.96563, 
    36.98615, 37.00647, 37.02661, 37.04655, 37.06631, 37.08587, 37.10524, 
    37.12442, 37.14341, 37.16221, 37.18081, 37.19923, 37.21745, 37.23547, 
    37.2533, 37.27094, 37.28839, 37.30564, 37.3227, 37.33957, 37.35623, 
    37.37271, 37.38899, 37.40508, 37.42097, 37.43666, 37.45216, 37.46746, 
    37.48257, 37.49749, 37.5122, 37.52672, 37.54105, 37.55518, 37.5691, 
    37.58284, 37.59637, 37.60971, 37.62286, 37.6358, 37.64854, 37.66109, 
    37.67344, 37.6856, 37.69755, 37.7093, 37.72086, 37.73222, 37.74338, 
    37.75434, 37.7651, 37.77567, 37.78603, 37.79619, 37.80615, 37.81592, 
    37.82548, 37.83485, 37.84401, 37.85297, 37.86174, 37.8703, 37.87866, 
    37.88683, 37.89479, 37.90255, 37.91011, 37.91747, 37.92463, 37.93158, 
    37.93834, 37.94489, 37.95124, 37.9574, 37.96334, 37.96909, 37.97464, 
    37.97999, 37.98513, 37.99007, 37.99481, 37.99935, 38.00368, 38.00782, 
    38.01175, 38.01548, 38.019, 38.02233, 38.02545, 38.02837, 38.03109, 
    38.03361, 38.03592, 38.03803, 38.03994, 38.04165, 38.04315, 38.04445, 
    38.04555, 38.04644, 38.04713, 38.04763, 38.04791, 38.048, 38.04788, 
    38.04756, 38.04704, 38.04631, 38.04539, 38.04426, 38.04292, 38.04139, 
    38.03965, 38.03771, 38.03557, 38.03322, 38.03067, 38.02792, 38.02497, 
    38.02182, 38.01846, 38.0149, 38.01114, 38.00718, 38.00301, 37.99865, 
    37.99408, 37.9893, 37.98433, 37.97915, 37.97378, 37.9682, 37.96242, 
    37.95644, 37.95025, 37.94387, 37.93728, 37.9305, 37.92351, 37.91632, 
    37.90892, 37.90133, 37.89354, 37.88555, 37.87735, 37.86896, 37.86036, 
    37.85157, 37.84258, 37.83338, 37.82398, 37.81438, 37.80459, 37.79459, 
    37.7844, 37.77401, 37.76341, 37.75262, 37.74163, 37.73044, 37.71905, 
    37.70746, 37.69567, 37.68369, 37.6715, 37.65912, 37.64654, 37.63377, 
    37.62079, 37.60762, 37.59425, 37.58068, 37.56691, 37.55295, 37.5388, 
    37.52444, 37.50989, 37.49514, 37.4802, 37.46506, 37.44972, 37.43419, 
    37.41846, 37.40254, 37.38643, 37.37012, 37.35361, 37.33691, 37.32001, 
    37.30293, 37.28564, 37.26817, 37.2505, 37.23263, 37.21458, 37.19633, 
    37.17788, 37.15925, 37.14042, 37.1214, 37.10219, 37.08279, 37.0632, 
    37.04341, 37.02343, 37.00327, 36.98291, 36.96236, 36.94162, 36.9207, 
    36.89958, 36.87827, 36.85678, 36.83509, 36.81322, 36.79116, 36.76891, 
    36.74647, 36.72384, 36.70103, 36.67803, 36.65484, 36.63147, 36.60791, 
    36.58416, 36.56023, 36.53611, 36.5118, 36.48731, 36.46264, 36.43778, 
    36.41273, 36.38751, 36.3621, 36.3365, 36.31072, 36.28476, 36.25862, 
    36.23229, 36.20578, 36.17909, 36.15222, 36.12516, 36.09793, 36.07051, 
    36.04292, 36.01514, 35.98718, 35.95905, 35.93073, 35.90223, 35.87356, 
    35.84471, 35.81568, 35.78647, 35.75708, 35.72752, 35.69778, 35.66786, 
    35.63777, 35.6075, 35.57705, 35.54643, 35.51563, 35.48466, 35.45351, 
    35.42219, 35.3907, 35.35903, 35.32719, 35.29517, 35.26299, 35.23063, 
    35.19809, 35.16539,
  31.52521, 31.57247, 31.61959, 31.66657, 31.71341, 31.76011, 31.80666, 
    31.85307, 31.89935, 31.94547, 31.99146, 32.0373, 32.083, 32.12856, 
    32.17397, 32.21923, 32.26435, 32.30933, 32.35416, 32.39884, 32.44338, 
    32.48777, 32.53201, 32.57611, 32.62006, 32.66386, 32.7075, 32.75101, 
    32.79436, 32.83756, 32.88062, 32.92352, 32.96627, 33.00887, 33.05132, 
    33.09362, 33.13577, 33.17776, 33.2196, 33.26128, 33.30282, 33.3442, 
    33.38542, 33.42649, 33.46741, 33.50817, 33.54877, 33.58922, 33.62951, 
    33.66965, 33.70963, 33.74945, 33.78911, 33.82862, 33.86797, 33.90715, 
    33.94619, 33.98505, 34.02377, 34.06231, 34.1007, 34.13893, 34.177, 
    34.2149, 34.25265, 34.29023, 34.32765, 34.36491, 34.402, 34.43893, 
    34.4757, 34.5123, 34.54874, 34.58501, 34.62112, 34.65705, 34.69283, 
    34.72844, 34.76389, 34.79916, 34.83427, 34.86921, 34.90398, 34.93859, 
    34.97303, 35.00729, 35.04139, 35.07532, 35.10908, 35.14267, 35.17609, 
    35.20933, 35.24241, 35.27531, 35.30805, 35.34061, 35.373, 35.40521, 
    35.43726, 35.46913, 35.50082, 35.53234, 35.56369, 35.59486, 35.62586, 
    35.65668, 35.68733, 35.7178, 35.7481, 35.77822, 35.80816, 35.83792, 
    35.86752, 35.89692, 35.92616, 35.95521, 35.98409, 36.01278, 36.0413, 
    36.06964, 36.0978, 36.12577, 36.15357, 36.18119, 36.20863, 36.23588, 
    36.26295, 36.28985, 36.31656, 36.34309, 36.36943, 36.39559, 36.42157, 
    36.44737, 36.47298, 36.49841, 36.52365, 36.54871, 36.57359, 36.59828, 
    36.62278, 36.6471, 36.67123, 36.69518, 36.71894, 36.74252, 36.7659, 
    36.7891, 36.81212, 36.83494, 36.85758, 36.88003, 36.90229, 36.92437, 
    36.94625, 36.96795, 36.98945, 37.01077, 37.03189, 37.05283, 37.07357, 
    37.09413, 37.11449, 37.13467, 37.15465, 37.17444, 37.19404, 37.21345, 
    37.23267, 37.25169, 37.27052, 37.28916, 37.30761, 37.32586, 37.34392, 
    37.36179, 37.37946, 37.39694, 37.41422, 37.43131, 37.44821, 37.46491, 
    37.48142, 37.49773, 37.51384, 37.52977, 37.54549, 37.56102, 37.57635, 
    37.59149, 37.60643, 37.62118, 37.63572, 37.65007, 37.66423, 37.67818, 
    37.69194, 37.70551, 37.71887, 37.73204, 37.74501, 37.75778, 37.77035, 
    37.78272, 37.7949, 37.80688, 37.81865, 37.83023, 37.84161, 37.85279, 
    37.86377, 37.87456, 37.88514, 37.89552, 37.9057, 37.91569, 37.92547, 
    37.93505, 37.94444, 37.95362, 37.9626, 37.97138, 37.97996, 37.98833, 
    37.99651, 38.00449, 38.01227, 38.01984, 38.02721, 38.03439, 38.04136, 
    38.04813, 38.05469, 38.06106, 38.06722, 38.07318, 38.07894, 38.0845, 
    38.08986, 38.09501, 38.09996, 38.10471, 38.10925, 38.1136, 38.11774, 
    38.12168, 38.12542, 38.12895, 38.13228, 38.13541, 38.13834, 38.14106, 
    38.14358, 38.1459, 38.14801, 38.14993, 38.15163, 38.15314, 38.15444, 
    38.15554, 38.15644, 38.15714, 38.15763, 38.15791, 38.158, 38.15788, 
    38.15756, 38.15704, 38.15631, 38.15538, 38.15425, 38.15292, 38.15137, 
    38.14964, 38.14769, 38.14554, 38.1432, 38.14064, 38.13789, 38.13493, 
    38.13177, 38.1284, 38.12484, 38.12107, 38.1171, 38.11293, 38.10855, 
    38.10397, 38.09919, 38.09421, 38.08902, 38.08363, 38.07804, 38.07225, 
    38.06626, 38.06006, 38.05367, 38.04707, 38.04027, 38.03326, 38.02606, 
    38.01866, 38.01105, 38.00324, 37.99524, 37.98702, 37.97861, 37.97, 
    37.96119, 37.95218, 37.94296, 37.93355, 37.92393, 37.91412, 37.90411, 
    37.89389, 37.88348, 37.87286, 37.86205, 37.85104, 37.83982, 37.82841, 
    37.8168, 37.805, 37.79299, 37.78078, 37.76838, 37.75577, 37.74297, 
    37.72997, 37.71677, 37.70338, 37.68978, 37.67599, 37.662, 37.64782, 
    37.63343, 37.61886, 37.60408, 37.58911, 37.57394, 37.55858, 37.54302, 
    37.52726, 37.51131, 37.49516, 37.47882, 37.46228, 37.44555, 37.42862, 
    37.4115, 37.39419, 37.37668, 37.35897, 37.34108, 37.32299, 37.3047, 
    37.28623, 37.26756, 37.2487, 37.22964, 37.2104, 37.19096, 37.17133, 
    37.1515, 37.13149, 37.11129, 37.09089, 37.0703, 37.04953, 37.02856, 
    37.00741, 36.98606, 36.96452, 36.9428, 36.92089, 36.89878, 36.87649, 
    36.85401, 36.83134, 36.80849, 36.78545, 36.76222, 36.7388, 36.71519, 
    36.69141, 36.66743, 36.64326, 36.61892, 36.59438, 36.56966, 36.54476, 
    36.51967, 36.4944, 36.46894, 36.4433, 36.41748, 36.39147, 36.36528, 
    36.3389, 36.31234, 36.28561, 36.25869, 36.23158, 36.2043, 36.17683, 
    36.14919, 36.12136, 36.09335, 36.06517, 36.0368, 36.00826, 35.97953, 
    35.95063, 35.92154, 35.89228, 35.86285, 35.83323, 35.80344, 35.77347, 
    35.74332, 35.713, 35.6825, 35.65182, 35.62097, 35.58995, 35.55875, 
    35.52737, 35.49582, 35.4641, 35.4322, 35.40013, 35.36789, 35.33547, 
    35.30288, 35.27012,
  31.62393, 31.67126, 31.71845, 31.7655, 31.81241, 31.85917, 31.9058, 
    31.95228, 31.99862, 32.04482, 32.09088, 32.13679, 32.18256, 32.22818, 
    32.27366, 32.319, 32.36419, 32.40923, 32.45413, 32.49888, 32.54349, 
    32.58795, 32.63226, 32.67642, 32.72044, 32.76431, 32.80803, 32.85159, 
    32.89502, 32.93829, 32.98141, 33.02438, 33.0672, 33.10986, 33.15238, 
    33.19474, 33.23695, 33.27901, 33.32092, 33.36267, 33.40427, 33.44572, 
    33.48701, 33.52814, 33.56913, 33.60995, 33.65062, 33.69114, 33.73149, 
    33.77169, 33.81174, 33.85162, 33.89135, 33.93092, 33.97033, 34.00959, 
    34.04868, 34.08761, 34.12638, 34.165, 34.20345, 34.24174, 34.27987, 
    34.31784, 34.35565, 34.3933, 34.43077, 34.46809, 34.50525, 34.54224, 
    34.57907, 34.61573, 34.65223, 34.68856, 34.72473, 34.76073, 34.79657, 
    34.83224, 34.86774, 34.90307, 34.93824, 34.97324, 35.00808, 35.04274, 
    35.07723, 35.11156, 35.14572, 35.1797, 35.21352, 35.24717, 35.28064, 
    35.31395, 35.34708, 35.38004, 35.41283, 35.44545, 35.47789, 35.51017, 
    35.54226, 35.57419, 35.60594, 35.63752, 35.66892, 35.70015, 35.7312, 
    35.76207, 35.79278, 35.8233, 35.85365, 35.88382, 35.91382, 35.94363, 
    35.97327, 36.00274, 36.03202, 36.06113, 36.09005, 36.1188, 36.14737, 
    36.17575, 36.20396, 36.23199, 36.25984, 36.28751, 36.31499, 36.3423, 
    36.36942, 36.39636, 36.42312, 36.44969, 36.47609, 36.5023, 36.52832, 
    36.55416, 36.57982, 36.6053, 36.63059, 36.65569, 36.68061, 36.70535, 
    36.7299, 36.75426, 36.77844, 36.80243, 36.82623, 36.84985, 36.87328, 
    36.89652, 36.91958, 36.94244, 36.96513, 36.98762, 37.00992, 37.03203, 
    37.05396, 37.07569, 37.09724, 37.11859, 37.13976, 37.16073, 37.18152, 
    37.20211, 37.22252, 37.24273, 37.26274, 37.28257, 37.30221, 37.32166, 
    37.34091, 37.35997, 37.37883, 37.39751, 37.41599, 37.43428, 37.45237, 
    37.47027, 37.48798, 37.50549, 37.5228, 37.53992, 37.55685, 37.57359, 
    37.59012, 37.60646, 37.62261, 37.63856, 37.65432, 37.66988, 37.68524, 
    37.70041, 37.71537, 37.73014, 37.74472, 37.7591, 37.77328, 37.78727, 
    37.80105, 37.81464, 37.82803, 37.84122, 37.85421, 37.86701, 37.8796, 
    37.892, 37.9042, 37.9162, 37.928, 37.9396, 37.951, 37.9622, 37.97321, 
    37.98401, 37.99461, 38.00502, 38.01522, 38.02522, 38.03502, 38.04462, 
    38.05402, 38.06322, 38.07222, 38.08102, 38.08961, 38.09801, 38.1062, 
    38.11419, 38.12199, 38.12957, 38.13696, 38.14415, 38.15113, 38.15791, 
    38.16449, 38.17087, 38.17704, 38.18302, 38.18879, 38.19436, 38.19972, 
    38.20489, 38.20985, 38.2146, 38.21916, 38.22351, 38.22766, 38.23161, 
    38.23535, 38.2389, 38.24223, 38.24537, 38.2483, 38.25103, 38.25355, 
    38.25587, 38.25799, 38.25991, 38.26162, 38.26313, 38.26443, 38.26554, 
    38.26644, 38.26713, 38.26762, 38.26791, 38.268, 38.26788, 38.26756, 
    38.26704, 38.26631, 38.26538, 38.26424, 38.26291, 38.26136, 38.25962, 
    38.25767, 38.25552, 38.25317, 38.25061, 38.24785, 38.24488, 38.24172, 
    38.23835, 38.23478, 38.231, 38.22702, 38.22284, 38.21845, 38.21387, 
    38.20908, 38.20408, 38.19889, 38.19349, 38.18789, 38.18209, 38.17608, 
    38.16988, 38.16346, 38.15685, 38.15004, 38.14302, 38.13581, 38.12839, 
    38.12077, 38.11294, 38.10492, 38.09669, 38.08827, 38.07964, 38.07081, 
    38.06178, 38.05255, 38.04312, 38.03349, 38.02365, 38.01362, 38.00338, 
    37.99295, 37.98232, 37.97148, 37.96045, 37.94921, 37.93778, 37.92615, 
    37.91431, 37.90228, 37.89005, 37.87762, 37.865, 37.85217, 37.83915, 
    37.82592, 37.8125, 37.79888, 37.78506, 37.77105, 37.75684, 37.74243, 
    37.72782, 37.71302, 37.69802, 37.68282, 37.66743, 37.65184, 37.63605, 
    37.62007, 37.60389, 37.58752, 37.57095, 37.55419, 37.53723, 37.52008, 
    37.50273, 37.48519, 37.46745, 37.44952, 37.4314, 37.41308, 37.39457, 
    37.37586, 37.35696, 37.33788, 37.31859, 37.29912, 37.27945, 37.25959, 
    37.23954, 37.2193, 37.19887, 37.17824, 37.15743, 37.13642, 37.11523, 
    37.09384, 37.07227, 37.0505, 37.02855, 37.0064, 36.98407, 36.96155, 
    36.93884, 36.91594, 36.89286, 36.86959, 36.84613, 36.82248, 36.79865, 
    36.77462, 36.75042, 36.72602, 36.70145, 36.67668, 36.65173, 36.6266, 
    36.60128, 36.57578, 36.55009, 36.52422, 36.49816, 36.47192, 36.4455, 
    36.4189, 36.39211, 36.36514, 36.33799, 36.31066, 36.28314, 36.25545, 
    36.22757, 36.19951, 36.17128, 36.14286, 36.11427, 36.08549, 36.05653, 
    36.0274, 35.99809, 35.9686, 35.93893, 35.90908, 35.87906, 35.84886, 
    35.81849, 35.78793, 35.7572, 35.7263, 35.69522, 35.66396, 35.63253, 
    35.60093, 35.56915, 35.5372, 35.50507, 35.47277, 35.4403, 35.40766, 
    35.37484,
  31.72263, 31.77003, 31.81729, 31.86441, 31.91138, 31.95822, 32.00492, 
    32.05147, 32.09788, 32.14415, 32.19027, 32.23626, 32.28209, 32.32779, 
    32.37334, 32.41874, 32.464, 32.50911, 32.55408, 32.5989, 32.64358, 
    32.6881, 32.73248, 32.77671, 32.8208, 32.86473, 32.90852, 32.95216, 
    32.99565, 33.03899, 33.08217, 33.12521, 33.1681, 33.21083, 33.25341, 
    33.29585, 33.33812, 33.38025, 33.42223, 33.46404, 33.50571, 33.54722, 
    33.58858, 33.62978, 33.67083, 33.71172, 33.75245, 33.79303, 33.83345, 
    33.87372, 33.91383, 33.95378, 33.99357, 34.03321, 34.07268, 34.112, 
    34.15116, 34.19016, 34.22899, 34.26767, 34.30618, 34.34454, 34.38273, 
    34.42076, 34.45863, 34.49634, 34.53388, 34.57126, 34.60848, 34.64553, 
    34.68242, 34.71914, 34.7557, 34.7921, 34.82833, 34.86439, 34.90028, 
    34.93601, 34.97158, 35.00697, 35.0422, 35.07726, 35.11215, 35.14687, 
    35.18143, 35.21581, 35.25003, 35.28407, 35.31795, 35.35165, 35.38519, 
    35.41854, 35.45174, 35.48475, 35.5176, 35.55027, 35.58278, 35.6151, 
    35.64726, 35.67924, 35.71104, 35.74268, 35.77413, 35.80542, 35.83652, 
    35.86745, 35.89821, 35.92879, 35.95919, 35.98941, 36.01946, 36.04933, 
    36.07902, 36.10854, 36.13787, 36.16703, 36.19601, 36.2248, 36.25343, 
    36.28186, 36.31012, 36.3382, 36.3661, 36.39381, 36.42135, 36.4487, 
    36.47587, 36.50286, 36.52967, 36.55629, 36.58273, 36.60899, 36.63506, 
    36.66095, 36.68666, 36.71218, 36.73751, 36.76266, 36.78763, 36.81241, 
    36.837, 36.86141, 36.88563, 36.90967, 36.93351, 36.95718, 36.98065, 
    37.00393, 37.02703, 37.04994, 37.07266, 37.0952, 37.11754, 37.13969, 
    37.16166, 37.18343, 37.20502, 37.22641, 37.24762, 37.26863, 37.28946, 
    37.31009, 37.33053, 37.35078, 37.37083, 37.3907, 37.41037, 37.42985, 
    37.44914, 37.46824, 37.48714, 37.50585, 37.52436, 37.54268, 37.56081, 
    37.57874, 37.59649, 37.61403, 37.63138, 37.64853, 37.66549, 37.68225, 
    37.69883, 37.7152, 37.73138, 37.74736, 37.76314, 37.77873, 37.79412, 
    37.80931, 37.82431, 37.83911, 37.85372, 37.86812, 37.88233, 37.89634, 
    37.91015, 37.92376, 37.93718, 37.9504, 37.96342, 37.97623, 37.98886, 
    38.00128, 38.0135, 38.02552, 38.03735, 38.04897, 38.06039, 38.07161, 
    38.08264, 38.09346, 38.10408, 38.11451, 38.12473, 38.13475, 38.14457, 
    38.15419, 38.16361, 38.17282, 38.18184, 38.19065, 38.19927, 38.20768, 
    38.21589, 38.2239, 38.2317, 38.23931, 38.24671, 38.25391, 38.2609, 
    38.2677, 38.27429, 38.28068, 38.28687, 38.29285, 38.29863, 38.30421, 
    38.30959, 38.31476, 38.31973, 38.3245, 38.32906, 38.33343, 38.33759, 
    38.34154, 38.34529, 38.34884, 38.35218, 38.35532, 38.35826, 38.36099, 
    38.36352, 38.36585, 38.36797, 38.36989, 38.37161, 38.37312, 38.37443, 
    38.37553, 38.37643, 38.37713, 38.37762, 38.37791, 38.378, 38.37788, 
    38.37756, 38.37703, 38.3763, 38.37537, 38.37423, 38.37289, 38.37135, 
    38.3696, 38.36765, 38.36549, 38.36314, 38.36057, 38.35781, 38.35484, 
    38.35167, 38.34829, 38.34471, 38.34093, 38.33694, 38.33275, 38.32836, 
    38.32376, 38.31896, 38.31396, 38.30875, 38.30334, 38.29773, 38.29192, 
    38.2859, 38.27969, 38.27326, 38.26664, 38.25981, 38.25278, 38.24555, 
    38.23812, 38.23048, 38.22264, 38.2146, 38.20636, 38.19792, 38.18927, 
    38.18043, 38.17138, 38.16213, 38.15268, 38.14303, 38.13318, 38.12313, 
    38.11287, 38.10242, 38.09176, 38.08091, 38.06985, 38.0586, 38.04714, 
    38.03549, 38.02363, 38.01158, 37.99932, 37.98687, 37.97422, 37.96137, 
    37.94832, 37.93507, 37.92162, 37.90798, 37.89414, 37.8801, 37.86586, 
    37.85142, 37.83678, 37.82195, 37.80692, 37.7917, 37.77628, 37.76066, 
    37.74484, 37.72883, 37.71262, 37.69622, 37.67962, 37.66282, 37.64583, 
    37.62865, 37.61127, 37.59369, 37.57592, 37.55796, 37.5398, 37.52145, 
    37.5029, 37.48416, 37.46523, 37.4461, 37.42678, 37.40727, 37.38757, 
    37.36767, 37.34758, 37.3273, 37.30684, 37.28617, 37.26532, 37.24427, 
    37.22304, 37.20161, 37.18, 37.1582, 37.1362, 37.11402, 37.09164, 
    37.06908, 37.04633, 37.02339, 37.00026, 36.97695, 36.95345, 36.92975, 
    36.90588, 36.88181, 36.85756, 36.83312, 36.8085, 36.78369, 36.7587, 
    36.73352, 36.70815, 36.6826, 36.65687, 36.63095, 36.60485, 36.57856, 
    36.55209, 36.52544, 36.4986, 36.47159, 36.44439, 36.417, 36.38944, 
    36.3617, 36.33377, 36.30566, 36.27738, 36.24891, 36.22026, 36.19144, 
    36.16243, 36.13324, 36.10388, 36.07434, 36.04462, 36.01472, 35.98464, 
    35.95439, 35.92396, 35.89335, 35.86257, 35.83161, 35.80048, 35.76917, 
    35.73768, 35.70602, 35.67419, 35.64218, 35.61, 35.57764, 35.54512, 
    35.51242, 35.47954,
  31.8213, 31.86877, 31.9161, 31.96329, 32.01033, 32.05724, 32.10401, 
    32.15063, 32.19711, 32.24345, 32.28965, 32.3357, 32.3816, 32.42737, 
    32.47298, 32.51846, 32.56379, 32.60897, 32.65401, 32.6989, 32.74364, 
    32.78823, 32.83268, 32.87698, 32.92114, 32.96514, 33.009, 33.0527, 
    33.09626, 33.13966, 33.18292, 33.22602, 33.26898, 33.31178, 33.35443, 
    33.39693, 33.43927, 33.48147, 33.52351, 33.56539, 33.60712, 33.6487, 
    33.69012, 33.73139, 33.77251, 33.81347, 33.85426, 33.89491, 33.9354, 
    33.97573, 34.0159, 34.05592, 34.09577, 34.13547, 34.17501, 34.21439, 
    34.25361, 34.29268, 34.33158, 34.37032, 34.40889, 34.44731, 34.48557, 
    34.52366, 34.5616, 34.59937, 34.63697, 34.67441, 34.71169, 34.74881, 
    34.78576, 34.82254, 34.85916, 34.89562, 34.93191, 34.96803, 35.00399, 
    35.03978, 35.0754, 35.11086, 35.14614, 35.18126, 35.21621, 35.25099, 
    35.28561, 35.32005, 35.35432, 35.38842, 35.42236, 35.45612, 35.48971, 
    35.52313, 35.55638, 35.58945, 35.62236, 35.65509, 35.68764, 35.72003, 
    35.75224, 35.78427, 35.81614, 35.84782, 35.87933, 35.91067, 35.94183, 
    35.97282, 36.00362, 36.03426, 36.06471, 36.09499, 36.12509, 36.15501, 
    36.18476, 36.21432, 36.24371, 36.27292, 36.30195, 36.3308, 36.35947, 
    36.38796, 36.41627, 36.4444, 36.47234, 36.50011, 36.52769, 36.5551, 
    36.58232, 36.60936, 36.63621, 36.66288, 36.68937, 36.71567, 36.74179, 
    36.76773, 36.79348, 36.81905, 36.84443, 36.86963, 36.89464, 36.91946, 
    36.9441, 36.96855, 36.99282, 37.0169, 37.04079, 37.06449, 37.08801, 
    37.11134, 37.13448, 37.15743, 37.18019, 37.20277, 37.22515, 37.24734, 
    37.26935, 37.29116, 37.31279, 37.33422, 37.35547, 37.37652, 37.39738, 
    37.41806, 37.43853, 37.45882, 37.47892, 37.49882, 37.51853, 37.53804, 
    37.55737, 37.5765, 37.59544, 37.61418, 37.63273, 37.65109, 37.66925, 
    37.68722, 37.70499, 37.72256, 37.73995, 37.75714, 37.77413, 37.79092, 
    37.80752, 37.82393, 37.84013, 37.85615, 37.87196, 37.88758, 37.903, 
    37.91822, 37.93325, 37.94808, 37.96271, 37.97714, 37.99137, 38.00541, 
    38.01925, 38.03289, 38.04633, 38.05957, 38.07262, 38.08546, 38.09811, 
    38.11055, 38.1228, 38.13484, 38.14669, 38.15833, 38.16978, 38.18102, 
    38.19207, 38.20291, 38.21355, 38.224, 38.23424, 38.24428, 38.25412, 
    38.26376, 38.27319, 38.28243, 38.29146, 38.30029, 38.30892, 38.31735, 
    38.32557, 38.3336, 38.34142, 38.34904, 38.35645, 38.36367, 38.37068, 
    38.37748, 38.38409, 38.39049, 38.39669, 38.40269, 38.40848, 38.41407, 
    38.41946, 38.42464, 38.42962, 38.4344, 38.43897, 38.44334, 38.44751, 
    38.45147, 38.45523, 38.45878, 38.46213, 38.46528, 38.46822, 38.47096, 
    38.4735, 38.47583, 38.47795, 38.47988, 38.48159, 38.48311, 38.48442, 
    38.48553, 38.48643, 38.48713, 38.48763, 38.48792, 38.488, 38.48788, 
    38.48756, 38.48703, 38.4863, 38.48537, 38.48423, 38.48288, 38.48134, 
    38.47959, 38.47763, 38.47547, 38.47311, 38.47054, 38.46777, 38.46479, 
    38.46162, 38.45823, 38.45464, 38.45086, 38.44686, 38.44266, 38.43826, 
    38.43365, 38.42885, 38.42384, 38.41862, 38.4132, 38.40758, 38.40175, 
    38.39573, 38.38949, 38.38306, 38.37642, 38.36958, 38.36254, 38.35529, 
    38.34785, 38.34019, 38.33234, 38.32429, 38.31603, 38.30757, 38.29891, 
    38.29005, 38.28098, 38.27171, 38.26225, 38.25257, 38.24271, 38.23263, 
    38.22236, 38.21188, 38.20121, 38.19033, 38.17926, 38.16798, 38.1565, 
    38.14482, 38.13295, 38.12087, 38.10859, 38.09612, 38.08344, 38.07057, 
    38.05749, 38.04422, 38.03075, 38.01707, 38.0032, 37.98914, 37.97487, 
    37.96041, 37.94574, 37.93089, 37.91583, 37.90057, 37.88512, 37.86947, 
    37.85363, 37.83759, 37.82135, 37.80491, 37.78828, 37.77145, 37.75443, 
    37.73721, 37.7198, 37.70219, 37.68439, 37.66639, 37.6482, 37.62981, 
    37.61123, 37.59246, 37.57349, 37.55433, 37.53497, 37.51542, 37.49568, 
    37.47575, 37.45562, 37.43531, 37.4148, 37.3941, 37.37321, 37.35212, 
    37.33085, 37.30938, 37.28773, 37.26588, 37.24385, 37.22162, 37.19921, 
    37.17661, 37.15381, 37.13083, 37.10766, 37.0843, 37.06076, 37.03702, 
    37.0131, 36.98899, 36.96469, 36.94022, 36.91555, 36.89069, 36.86565, 
    36.84043, 36.81501, 36.78942, 36.76364, 36.73767, 36.71152, 36.68519, 
    36.65867, 36.63197, 36.60509, 36.57802, 36.55077, 36.52334, 36.49573, 
    36.46794, 36.43996, 36.4118, 36.38346, 36.35495, 36.32625, 36.29737, 
    36.26831, 36.23907, 36.20966, 36.18007, 36.15029, 36.12034, 36.09021, 
    36.05991, 36.02942, 35.99876, 35.96793, 35.93691, 35.90572, 35.87436, 
    35.84282, 35.81111, 35.77922, 35.74715, 35.71492, 35.68251, 35.64992, 
    35.61716, 35.58423,
  31.91994, 31.96748, 32.01488, 32.06214, 32.10926, 32.15624, 32.20308, 
    32.24977, 32.29632, 32.34273, 32.38899, 32.43511, 32.48109, 32.52692, 
    32.57261, 32.61815, 32.66355, 32.70881, 32.75391, 32.79887, 32.84368, 
    32.88834, 32.93286, 32.97723, 33.02145, 33.06553, 33.10945, 33.15322, 
    33.19685, 33.24032, 33.28364, 33.32681, 33.36983, 33.4127, 33.45542, 
    33.49799, 33.5404, 33.58266, 33.62477, 33.66672, 33.70852, 33.75016, 
    33.79165, 33.83298, 33.87416, 33.91519, 33.95605, 33.99677, 34.03732, 
    34.07771, 34.11795, 34.15803, 34.19796, 34.23772, 34.27732, 34.31677, 
    34.35605, 34.39518, 34.43414, 34.47295, 34.51159, 34.55007, 34.58839, 
    34.62654, 34.66454, 34.70237, 34.74004, 34.77755, 34.81489, 34.85206, 
    34.88908, 34.92592, 34.9626, 34.99912, 35.03547, 35.07166, 35.10767, 
    35.14352, 35.1792, 35.21472, 35.25006, 35.28524, 35.32026, 35.35509, 
    35.38977, 35.42427, 35.4586, 35.49276, 35.52675, 35.56057, 35.59422, 
    35.6277, 35.661, 35.69414, 35.7271, 35.75988, 35.7925, 35.82494, 35.8572, 
    35.88929, 35.92121, 35.95295, 35.98452, 36.01591, 36.04713, 36.07817, 
    36.10903, 36.13972, 36.17023, 36.20056, 36.23071, 36.26068, 36.29049, 
    36.3201, 36.34954, 36.3788, 36.40788, 36.43679, 36.46551, 36.49405, 
    36.52241, 36.55058, 36.57858, 36.6064, 36.63403, 36.66148, 36.68875, 
    36.71584, 36.74274, 36.76946, 36.79599, 36.82235, 36.84851, 36.8745, 
    36.9003, 36.92591, 36.95134, 36.97658, 37.00164, 37.0265, 37.05119, 
    37.07569, 37.09999, 37.12412, 37.14806, 37.1718, 37.19536, 37.21873, 
    37.24192, 37.26491, 37.28772, 37.31033, 37.33276, 37.35499, 37.37704, 
    37.3989, 37.42056, 37.44203, 37.46332, 37.48441, 37.50531, 37.52602, 
    37.54654, 37.56686, 37.58699, 37.60693, 37.62668, 37.64623, 37.66559, 
    37.68476, 37.70373, 37.72251, 37.7411, 37.75949, 37.77768, 37.79568, 
    37.81349, 37.8311, 37.84851, 37.86573, 37.88276, 37.89959, 37.91622, 
    37.93265, 37.94889, 37.96493, 37.98078, 37.99643, 38.01188, 38.02713, 
    38.04218, 38.05704, 38.0717, 38.08615, 38.10042, 38.11448, 38.12835, 
    38.14201, 38.15548, 38.16875, 38.18182, 38.19468, 38.20735, 38.21982, 
    38.23209, 38.24416, 38.25603, 38.2677, 38.27916, 38.29043, 38.30149, 
    38.31236, 38.32302, 38.33348, 38.34375, 38.35381, 38.36367, 38.37332, 
    38.38278, 38.39203, 38.40108, 38.40993, 38.41858, 38.42702, 38.43526, 
    38.4433, 38.45113, 38.45877, 38.4662, 38.47342, 38.48045, 38.48727, 
    38.49389, 38.5003, 38.50652, 38.51252, 38.51833, 38.52393, 38.52932, 
    38.53452, 38.53951, 38.54429, 38.54887, 38.55325, 38.55743, 38.5614, 
    38.56516, 38.56872, 38.57208, 38.57523, 38.57818, 38.58093, 38.58347, 
    38.5858, 38.58793, 38.58986, 38.59158, 38.5931, 38.59441, 38.59552, 
    38.59643, 38.59713, 38.59762, 38.59791, 38.598, 38.59788, 38.59756, 
    38.59703, 38.5963, 38.59536, 38.59422, 38.59288, 38.59132, 38.58957, 
    38.58761, 38.58545, 38.58308, 38.58051, 38.57773, 38.57475, 38.57156, 
    38.56817, 38.56458, 38.56078, 38.55678, 38.55257, 38.54816, 38.54355, 
    38.53873, 38.53371, 38.52848, 38.52306, 38.51742, 38.51159, 38.50555, 
    38.4993, 38.49286, 38.48621, 38.47935, 38.47229, 38.46503, 38.45757, 
    38.44991, 38.44204, 38.43397, 38.4257, 38.41722, 38.40854, 38.39966, 
    38.39058, 38.38129, 38.37181, 38.36212, 38.35223, 38.34214, 38.33184, 
    38.32135, 38.31065, 38.29976, 38.28866, 38.27736, 38.26586, 38.25416, 
    38.24226, 38.23016, 38.21786, 38.20536, 38.19266, 38.17976, 38.16666, 
    38.15336, 38.13987, 38.12617, 38.11227, 38.09818, 38.08388, 38.06939, 
    38.0547, 38.03981, 38.02473, 38.00944, 37.99396, 37.97828, 37.96241, 
    37.94633, 37.93007, 37.9136, 37.89694, 37.88008, 37.86302, 37.84577, 
    37.82833, 37.81068, 37.79285, 37.77482, 37.75659, 37.73817, 37.71955, 
    37.70074, 37.68174, 37.66254, 37.64315, 37.62357, 37.60379, 37.58382, 
    37.56366, 37.5433, 37.52275, 37.50201, 37.48109, 37.45996, 37.43865, 
    37.41714, 37.39545, 37.37356, 37.35149, 37.32922, 37.30677, 37.28412, 
    37.26128, 37.23826, 37.21505, 37.19165, 37.16806, 37.14428, 37.12032, 
    37.09616, 37.07182, 37.0473, 37.02258, 36.99768, 36.9726, 36.94733, 
    36.92187, 36.89623, 36.8704, 36.84439, 36.81819, 36.79181, 36.76524, 
    36.73849, 36.71156, 36.68445, 36.65715, 36.62967, 36.60201, 36.57417, 
    36.54614, 36.51793, 36.48954, 36.46098, 36.43222, 36.4033, 36.37419, 
    36.3449, 36.31543, 36.28578, 36.25596, 36.22595, 36.19577, 36.16541, 
    36.13488, 36.10416, 36.07327, 36.0422, 36.01096, 35.97954, 35.94794, 
    35.91618, 35.88423, 35.85211, 35.81982, 35.78735, 35.75471, 35.72189, 
    35.68891,
  32.01856, 32.06617, 32.11364, 32.16097, 32.20816, 32.25521, 32.30212, 
    32.34888, 32.3955, 32.44198, 32.48832, 32.5345, 32.58055, 32.62645, 
    32.67221, 32.71782, 32.76329, 32.80861, 32.85379, 32.89882, 32.9437, 
    32.98843, 33.03302, 33.07745, 33.12174, 33.16588, 33.20988, 33.25372, 
    33.29741, 33.34095, 33.38434, 33.42758, 33.47067, 33.51361, 33.55639, 
    33.59903, 33.64151, 33.68383, 33.72601, 33.76802, 33.80989, 33.8516, 
    33.89316, 33.93456, 33.9758, 34.01689, 34.05782, 34.0986, 34.13922, 
    34.17968, 34.21998, 34.26013, 34.30012, 34.33994, 34.37961, 34.41912, 
    34.45847, 34.49766, 34.53669, 34.57556, 34.61426, 34.65281, 34.69119, 
    34.72941, 34.76747, 34.80536, 34.84309, 34.88066, 34.91806, 34.9553, 
    34.99237, 35.02929, 35.06603, 35.1026, 35.13902, 35.17526, 35.21134, 
    35.24725, 35.28299, 35.31857, 35.35398, 35.38921, 35.42428, 35.45918, 
    35.49392, 35.52848, 35.56287, 35.59709, 35.63114, 35.66501, 35.69872, 
    35.73225, 35.76562, 35.79881, 35.83183, 35.86467, 35.89734, 35.92983, 
    35.96215, 35.9943, 36.02628, 36.05807, 36.08969, 36.12114, 36.15241, 
    36.18351, 36.21442, 36.24516, 36.27573, 36.30611, 36.33632, 36.36635, 
    36.3962, 36.42587, 36.45536, 36.48467, 36.51381, 36.54276, 36.57153, 
    36.60012, 36.62853, 36.65676, 36.68481, 36.71267, 36.74036, 36.76786, 
    36.79517, 36.82231, 36.84926, 36.87603, 36.90261, 36.92901, 36.95523, 
    36.98126, 37.0071, 37.03276, 37.05824, 37.08352, 37.10863, 37.13354, 
    37.15827, 37.18281, 37.20717, 37.23133, 37.25531, 37.2791, 37.30271, 
    37.32612, 37.34935, 37.37238, 37.39523, 37.41788, 37.44035, 37.46263, 
    37.48472, 37.50661, 37.52832, 37.54984, 37.57116, 37.59229, 37.61323, 
    37.63398, 37.65453, 37.67489, 37.69506, 37.71504, 37.73483, 37.75441, 
    37.77381, 37.79301, 37.81202, 37.83084, 37.84946, 37.86788, 37.88611, 
    37.90414, 37.92199, 37.93963, 37.95708, 37.97433, 37.99139, 38.00824, 
    38.02491, 38.04137, 38.05764, 38.07372, 38.08959, 38.10527, 38.12075, 
    38.13603, 38.15111, 38.166, 38.18068, 38.19517, 38.20946, 38.22355, 
    38.23744, 38.25113, 38.26463, 38.27792, 38.29101, 38.30391, 38.3166, 
    38.32909, 38.34138, 38.35347, 38.36536, 38.37706, 38.38855, 38.39983, 
    38.41092, 38.42181, 38.43249, 38.44297, 38.45325, 38.46333, 38.47321, 
    38.48289, 38.49236, 38.50163, 38.5107, 38.51956, 38.52822, 38.53669, 
    38.54494, 38.553, 38.56085, 38.5685, 38.57594, 38.58318, 38.59022, 
    38.59705, 38.60369, 38.61011, 38.61634, 38.62236, 38.62817, 38.63378, 
    38.63919, 38.64439, 38.64939, 38.65419, 38.65878, 38.66317, 38.66735, 
    38.67133, 38.6751, 38.67867, 38.68203, 38.68519, 38.68814, 38.6909, 
    38.69344, 38.69578, 38.69791, 38.69984, 38.70157, 38.70309, 38.70441, 
    38.70552, 38.70642, 38.70713, 38.70762, 38.70791, 38.708, 38.70788, 
    38.70756, 38.70703, 38.7063, 38.70536, 38.70421, 38.70287, 38.70131, 
    38.69955, 38.69759, 38.69542, 38.69305, 38.69047, 38.68769, 38.6847, 
    38.68151, 38.67812, 38.67451, 38.67071, 38.6667, 38.66249, 38.65807, 
    38.65344, 38.64862, 38.64359, 38.63835, 38.63291, 38.62727, 38.62142, 
    38.61536, 38.60911, 38.60265, 38.59599, 38.58912, 38.58205, 38.57478, 
    38.5673, 38.55962, 38.55174, 38.54365, 38.53536, 38.52687, 38.51817, 
    38.50928, 38.50018, 38.49088, 38.48137, 38.47166, 38.46175, 38.45164, 
    38.44133, 38.43081, 38.4201, 38.40918, 38.39806, 38.38674, 38.37522, 
    38.3635, 38.35157, 38.33945, 38.32713, 38.3146, 38.30188, 38.28895, 
    38.27583, 38.2625, 38.24898, 38.23526, 38.22133, 38.20721, 38.19289, 
    38.17837, 38.16365, 38.14874, 38.13362, 38.11831, 38.1028, 38.08709, 
    38.07119, 38.05508, 38.03878, 38.02229, 38.00559, 37.9887, 37.97161, 
    37.95433, 37.93685, 37.91918, 37.90131, 37.88324, 37.86498, 37.84652, 
    37.82787, 37.80903, 37.78999, 37.77076, 37.75133, 37.73171, 37.71189, 
    37.69189, 37.67168, 37.65129, 37.63071, 37.60993, 37.58896, 37.5678, 
    37.54644, 37.5249, 37.50316, 37.48124, 37.45912, 37.43681, 37.41431, 
    37.39163, 37.36875, 37.34568, 37.32243, 37.29898, 37.27535, 37.25153, 
    37.22752, 37.20333, 37.17894, 37.15437, 37.12961, 37.10467, 37.07954, 
    37.05422, 37.02872, 37.00303, 36.97715, 36.95109, 36.92485, 36.89842, 
    36.87181, 36.84501, 36.81803, 36.79087, 36.76352, 36.73599, 36.70828, 
    36.68038, 36.65231, 36.62405, 36.59561, 36.56699, 36.53819, 36.50921, 
    36.48005, 36.45071, 36.42119, 36.39149, 36.36161, 36.33155, 36.30132, 
    36.2709, 36.24031, 36.20955, 36.1786, 36.14748, 36.11618, 36.08471, 
    36.05305, 36.02123, 35.98923, 35.95705, 35.92471, 35.89218, 35.85949, 
    35.82661, 35.79357,
  32.11715, 32.16483, 32.21238, 32.25978, 32.30704, 32.35416, 32.40113, 
    32.44797, 32.49466, 32.54121, 32.58761, 32.63387, 32.67999, 32.72596, 
    32.77179, 32.81747, 32.86301, 32.9084, 32.95364, 32.99874, 33.04369, 
    33.08849, 33.13315, 33.17765, 33.22201, 33.26622, 33.31028, 33.35419, 
    33.39795, 33.44156, 33.48502, 33.52833, 33.57148, 33.61449, 33.65734, 
    33.70004, 33.74259, 33.78498, 33.82722, 33.86931, 33.91124, 33.95302, 
    33.99464, 34.03611, 34.07742, 34.11858, 34.15957, 34.20042, 34.2411, 
    34.28163, 34.32199, 34.36221, 34.40226, 34.44215, 34.48188, 34.52146, 
    34.56087, 34.60012, 34.63922, 34.67815, 34.71692, 34.75553, 34.79397, 
    34.83226, 34.87038, 34.90833, 34.94613, 34.98376, 35.02122, 35.05853, 
    35.09566, 35.13263, 35.16944, 35.20607, 35.24255, 35.27885, 35.31499, 
    35.35096, 35.38677, 35.4224, 35.45787, 35.49317, 35.5283, 35.56326, 
    35.59805, 35.63267, 35.66712, 35.7014, 35.7355, 35.76944, 35.8032, 
    35.8368, 35.87022, 35.90346, 35.93653, 35.96944, 36.00216, 36.03472, 
    36.0671, 36.0993, 36.13133, 36.16318, 36.19486, 36.22636, 36.25768, 
    36.28883, 36.31981, 36.3506, 36.38121, 36.41165, 36.44191, 36.472, 
    36.5019, 36.53162, 36.56116, 36.59053, 36.61972, 36.64872, 36.67754, 
    36.70618, 36.73465, 36.76292, 36.79102, 36.81894, 36.84667, 36.87422, 
    36.90159, 36.92877, 36.95577, 36.98259, 37.00922, 37.03567, 37.06193, 
    37.08801, 37.1139, 37.13961, 37.16513, 37.19046, 37.21561, 37.24057, 
    37.26534, 37.28993, 37.31433, 37.33854, 37.36256, 37.3864, 37.41005, 
    37.4335, 37.45677, 37.47985, 37.50274, 37.52544, 37.54795, 37.57026, 
    37.59239, 37.61433, 37.63607, 37.65763, 37.67899, 37.70016, 37.72114, 
    37.74193, 37.76252, 37.78292, 37.80313, 37.82314, 37.84296, 37.86259, 
    37.88202, 37.90126, 37.92031, 37.93916, 37.95781, 37.97627, 37.99453, 
    38.0126, 38.03048, 38.04815, 38.06564, 38.08292, 38.10001, 38.1169, 
    38.13359, 38.15009, 38.16639, 38.1825, 38.1984, 38.2141, 38.22961, 
    38.24492, 38.26004, 38.27495, 38.28967, 38.30418, 38.3185, 38.33261, 
    38.34653, 38.36025, 38.37377, 38.38708, 38.4002, 38.41312, 38.42584, 
    38.43835, 38.45067, 38.46279, 38.4747, 38.48642, 38.49792, 38.50924, 
    38.52034, 38.53125, 38.54196, 38.55246, 38.56276, 38.57286, 38.58276, 
    38.59245, 38.60194, 38.61123, 38.62032, 38.6292, 38.63788, 38.64635, 
    38.65462, 38.6627, 38.67056, 38.67823, 38.68568, 38.69294, 38.69999, 
    38.70684, 38.71348, 38.71992, 38.72616, 38.73219, 38.73801, 38.74364, 
    38.74906, 38.75427, 38.75928, 38.76408, 38.76868, 38.77308, 38.77727, 
    38.78125, 38.78503, 38.78861, 38.79198, 38.79514, 38.7981, 38.80086, 
    38.80341, 38.80576, 38.8079, 38.80983, 38.81156, 38.81308, 38.8144, 
    38.81551, 38.81642, 38.81712, 38.81762, 38.81791, 38.818, 38.81788, 
    38.81755, 38.81703, 38.81629, 38.81535, 38.81421, 38.81285, 38.8113, 
    38.80954, 38.80757, 38.8054, 38.80302, 38.80044, 38.79765, 38.79466, 
    38.79146, 38.78806, 38.78445, 38.78064, 38.77662, 38.7724, 38.76797, 
    38.76334, 38.7585, 38.75346, 38.74821, 38.74276, 38.73711, 38.73125, 
    38.72519, 38.71892, 38.71244, 38.70577, 38.69889, 38.69181, 38.68452, 
    38.67702, 38.66933, 38.66143, 38.65333, 38.64503, 38.63652, 38.6278, 
    38.61889, 38.60977, 38.60045, 38.59093, 38.5812, 38.57127, 38.56115, 
    38.55081, 38.54028, 38.52954, 38.5186, 38.50746, 38.49612, 38.48457, 
    38.47283, 38.46088, 38.44874, 38.43639, 38.42384, 38.41109, 38.39814, 
    38.38499, 38.37164, 38.35809, 38.34435, 38.33039, 38.31625, 38.3019, 
    38.28735, 38.27261, 38.25766, 38.24252, 38.22717, 38.21164, 38.1959, 
    38.17996, 38.16383, 38.1475, 38.13097, 38.11424, 38.09732, 38.0802, 
    38.06288, 38.04537, 38.02766, 38.00976, 37.99166, 37.97336, 37.95487, 
    37.93619, 37.91731, 37.89823, 37.87896, 37.8595, 37.83984, 37.81999, 
    37.79995, 37.77971, 37.75928, 37.73865, 37.71783, 37.69683, 37.67562, 
    37.65423, 37.63265, 37.61087, 37.58891, 37.56675, 37.5444, 37.52186, 
    37.49913, 37.47621, 37.4531, 37.42981, 37.40631, 37.38264, 37.35878, 
    37.33472, 37.31048, 37.28605, 37.26144, 37.23663, 37.21164, 37.18647, 
    37.1611, 37.13555, 37.10982, 37.0839, 37.05779, 37.0315, 37.00502, 
    36.97836, 36.95152, 36.92448, 36.89727, 36.86988, 36.8423, 36.81453, 
    36.78659, 36.75846, 36.73016, 36.70167, 36.673, 36.64414, 36.61511, 
    36.5859, 36.5565, 36.52693, 36.49718, 36.46725, 36.43714, 36.40685, 
    36.37638, 36.34574, 36.31491, 36.28392, 36.25274, 36.22139, 36.18986, 
    36.15815, 36.12627, 36.09422, 36.06199, 36.02958, 35.997, 35.96424, 
    35.93132, 35.89822,
  32.21572, 32.26347, 32.31108, 32.35855, 32.40589, 32.45308, 32.50012, 
    32.54703, 32.59379, 32.64041, 32.68688, 32.73322, 32.7794, 32.82544, 
    32.87134, 32.91709, 32.9627, 33.00816, 33.05347, 33.09864, 33.14366, 
    33.18853, 33.23325, 33.27783, 33.32226, 33.36654, 33.41066, 33.45464, 
    33.49847, 33.54215, 33.58567, 33.62905, 33.67228, 33.71535, 33.75827, 
    33.80104, 33.84365, 33.88611, 33.92842, 33.97057, 34.01257, 34.05442, 
    34.09611, 34.13764, 34.17902, 34.22024, 34.2613, 34.30221, 34.34296, 
    34.38355, 34.42398, 34.46426, 34.50438, 34.54434, 34.58414, 34.62378, 
    34.66325, 34.70257, 34.74173, 34.78072, 34.81956, 34.85823, 34.89674, 
    34.93509, 34.97327, 35.01129, 35.04914, 35.08684, 35.12437, 35.16173, 
    35.19893, 35.23596, 35.27283, 35.30952, 35.34606, 35.38243, 35.41862, 
    35.45466, 35.49052, 35.52622, 35.56174, 35.5971, 35.63229, 35.66731, 
    35.70216, 35.73684, 35.77135, 35.80569, 35.83986, 35.87385, 35.90767, 
    35.94132, 35.9748, 36.0081, 36.04123, 36.07419, 36.10698, 36.13958, 
    36.17202, 36.20428, 36.23636, 36.26827, 36.30001, 36.33156, 36.36294, 
    36.39415, 36.42517, 36.45602, 36.48669, 36.51718, 36.5475, 36.57763, 
    36.60759, 36.63736, 36.66696, 36.69638, 36.72561, 36.75467, 36.78354, 
    36.81224, 36.84075, 36.86908, 36.89723, 36.92519, 36.95298, 36.98058, 
    37.00799, 37.03522, 37.06227, 37.08914, 37.11582, 37.14231, 37.16862, 
    37.19475, 37.22069, 37.24644, 37.27201, 37.29739, 37.32258, 37.34759, 
    37.37241, 37.39704, 37.42148, 37.44574, 37.46981, 37.49369, 37.51738, 
    37.54087, 37.56419, 37.58731, 37.61024, 37.63298, 37.65553, 37.67789, 
    37.70006, 37.72203, 37.74382, 37.76542, 37.78682, 37.80803, 37.82905, 
    37.84987, 37.8705, 37.89094, 37.91119, 37.93124, 37.9511, 37.97076, 
    37.99023, 38.00951, 38.02859, 38.04747, 38.06616, 38.08466, 38.10295, 
    38.12106, 38.13897, 38.15667, 38.17419, 38.19151, 38.20863, 38.22555, 
    38.24228, 38.2588, 38.27514, 38.29127, 38.30721, 38.32294, 38.33848, 
    38.35382, 38.36896, 38.3839, 38.39864, 38.41319, 38.42753, 38.44168, 
    38.45562, 38.46936, 38.48291, 38.49625, 38.5094, 38.52234, 38.53508, 
    38.54762, 38.55996, 38.5721, 38.58404, 38.59577, 38.6073, 38.61864, 
    38.62977, 38.64069, 38.65142, 38.66195, 38.67226, 38.68238, 38.6923, 
    38.70201, 38.71152, 38.72083, 38.72993, 38.73883, 38.74752, 38.75602, 
    38.76431, 38.77239, 38.78027, 38.78795, 38.79543, 38.8027, 38.80976, 
    38.81662, 38.82328, 38.82973, 38.83598, 38.84202, 38.84786, 38.85349, 
    38.85892, 38.86415, 38.86916, 38.87398, 38.87859, 38.88299, 38.88719, 
    38.89118, 38.89497, 38.89855, 38.90193, 38.9051, 38.90807, 38.91083, 
    38.91338, 38.91573, 38.91787, 38.91981, 38.92155, 38.92307, 38.92439, 
    38.92551, 38.92642, 38.92712, 38.92762, 38.92791, 38.928, 38.92788, 
    38.92756, 38.92702, 38.92629, 38.92535, 38.9242, 38.92284, 38.92128, 
    38.91952, 38.91755, 38.91537, 38.91299, 38.9104, 38.90761, 38.90461, 
    38.90141, 38.898, 38.89438, 38.89056, 38.88654, 38.88231, 38.87787, 
    38.87323, 38.86839, 38.86333, 38.85808, 38.85262, 38.84695, 38.84108, 
    38.835, 38.82872, 38.82224, 38.81555, 38.80866, 38.80156, 38.79426, 
    38.78675, 38.77904, 38.77113, 38.76301, 38.75469, 38.74616, 38.73743, 
    38.7285, 38.71937, 38.71003, 38.70049, 38.69074, 38.6808, 38.67065, 
    38.66029, 38.64974, 38.63898, 38.62802, 38.61686, 38.6055, 38.59393, 
    38.58216, 38.57019, 38.55802, 38.54565, 38.53308, 38.52031, 38.50733, 
    38.49416, 38.48078, 38.46721, 38.45343, 38.43945, 38.42527, 38.4109, 
    38.39632, 38.38155, 38.36658, 38.35141, 38.33603, 38.32047, 38.3047, 
    38.28873, 38.27256, 38.2562, 38.23964, 38.22289, 38.20593, 38.18878, 
    38.17143, 38.15388, 38.13614, 38.11821, 38.10007, 38.08174, 38.06322, 
    38.0445, 38.02558, 38.00647, 37.98716, 37.96766, 37.94797, 37.92808, 
    37.908, 37.88772, 37.86725, 37.84659, 37.82573, 37.80469, 37.78345, 
    37.76201, 37.74039, 37.71857, 37.69656, 37.67437, 37.65198, 37.62939, 
    37.60662, 37.58366, 37.56051, 37.53717, 37.51364, 37.48992, 37.46601, 
    37.44191, 37.41763, 37.39315, 37.3685, 37.34365, 37.31861, 37.29338, 
    37.26797, 37.24238, 37.2166, 37.19063, 37.16447, 37.13813, 37.11161, 
    37.0849, 37.05801, 37.03093, 37.00367, 36.97622, 36.94859, 36.92078, 
    36.89279, 36.86461, 36.83625, 36.80771, 36.77899, 36.75008, 36.721, 
    36.69174, 36.66229, 36.63267, 36.60286, 36.57288, 36.54271, 36.51237, 
    36.48185, 36.45115, 36.42028, 36.38922, 36.35799, 36.32658, 36.295, 
    36.26324, 36.2313, 36.19919, 36.1669, 36.13444, 36.1018, 36.06899, 
    36.03601, 36.00285,
  32.31425, 32.36208, 32.40976, 32.45731, 32.50471, 32.55197, 32.59909, 
    32.64606, 32.69289, 32.73959, 32.78613, 32.83253, 32.87879, 32.9249, 
    32.97087, 33.01669, 33.06237, 33.10789, 33.15328, 33.19851, 33.2436, 
    33.28854, 33.33334, 33.37798, 33.42248, 33.46682, 33.51102, 33.55507, 
    33.59896, 33.64271, 33.68631, 33.72975, 33.77304, 33.81618, 33.85917, 
    33.90201, 33.94469, 33.98722, 34.02959, 34.07182, 34.11388, 34.15579, 
    34.19755, 34.23915, 34.28059, 34.32188, 34.36301, 34.40398, 34.4448, 
    34.48546, 34.52596, 34.5663, 34.60648, 34.6465, 34.68637, 34.72607, 
    34.76561, 34.805, 34.84422, 34.88328, 34.92217, 34.96091, 34.99948, 
    35.03789, 35.07614, 35.11422, 35.15214, 35.1899, 35.22749, 35.26492, 
    35.30217, 35.33927, 35.3762, 35.41296, 35.44955, 35.48598, 35.52224, 
    35.55834, 35.59426, 35.63002, 35.66561, 35.70103, 35.73627, 35.77135, 
    35.80626, 35.841, 35.87557, 35.90997, 35.94419, 35.97824, 36.01212, 
    36.04583, 36.07937, 36.11273, 36.14592, 36.17893, 36.21177, 36.24444, 
    36.27693, 36.30925, 36.34139, 36.37335, 36.40514, 36.43675, 36.46819, 
    36.49945, 36.53053, 36.56143, 36.59215, 36.6227, 36.65307, 36.68325, 
    36.71326, 36.7431, 36.77274, 36.80221, 36.8315, 36.86061, 36.88953, 
    36.91828, 36.94684, 36.97522, 37.00342, 37.03144, 37.05927, 37.08692, 
    37.11439, 37.14167, 37.16877, 37.19568, 37.22241, 37.24895, 37.27531, 
    37.30148, 37.32747, 37.35327, 37.37888, 37.40431, 37.42955, 37.4546, 
    37.47946, 37.50414, 37.52863, 37.55293, 37.57704, 37.60096, 37.62469, 
    37.64824, 37.67159, 37.69476, 37.71773, 37.74052, 37.76311, 37.78551, 
    37.80772, 37.82974, 37.85156, 37.8732, 37.89464, 37.91589, 37.93695, 
    37.95781, 37.97848, 37.99896, 38.01924, 38.03933, 38.05923, 38.07893, 
    38.09843, 38.11774, 38.13686, 38.15578, 38.17451, 38.19304, 38.21137, 
    38.22951, 38.24745, 38.26519, 38.28274, 38.30009, 38.31724, 38.3342, 
    38.35096, 38.36752, 38.38388, 38.40004, 38.416, 38.43177, 38.44734, 
    38.46271, 38.47788, 38.49285, 38.50762, 38.52219, 38.53656, 38.55074, 
    38.5647, 38.57848, 38.59204, 38.60542, 38.61858, 38.63155, 38.64432, 
    38.65688, 38.66925, 38.68141, 38.69337, 38.70513, 38.71668, 38.72803, 
    38.73919, 38.75014, 38.76088, 38.77143, 38.78177, 38.7919, 38.80184, 
    38.81157, 38.8211, 38.83042, 38.83954, 38.84846, 38.85717, 38.86568, 
    38.87399, 38.88209, 38.88999, 38.89768, 38.90517, 38.91245, 38.91953, 
    38.92641, 38.93307, 38.93954, 38.9458, 38.95185, 38.9577, 38.96335, 
    38.96879, 38.97402, 38.97905, 38.98387, 38.98849, 38.9929, 38.99711, 
    39.00111, 39.00491, 39.0085, 39.01188, 39.01506, 39.01803, 39.02079, 
    39.02335, 39.02571, 39.02785, 39.0298, 39.03153, 39.03306, 39.03439, 
    39.0355, 39.03642, 39.03712, 39.03762, 39.03791, 39.038, 39.03788, 
    39.03756, 39.03702, 39.03629, 39.03534, 39.03419, 39.03283, 39.03127, 
    39.0295, 39.02753, 39.02535, 39.02296, 39.02037, 39.01757, 39.01457, 
    39.01136, 39.00794, 39.00432, 39.00049, 38.99646, 38.99222, 38.98777, 
    38.98312, 38.97827, 38.97321, 38.96794, 38.96247, 38.95679, 38.95091, 
    38.94482, 38.93853, 38.93203, 38.92533, 38.91843, 38.91131, 38.904, 
    38.89648, 38.88875, 38.88082, 38.87269, 38.86435, 38.85581, 38.84706, 
    38.83812, 38.82896, 38.81961, 38.81004, 38.80028, 38.79031, 38.78014, 
    38.76977, 38.7592, 38.74842, 38.73744, 38.72625, 38.71487, 38.70328, 
    38.69149, 38.6795, 38.6673, 38.65491, 38.64231, 38.62951, 38.61652, 
    38.60331, 38.58991, 38.57631, 38.56251, 38.54851, 38.5343, 38.5199, 
    38.5053, 38.49049, 38.47549, 38.46029, 38.44489, 38.42929, 38.41349, 
    38.3975, 38.3813, 38.36491, 38.34832, 38.33153, 38.31454, 38.29736, 
    38.27998, 38.2624, 38.24462, 38.22665, 38.20848, 38.19012, 38.17156, 
    38.1528, 38.13385, 38.1147, 38.09536, 38.07582, 38.05609, 38.03617, 
    38.01604, 37.99573, 37.97522, 37.95452, 37.93363, 37.91254, 37.89126, 
    37.86979, 37.84813, 37.82627, 37.80422, 37.78198, 37.75955, 37.73692, 
    37.71411, 37.69111, 37.66791, 37.64453, 37.62096, 37.59719, 37.57324, 
    37.5491, 37.52477, 37.50025, 37.47554, 37.45065, 37.42557, 37.4003, 
    37.37484, 37.3492, 37.32337, 37.29735, 37.27115, 37.24476, 37.21819, 
    37.19143, 37.16449, 37.13736, 37.11005, 37.08256, 37.05488, 37.02702, 
    36.99897, 36.97075, 36.94234, 36.91375, 36.88497, 36.85602, 36.82688, 
    36.79756, 36.76807, 36.73839, 36.70853, 36.67849, 36.64827, 36.61788, 
    36.58731, 36.55655, 36.52562, 36.49451, 36.46323, 36.43176, 36.40012, 
    36.36831, 36.33632, 36.30415, 36.2718, 36.23928, 36.20659, 36.17372, 
    36.14068, 36.10746,
  32.41277, 32.46066, 32.50842, 32.55603, 32.60351, 32.65084, 32.69802, 
    32.74507, 32.79198, 32.83873, 32.88535, 32.93182, 32.97815, 33.02433, 
    33.07037, 33.11626, 33.16201, 33.20761, 33.25306, 33.29837, 33.34352, 
    33.38853, 33.4334, 33.47811, 33.52267, 33.56709, 33.61136, 33.65547, 
    33.69944, 33.74326, 33.78692, 33.83043, 33.87379, 33.917, 33.96006, 
    34.00296, 34.04571, 34.08831, 34.13075, 34.17303, 34.21517, 34.25714, 
    34.29897, 34.34063, 34.38214, 34.4235, 34.46469, 34.50574, 34.54662, 
    34.58734, 34.62791, 34.66832, 34.70856, 34.74865, 34.78858, 34.82835, 
    34.86795, 34.9074, 34.94669, 34.98581, 35.02477, 35.06357, 35.10221, 
    35.14068, 35.17899, 35.21714, 35.25512, 35.29294, 35.33059, 35.36808, 
    35.40541, 35.44256, 35.47955, 35.51638, 35.55304, 35.58952, 35.62585, 
    35.662, 35.69799, 35.7338, 35.76945, 35.80493, 35.84024, 35.87538, 
    35.91035, 35.94514, 35.97977, 36.01423, 36.04851, 36.08262, 36.11656, 
    36.15033, 36.18392, 36.21734, 36.25059, 36.28366, 36.31656, 36.34928, 
    36.38183, 36.4142, 36.4464, 36.47842, 36.51026, 36.54193, 36.57342, 
    36.60473, 36.63587, 36.66682, 36.69761, 36.7282, 36.75863, 36.78887, 
    36.81893, 36.84881, 36.87851, 36.90804, 36.93738, 36.96654, 36.99551, 
    37.02431, 37.05293, 37.08136, 37.1096, 37.13767, 37.16555, 37.19325, 
    37.22077, 37.2481, 37.27525, 37.30221, 37.32899, 37.35558, 37.38198, 
    37.4082, 37.43423, 37.46008, 37.48574, 37.51122, 37.5365, 37.5616, 
    37.58651, 37.61123, 37.63577, 37.66011, 37.68427, 37.70823, 37.73201, 
    37.7556, 37.779, 37.8022, 37.82522, 37.84805, 37.87068, 37.89312, 
    37.91537, 37.93743, 37.9593, 37.98097, 38.00246, 38.02375, 38.04484, 
    38.06574, 38.08645, 38.10697, 38.12729, 38.14742, 38.16735, 38.18709, 
    38.20663, 38.22598, 38.24513, 38.26408, 38.28284, 38.30141, 38.31978, 
    38.33795, 38.35592, 38.3737, 38.39128, 38.40866, 38.42585, 38.44284, 
    38.45963, 38.47622, 38.49261, 38.50881, 38.5248, 38.5406, 38.5562, 
    38.5716, 38.5868, 38.6018, 38.61659, 38.63119, 38.64559, 38.65979, 
    38.67379, 38.68758, 38.70118, 38.71458, 38.72777, 38.74076, 38.75356, 
    38.76614, 38.77853, 38.79071, 38.8027, 38.81448, 38.82606, 38.83743, 
    38.84861, 38.85958, 38.87034, 38.88091, 38.89127, 38.90142, 38.91138, 
    38.92113, 38.93068, 38.94002, 38.94916, 38.95809, 38.96682, 38.97535, 
    38.98367, 38.99179, 38.9997, 39.0074, 39.01491, 39.02221, 39.0293, 
    39.03619, 39.04287, 39.04935, 39.05562, 39.06169, 39.06755, 39.0732, 
    39.07865, 39.0839, 39.08894, 39.09377, 39.09839, 39.10281, 39.10703, 
    39.11104, 39.11484, 39.11843, 39.12183, 39.12501, 39.12799, 39.13076, 
    39.13332, 39.13568, 39.13784, 39.13978, 39.14152, 39.14305, 39.14438, 
    39.1455, 39.14641, 39.14712, 39.14762, 39.14791, 39.148, 39.14788, 
    39.14755, 39.14702, 39.14628, 39.14534, 39.14418, 39.14283, 39.14126, 
    39.13949, 39.13751, 39.13532, 39.13293, 39.13034, 39.12753, 39.12452, 
    39.1213, 39.11788, 39.11425, 39.11042, 39.10638, 39.10213, 39.09768, 
    39.09302, 39.08815, 39.08308, 39.0778, 39.07232, 39.06664, 39.06074, 
    39.05464, 39.04834, 39.04183, 39.03511, 39.02819, 39.02106, 39.01374, 
    39.0062, 38.99846, 38.99052, 38.98236, 38.97401, 38.96545, 38.95669, 
    38.94772, 38.93855, 38.92918, 38.9196, 38.90982, 38.89983, 38.88964, 
    38.87925, 38.86865, 38.85785, 38.84685, 38.83565, 38.82424, 38.81263, 
    38.80082, 38.7888, 38.77658, 38.76416, 38.75154, 38.73872, 38.7257, 
    38.71247, 38.69904, 38.68542, 38.67159, 38.65756, 38.64333, 38.62889, 
    38.61427, 38.59943, 38.5844, 38.56918, 38.55375, 38.53812, 38.52229, 
    38.50626, 38.49003, 38.47361, 38.45699, 38.44017, 38.42315, 38.40593, 
    38.38852, 38.3709, 38.3531, 38.33509, 38.31689, 38.29849, 38.27989, 
    38.2611, 38.24211, 38.22293, 38.20355, 38.18398, 38.16421, 38.14425, 
    38.12409, 38.10374, 38.08319, 38.06245, 38.04152, 38.02039, 37.99907, 
    37.97756, 37.95585, 37.93396, 37.91187, 37.88958, 37.86711, 37.84444, 
    37.82159, 37.79854, 37.77531, 37.75188, 37.72826, 37.70446, 37.68046, 
    37.65627, 37.6319, 37.60733, 37.58258, 37.55764, 37.53252, 37.5072, 
    37.4817, 37.45601, 37.43013, 37.40407, 37.37782, 37.35138, 37.32476, 
    37.29795, 37.27097, 37.24379, 37.21643, 37.18888, 37.16116, 37.13324, 
    37.10515, 37.07687, 37.04841, 37.01977, 36.99094, 36.96194, 36.93275, 
    36.90338, 36.87383, 36.8441, 36.81419, 36.7841, 36.75383, 36.72338, 
    36.69275, 36.66194, 36.63095, 36.59979, 36.56845, 36.53693, 36.50524, 
    36.47337, 36.44131, 36.40909, 36.37669, 36.34412, 36.31137, 36.27844, 
    36.24534, 36.21207,
  32.51125, 32.55922, 32.60705, 32.65474, 32.70228, 32.74968, 32.79694, 
    32.84406, 32.89103, 32.93786, 32.98455, 33.03109, 33.07749, 33.12374, 
    33.16985, 33.21581, 33.26162, 33.30729, 33.35282, 33.39819, 33.44342, 
    33.4885, 33.53343, 33.57822, 33.62285, 33.66734, 33.71167, 33.75586, 
    33.79989, 33.84377, 33.8875, 33.93109, 33.97451, 34.01779, 34.06092, 
    34.10389, 34.14671, 34.18937, 34.23188, 34.27423, 34.31643, 34.35848, 
    34.40037, 34.4421, 34.48368, 34.5251, 34.56636, 34.60747, 34.64841, 
    34.68921, 34.72984, 34.77031, 34.81062, 34.85078, 34.89077, 34.9306, 
    34.97028, 35.00979, 35.04914, 35.08833, 35.12735, 35.16622, 35.20492, 
    35.24345, 35.28183, 35.32004, 35.35809, 35.39597, 35.43368, 35.47123, 
    35.50862, 35.54584, 35.58289, 35.61978, 35.65649, 35.69305, 35.72943, 
    35.76564, 35.80169, 35.83757, 35.87328, 35.90882, 35.94419, 35.97939, 
    36.01442, 36.04927, 36.08396, 36.11847, 36.15282, 36.18699, 36.22099, 
    36.25481, 36.28846, 36.32194, 36.35524, 36.38837, 36.42133, 36.45411, 
    36.48671, 36.51914, 36.55139, 36.58347, 36.61537, 36.64709, 36.67864, 
    36.71001, 36.7412, 36.77221, 36.80304, 36.83369, 36.86417, 36.89447, 
    36.92458, 36.95452, 36.98427, 37.01385, 37.04324, 37.07245, 37.10148, 
    37.13033, 37.159, 37.18748, 37.21578, 37.24389, 37.27183, 37.29958, 
    37.32714, 37.35452, 37.38172, 37.40873, 37.43555, 37.46219, 37.48865, 
    37.51492, 37.541, 37.56689, 37.5926, 37.61812, 37.64345, 37.66859, 
    37.69355, 37.71832, 37.7429, 37.76728, 37.79148, 37.81549, 37.83932, 
    37.86295, 37.88639, 37.90964, 37.9327, 37.95557, 37.97824, 38.00072, 
    38.02302, 38.04512, 38.06703, 38.08874, 38.11026, 38.13159, 38.15273, 
    38.17367, 38.19442, 38.21497, 38.23533, 38.2555, 38.27547, 38.29524, 
    38.31482, 38.33421, 38.35339, 38.37239, 38.39118, 38.40978, 38.42818, 
    38.44639, 38.4644, 38.48221, 38.49982, 38.51724, 38.53446, 38.55148, 
    38.5683, 38.58492, 38.60135, 38.61757, 38.6336, 38.64943, 38.66505, 
    38.68048, 38.69571, 38.71074, 38.72556, 38.74019, 38.75462, 38.76884, 
    38.78287, 38.79669, 38.81031, 38.82373, 38.83695, 38.84997, 38.86279, 
    38.8754, 38.88781, 38.90002, 38.91203, 38.92383, 38.93543, 38.94683, 
    38.95802, 38.96901, 38.9798, 38.99039, 39.00077, 39.01094, 39.02092, 
    39.03069, 39.04025, 39.04961, 39.05877, 39.06772, 39.07647, 39.08501, 
    39.09335, 39.10148, 39.10941, 39.11713, 39.12465, 39.13196, 39.13907, 
    39.14597, 39.15266, 39.15915, 39.16544, 39.17152, 39.17739, 39.18306, 
    39.18851, 39.19377, 39.19882, 39.20366, 39.2083, 39.21273, 39.21695, 
    39.22097, 39.22477, 39.22838, 39.23178, 39.23497, 39.23795, 39.24073, 
    39.2433, 39.24566, 39.24781, 39.24976, 39.25151, 39.25304, 39.25437, 
    39.25549, 39.25641, 39.25712, 39.25762, 39.25791, 39.258, 39.25788, 
    39.25755, 39.25702, 39.25628, 39.25533, 39.25418, 39.25282, 39.25125, 
    39.24947, 39.24749, 39.2453, 39.2429, 39.2403, 39.23749, 39.23447, 
    39.23125, 39.22782, 39.22419, 39.22034, 39.21629, 39.21204, 39.20758, 
    39.20291, 39.19803, 39.19296, 39.18767, 39.18217, 39.17648, 39.17057, 
    39.16446, 39.15814, 39.15162, 39.14489, 39.13796, 39.13082, 39.12347, 
    39.11592, 39.10817, 39.10021, 39.09204, 39.08367, 39.0751, 39.06632, 
    39.05733, 39.04815, 39.03875, 39.02916, 39.01936, 39.00935, 38.99914, 
    38.98873, 38.97811, 38.96729, 38.95626, 38.94504, 38.93361, 38.92198, 
    38.91014, 38.8981, 38.88586, 38.87342, 38.86077, 38.84793, 38.83488, 
    38.82162, 38.80817, 38.79452, 38.78066, 38.76661, 38.75235, 38.73789, 
    38.72323, 38.70837, 38.69331, 38.67805, 38.66259, 38.64693, 38.63108, 
    38.61502, 38.59876, 38.58231, 38.56565, 38.5488, 38.53175, 38.5145, 
    38.49705, 38.4794, 38.46156, 38.44352, 38.42529, 38.40685, 38.38822, 
    38.36939, 38.35037, 38.33115, 38.31174, 38.29213, 38.27232, 38.25232, 
    38.23212, 38.21173, 38.19115, 38.17037, 38.1494, 38.12823, 38.10687, 
    38.08532, 38.06358, 38.04163, 38.0195, 37.99718, 37.97467, 37.95196, 
    37.92906, 37.90597, 37.88269, 37.85922, 37.83556, 37.81171, 37.78767, 
    37.76344, 37.73902, 37.71441, 37.68961, 37.66463, 37.63945, 37.61409, 
    37.58854, 37.56281, 37.53688, 37.51077, 37.48447, 37.45799, 37.43132, 
    37.40447, 37.37743, 37.3502, 37.32279, 37.2952, 37.26742, 37.23946, 
    37.21132, 37.18298, 37.15447, 37.12578, 37.0969, 37.06784, 37.0386, 
    37.00918, 36.97958, 36.94979, 36.91983, 36.88969, 36.85936, 36.82886, 
    36.79818, 36.76731, 36.73627, 36.70506, 36.67366, 36.64209, 36.61034, 
    36.57841, 36.5463, 36.51402, 36.48157, 36.44893, 36.41613, 36.38314, 
    36.34999, 36.31665,
  32.60971, 32.65775, 32.70565, 32.75341, 32.80102, 32.8485, 32.89583, 
    32.94302, 32.99006, 33.03696, 33.08372, 33.13033, 33.1768, 33.22312, 
    33.2693, 33.31533, 33.36122, 33.40696, 33.45255, 33.49799, 33.54329, 
    33.58844, 33.63344, 33.6783, 33.723, 33.76755, 33.81196, 33.85621, 
    33.90031, 33.94427, 33.98807, 34.03172, 34.07521, 34.11856, 34.16175, 
    34.20479, 34.24768, 34.29041, 34.33298, 34.37541, 34.41768, 34.45979, 
    34.50174, 34.54354, 34.58519, 34.62667, 34.66801, 34.70918, 34.75019, 
    34.79105, 34.83175, 34.87228, 34.91266, 34.95288, 34.99294, 35.03284, 
    35.07258, 35.11216, 35.15157, 35.19082, 35.22991, 35.26884, 35.30761, 
    35.34621, 35.38464, 35.42292, 35.46103, 35.49897, 35.53675, 35.57436, 
    35.61181, 35.64909, 35.68621, 35.72316, 35.75994, 35.79655, 35.833, 
    35.86927, 35.90538, 35.94132, 35.97709, 36.01269, 36.04812, 36.08338, 
    36.11847, 36.15339, 36.18813, 36.22271, 36.25711, 36.29134, 36.32539, 
    36.35928, 36.39299, 36.42652, 36.45988, 36.49307, 36.52608, 36.55892, 
    36.59158, 36.62407, 36.65638, 36.68851, 36.72046, 36.75224, 36.78384, 
    36.81527, 36.84651, 36.87758, 36.90847, 36.93917, 36.9697, 37.00005, 
    37.03022, 37.06021, 37.09002, 37.11965, 37.14909, 37.17836, 37.20744, 
    37.23634, 37.26505, 37.29359, 37.32194, 37.35011, 37.37809, 37.40589, 
    37.4335, 37.46093, 37.48818, 37.51524, 37.54211, 37.5688, 37.5953, 
    37.62162, 37.64775, 37.67369, 37.69944, 37.72501, 37.75039, 37.77558, 
    37.80058, 37.82539, 37.85002, 37.87445, 37.8987, 37.92275, 37.94662, 
    37.97029, 37.99377, 38.01707, 38.04017, 38.06308, 38.0858, 38.10832, 
    38.13066, 38.1528, 38.17475, 38.1965, 38.21807, 38.23943, 38.26061, 
    38.28159, 38.30238, 38.32297, 38.34337, 38.36357, 38.38358, 38.40339, 
    38.42301, 38.44243, 38.46165, 38.48068, 38.49951, 38.51815, 38.53658, 
    38.55482, 38.57286, 38.59071, 38.60836, 38.62581, 38.64306, 38.66011, 
    38.67696, 38.69362, 38.71008, 38.72633, 38.74239, 38.75825, 38.7739, 
    38.78936, 38.80462, 38.81968, 38.83453, 38.84919, 38.86364, 38.87789, 
    38.89194, 38.9058, 38.91945, 38.93289, 38.94614, 38.95918, 38.97202, 
    38.98466, 38.99709, 39.00932, 39.02135, 39.03318, 39.0448, 39.05622, 
    39.06744, 39.07845, 39.08926, 39.09986, 39.11027, 39.12046, 39.13046, 
    39.14024, 39.14983, 39.15921, 39.16838, 39.17735, 39.18611, 39.19467, 
    39.20303, 39.21117, 39.21912, 39.22686, 39.23439, 39.24171, 39.24884, 
    39.25575, 39.26246, 39.26896, 39.27526, 39.28135, 39.28723, 39.29291, 
    39.29838, 39.30365, 39.3087, 39.31355, 39.3182, 39.32264, 39.32687, 
    39.33089, 39.33471, 39.33832, 39.34172, 39.34492, 39.34791, 39.35069, 
    39.35327, 39.35564, 39.3578, 39.35975, 39.3615, 39.36303, 39.36436, 
    39.36549, 39.36641, 39.36712, 39.36762, 39.36791, 39.368, 39.36788, 
    39.36755, 39.36702, 39.36628, 39.36533, 39.36417, 39.3628, 39.36123, 
    39.35946, 39.35747, 39.35527, 39.35287, 39.35027, 39.34745, 39.34443, 
    39.3412, 39.33776, 39.33412, 39.33027, 39.32621, 39.32195, 39.31748, 
    39.3128, 39.30791, 39.30283, 39.29753, 39.29203, 39.28632, 39.2804, 
    39.27428, 39.26794, 39.26141, 39.25467, 39.24772, 39.24057, 39.23321, 
    39.22565, 39.21788, 39.2099, 39.20172, 39.19333, 39.18474, 39.17595, 
    39.16694, 39.15773, 39.14832, 39.13871, 39.12889, 39.11886, 39.10863, 
    39.0982, 39.08756, 39.07672, 39.06568, 39.05443, 39.04298, 39.03132, 
    39.01946, 39.0074, 38.99514, 38.98267, 38.97, 38.95713, 38.94405, 
    38.93077, 38.9173, 38.90362, 38.88974, 38.87565, 38.86137, 38.84688, 
    38.8322, 38.81731, 38.80222, 38.78693, 38.77144, 38.75575, 38.73986, 
    38.72377, 38.70749, 38.691, 38.67431, 38.65743, 38.64034, 38.62306, 
    38.60558, 38.5879, 38.57003, 38.55195, 38.53368, 38.51521, 38.49654, 
    38.47768, 38.45862, 38.43937, 38.41992, 38.40027, 38.38043, 38.36039, 
    38.34016, 38.31973, 38.2991, 38.27829, 38.25727, 38.23607, 38.21467, 
    38.19307, 38.17129, 38.14931, 38.12714, 38.10477, 38.08221, 38.05947, 
    38.03653, 38.01339, 37.99007, 37.96656, 37.94285, 37.91896, 37.89487, 
    37.8706, 37.84613, 37.82148, 37.79664, 37.77161, 37.74638, 37.72098, 
    37.69538, 37.6696, 37.64363, 37.61747, 37.59112, 37.56459, 37.53787, 
    37.51097, 37.48388, 37.45661, 37.42915, 37.4015, 37.37368, 37.34566, 
    37.31747, 37.28909, 37.26052, 37.23178, 37.20285, 37.17374, 37.14445, 
    37.11497, 37.08532, 37.05548, 37.02546, 36.99527, 36.96489, 36.93433, 
    36.90359, 36.87268, 36.84158, 36.81031, 36.77886, 36.74723, 36.71542, 
    36.68344, 36.65128, 36.61894, 36.58643, 36.55374, 36.52087, 36.48783, 
    36.45462, 36.42123,
  32.70815, 32.75626, 32.80423, 32.85205, 32.89974, 32.94728, 32.99469, 
    33.04195, 33.08906, 33.13603, 33.18286, 33.22955, 33.27608, 33.32248, 
    33.36872, 33.41483, 33.46078, 33.50659, 33.55226, 33.59777, 33.64314, 
    33.68836, 33.73343, 33.77835, 33.82312, 33.86775, 33.91222, 33.95654, 
    34.00072, 34.04474, 34.08861, 34.13232, 34.17589, 34.21931, 34.26257, 
    34.30567, 34.34863, 34.39143, 34.43407, 34.47656, 34.5189, 34.56108, 
    34.6031, 34.64497, 34.68668, 34.72823, 34.76963, 34.81087, 34.85195, 
    34.89287, 34.93364, 34.97424, 35.01468, 35.05497, 35.09509, 35.13506, 
    35.17486, 35.2145, 35.25398, 35.2933, 35.33245, 35.37144, 35.41027, 
    35.44894, 35.48744, 35.52578, 35.56395, 35.60196, 35.6398, 35.67748, 
    35.71499, 35.75233, 35.78951, 35.82652, 35.86337, 35.90004, 35.93655, 
    35.97289, 36.00905, 36.04506, 36.08088, 36.11655, 36.15203, 36.18736, 
    36.2225, 36.25748, 36.29229, 36.32692, 36.36138, 36.39567, 36.42978, 
    36.46373, 36.49749, 36.53109, 36.56451, 36.59775, 36.63082, 36.66372, 
    36.69643, 36.72898, 36.76134, 36.79353, 36.82554, 36.85738, 36.88903, 
    36.92051, 36.95181, 36.98294, 37.01388, 37.04464, 37.07523, 37.10563, 
    37.13585, 37.16589, 37.19576, 37.22543, 37.25493, 37.28425, 37.31338, 
    37.34233, 37.3711, 37.39969, 37.42809, 37.45631, 37.48434, 37.51219, 
    37.53986, 37.56734, 37.59463, 37.62174, 37.64866, 37.6754, 37.70195, 
    37.72831, 37.75449, 37.78048, 37.80628, 37.83189, 37.85732, 37.88255, 
    37.9076, 37.93246, 37.95713, 37.98161, 38.0059, 38.03, 38.05391, 
    38.07763, 38.10115, 38.12449, 38.14763, 38.17059, 38.19334, 38.21591, 
    38.23829, 38.26047, 38.28246, 38.30426, 38.32586, 38.34727, 38.36848, 
    38.38951, 38.41033, 38.43096, 38.4514, 38.47164, 38.49168, 38.51154, 
    38.53119, 38.55064, 38.5699, 38.58897, 38.60784, 38.62651, 38.64498, 
    38.66325, 38.68133, 38.69921, 38.71689, 38.73437, 38.75166, 38.76874, 
    38.78563, 38.80231, 38.8188, 38.83509, 38.85118, 38.86707, 38.88275, 
    38.89824, 38.91352, 38.92861, 38.94349, 38.95818, 38.97266, 38.98694, 
    39.00102, 39.0149, 39.02857, 39.04204, 39.05531, 39.06838, 39.08125, 
    39.09391, 39.10637, 39.11863, 39.13068, 39.14252, 39.15417, 39.16562, 
    39.17685, 39.18789, 39.19872, 39.20934, 39.21976, 39.22998, 39.23999, 
    39.2498, 39.2594, 39.2688, 39.27799, 39.28698, 39.29576, 39.30433, 
    39.3127, 39.32087, 39.32883, 39.33658, 39.34413, 39.35147, 39.3586, 
    39.36553, 39.37225, 39.37877, 39.38507, 39.39118, 39.39707, 39.40276, 
    39.40825, 39.41352, 39.41859, 39.42345, 39.4281, 39.43255, 39.43679, 
    39.44082, 39.44464, 39.44826, 39.45167, 39.45488, 39.45787, 39.46066, 
    39.46324, 39.46561, 39.46778, 39.46973, 39.47148, 39.47302, 39.47436, 
    39.47548, 39.4764, 39.47711, 39.47762, 39.47791, 39.478, 39.47788, 
    39.47755, 39.47702, 39.47627, 39.47532, 39.47416, 39.47279, 39.47122, 
    39.46944, 39.46745, 39.46525, 39.46284, 39.46023, 39.45741, 39.45438, 
    39.45115, 39.4477, 39.44405, 39.4402, 39.43613, 39.43186, 39.42738, 
    39.42269, 39.4178, 39.4127, 39.40739, 39.40187, 39.39615, 39.39022, 
    39.38409, 39.37775, 39.3712, 39.36445, 39.35749, 39.35032, 39.34295, 
    39.33537, 39.32758, 39.31959, 39.31139, 39.30299, 39.29438, 39.28557, 
    39.27655, 39.26733, 39.2579, 39.24826, 39.23842, 39.22838, 39.21813, 
    39.20767, 39.19702, 39.18615, 39.17509, 39.16382, 39.15234, 39.14067, 
    39.12878, 39.1167, 39.10441, 39.09192, 39.07922, 39.06633, 39.05323, 
    39.03992, 39.02642, 39.01271, 38.99881, 38.9847, 38.97038, 38.95587, 
    38.94115, 38.92624, 38.91112, 38.8958, 38.88028, 38.86456, 38.84864, 
    38.83253, 38.81621, 38.79969, 38.78297, 38.76605, 38.74894, 38.73162, 
    38.71411, 38.6964, 38.67849, 38.66038, 38.64207, 38.62357, 38.60487, 
    38.58597, 38.56687, 38.54758, 38.52809, 38.50841, 38.48853, 38.46845, 
    38.44818, 38.42771, 38.40705, 38.38619, 38.36514, 38.34389, 38.32246, 
    38.30082, 38.279, 38.25698, 38.23476, 38.21236, 38.18976, 38.16697, 
    38.14399, 38.12081, 38.09744, 38.07389, 38.05014, 38.0262, 38.00207, 
    37.97775, 37.95324, 37.92854, 37.90365, 37.87857, 37.85331, 37.82785, 
    37.80221, 37.77638, 37.75036, 37.72416, 37.69776, 37.67118, 37.64442, 
    37.61746, 37.59032, 37.563, 37.53549, 37.5078, 37.47992, 37.45185, 
    37.42361, 37.39518, 37.36656, 37.33776, 37.30878, 37.27962, 37.25028, 
    37.22075, 37.19104, 37.16115, 37.13108, 37.10083, 37.0704, 37.03979, 
    37.009, 36.97802, 36.94688, 36.91555, 36.88404, 36.85236, 36.82049, 
    36.78845, 36.75623, 36.72384, 36.69127, 36.65852, 36.6256, 36.59251, 
    36.55923, 36.52579,
  32.80655, 32.85474, 32.90277, 32.95068, 32.99843, 33.04605, 33.09352, 
    33.14085, 33.18804, 33.23508, 33.28198, 33.32874, 33.37534, 33.42181, 
    33.46813, 33.5143, 33.56033, 33.6062, 33.65194, 33.69753, 33.74296, 
    33.78825, 33.83339, 33.87838, 33.92323, 33.96792, 34.01246, 34.05685, 
    34.10109, 34.14518, 34.18913, 34.23291, 34.27655, 34.32003, 34.36336, 
    34.40653, 34.44955, 34.49242, 34.53513, 34.57769, 34.62009, 34.66234, 
    34.70443, 34.74637, 34.78815, 34.82977, 34.87123, 34.91254, 34.95368, 
    34.99467, 35.0355, 35.07617, 35.11668, 35.15703, 35.19722, 35.23725, 
    35.27712, 35.31683, 35.35637, 35.39576, 35.43497, 35.47403, 35.51292, 
    35.55165, 35.59022, 35.62862, 35.66686, 35.70493, 35.74284, 35.78057, 
    35.81815, 35.85556, 35.8928, 35.92987, 35.96677, 36.00351, 36.04008, 
    36.07648, 36.11271, 36.14877, 36.18466, 36.22038, 36.25594, 36.29131, 
    36.32652, 36.36156, 36.39642, 36.43112, 36.46564, 36.49998, 36.53416, 
    36.56816, 36.60199, 36.63564, 36.66912, 36.70242, 36.73555, 36.7685, 
    36.80127, 36.83387, 36.86629, 36.89854, 36.93061, 36.9625, 36.99421, 
    37.02575, 37.0571, 37.08828, 37.11928, 37.15009, 37.18073, 37.21119, 
    37.24147, 37.27156, 37.30148, 37.33121, 37.36076, 37.39013, 37.41932, 
    37.44832, 37.47714, 37.50578, 37.53423, 37.5625, 37.59058, 37.61848, 
    37.6462, 37.67373, 37.70107, 37.72823, 37.7552, 37.78199, 37.80858, 
    37.835, 37.86122, 37.88726, 37.91311, 37.93877, 37.96424, 37.98952, 
    38.01461, 38.03952, 38.06423, 38.08876, 38.11309, 38.13723, 38.16119, 
    38.18495, 38.20852, 38.2319, 38.25509, 38.27808, 38.30089, 38.3235, 
    38.34591, 38.36814, 38.39017, 38.41201, 38.43365, 38.4551, 38.47635, 
    38.49741, 38.51828, 38.53895, 38.55942, 38.5797, 38.59978, 38.61967, 
    38.63936, 38.65886, 38.67815, 38.69725, 38.71616, 38.73486, 38.75337, 
    38.77168, 38.78979, 38.8077, 38.82542, 38.84293, 38.86025, 38.87737, 
    38.89429, 38.911, 38.92752, 38.94384, 38.95996, 38.97588, 38.9916, 
    39.00711, 39.02243, 39.03754, 39.05246, 39.06717, 39.08168, 39.09599, 
    39.11009, 39.12399, 39.1377, 39.1512, 39.16449, 39.17758, 39.19047, 
    39.20316, 39.21564, 39.22792, 39.24, 39.25187, 39.26354, 39.275, 
    39.28626, 39.29732, 39.30817, 39.31882, 39.32926, 39.33949, 39.34953, 
    39.35935, 39.36897, 39.37839, 39.3876, 39.3966, 39.4054, 39.41399, 
    39.42238, 39.43056, 39.43853, 39.4463, 39.45387, 39.46122, 39.46837, 
    39.47531, 39.48204, 39.48857, 39.49489, 39.50101, 39.50691, 39.51262, 
    39.51811, 39.52339, 39.52847, 39.53334, 39.538, 39.54246, 39.54671, 
    39.55075, 39.55458, 39.5582, 39.56162, 39.56483, 39.56783, 39.57063, 
    39.57321, 39.57558, 39.57775, 39.57972, 39.58147, 39.58302, 39.58435, 
    39.58548, 39.5864, 39.58711, 39.58762, 39.58791, 39.588, 39.58788, 
    39.58755, 39.58701, 39.58627, 39.58532, 39.58415, 39.58278, 39.58121, 
    39.57942, 39.57743, 39.57523, 39.57281, 39.57019, 39.56737, 39.56433, 
    39.56109, 39.55764, 39.55399, 39.55012, 39.54605, 39.54177, 39.53728, 
    39.53259, 39.52768, 39.52257, 39.51725, 39.51173, 39.50599, 39.50005, 
    39.49391, 39.48755, 39.48099, 39.47422, 39.46725, 39.46007, 39.45268, 
    39.44509, 39.43729, 39.42928, 39.42107, 39.41265, 39.40402, 39.39519, 
    39.38615, 39.37691, 39.36746, 39.35781, 39.34795, 39.33789, 39.32762, 
    39.31715, 39.30647, 39.29558, 39.2845, 39.2732, 39.26171, 39.25001, 
    39.2381, 39.22599, 39.21368, 39.20116, 39.18845, 39.17553, 39.1624, 
    39.14907, 39.13554, 39.12181, 39.10787, 39.09373, 39.0794, 39.06485, 
    39.05011, 39.03516, 39.02002, 39.00467, 38.98912, 38.97337, 38.95742, 
    38.94127, 38.92492, 38.90837, 38.89162, 38.87467, 38.85752, 38.84018, 
    38.82263, 38.80488, 38.78694, 38.7688, 38.75045, 38.73191, 38.71318, 
    38.69424, 38.67511, 38.65578, 38.63626, 38.61654, 38.59662, 38.57651, 
    38.5562, 38.53569, 38.51499, 38.49409, 38.473, 38.45172, 38.43024, 
    38.40857, 38.3867, 38.36464, 38.34238, 38.31993, 38.29729, 38.27446, 
    38.25143, 38.22821, 38.20481, 38.18121, 38.15741, 38.13343, 38.10925, 
    38.08489, 38.06034, 38.03559, 38.01065, 37.98553, 37.96022, 37.93472, 
    37.90903, 37.88315, 37.85708, 37.83083, 37.80439, 37.77776, 37.75095, 
    37.72395, 37.69676, 37.66938, 37.64183, 37.61408, 37.58615, 37.55804, 
    37.52974, 37.50126, 37.47259, 37.44374, 37.41471, 37.38549, 37.3561, 
    37.32652, 37.29676, 37.26681, 37.23669, 37.20638, 37.1759, 37.14523, 
    37.11439, 37.08336, 37.05215, 37.02077, 36.98921, 36.95747, 36.92555, 
    36.89345, 36.86118, 36.82873, 36.7961, 36.7633, 36.73032, 36.69716, 
    36.66383, 36.63033,
  32.90493, 32.95319, 33.0013, 33.04927, 33.0971, 33.14479, 33.19233, 
    33.23973, 33.28699, 33.3341, 33.38107, 33.4279, 33.47458, 33.52111, 
    33.5675, 33.61375, 33.65984, 33.70579, 33.75159, 33.79725, 33.84276, 
    33.88812, 33.93333, 33.97839, 34.0233, 34.06807, 34.11268, 34.15714, 
    34.20145, 34.24561, 34.28962, 34.33347, 34.37717, 34.42073, 34.46412, 
    34.50737, 34.55046, 34.59339, 34.63617, 34.6788, 34.72127, 34.76358, 
    34.80574, 34.84775, 34.88959, 34.93128, 34.97281, 35.01418, 35.0554, 
    35.09645, 35.13735, 35.17809, 35.21866, 35.25908, 35.29933, 35.33943, 
    35.37936, 35.41913, 35.45874, 35.49819, 35.53748, 35.5766, 35.61555, 
    35.65435, 35.69298, 35.73145, 35.76974, 35.80788, 35.84585, 35.88365, 
    35.92129, 35.95876, 35.99606, 36.0332, 36.07016, 36.10696, 36.14359, 
    36.18005, 36.21635, 36.25247, 36.28842, 36.3242, 36.35982, 36.39526, 
    36.43053, 36.46562, 36.50055, 36.5353, 36.56988, 36.60429, 36.63852, 
    36.67258, 36.70647, 36.74018, 36.77371, 36.80707, 36.84026, 36.87327, 
    36.9061, 36.93876, 36.97124, 37.00354, 37.03566, 37.06761, 37.09938, 
    37.13097, 37.16238, 37.19361, 37.22466, 37.25554, 37.28623, 37.31674, 
    37.34707, 37.37722, 37.40718, 37.43697, 37.46658, 37.496, 37.52524, 
    37.55429, 37.58316, 37.61185, 37.64036, 37.66868, 37.69681, 37.72476, 
    37.75253, 37.78011, 37.8075, 37.83471, 37.86173, 37.88856, 37.91521, 
    37.94167, 37.96794, 37.99403, 38.01992, 38.04563, 38.07115, 38.09648, 
    38.12162, 38.14657, 38.17133, 38.1959, 38.22028, 38.24446, 38.26846, 
    38.29227, 38.31588, 38.33931, 38.36254, 38.38557, 38.40842, 38.43107, 
    38.45353, 38.4758, 38.49787, 38.51975, 38.54143, 38.56292, 38.58422, 
    38.60532, 38.62622, 38.64693, 38.66744, 38.68776, 38.70788, 38.7278, 
    38.74753, 38.76706, 38.7864, 38.80553, 38.82447, 38.84321, 38.86176, 
    38.8801, 38.89824, 38.91619, 38.93394, 38.95149, 38.96884, 38.98599, 
    39.00294, 39.01969, 39.03624, 39.05259, 39.06874, 39.08469, 39.10044, 
    39.11598, 39.13133, 39.14647, 39.16141, 39.17615, 39.19069, 39.20502, 
    39.21916, 39.23309, 39.24682, 39.26034, 39.27366, 39.28678, 39.2997, 
    39.31241, 39.32492, 39.33722, 39.34932, 39.36121, 39.37291, 39.38439, 
    39.39567, 39.40675, 39.41762, 39.42829, 39.43875, 39.44901, 39.45906, 
    39.4689, 39.47854, 39.48798, 39.4972, 39.50623, 39.51504, 39.52365, 
    39.53205, 39.54025, 39.54824, 39.55602, 39.5636, 39.57097, 39.57813, 
    39.58509, 39.59184, 39.59838, 39.60471, 39.61084, 39.61676, 39.62247, 
    39.62797, 39.63327, 39.63835, 39.64323, 39.6479, 39.65237, 39.65662, 
    39.66068, 39.66451, 39.66814, 39.67157, 39.67479, 39.67779, 39.68059, 
    39.68318, 39.68556, 39.68774, 39.6897, 39.69146, 39.693, 39.69434, 
    39.69547, 39.6964, 39.69711, 39.69762, 39.69791, 39.698, 39.69788, 
    39.69755, 39.69701, 39.69627, 39.69531, 39.69415, 39.69277, 39.69119, 
    39.6894, 39.6874, 39.6852, 39.68279, 39.68016, 39.67733, 39.67429, 
    39.67104, 39.66758, 39.66392, 39.66005, 39.65597, 39.65168, 39.64718, 
    39.64248, 39.63756, 39.63244, 39.62711, 39.62157, 39.61583, 39.60988, 
    39.60372, 39.59735, 39.59078, 39.584, 39.57701, 39.56982, 39.56242, 
    39.55481, 39.54699, 39.53897, 39.53074, 39.5223, 39.51366, 39.50481, 
    39.49576, 39.4865, 39.47703, 39.46736, 39.45748, 39.4474, 39.43711, 
    39.42662, 39.41592, 39.40501, 39.3939, 39.38259, 39.37107, 39.35934, 
    39.34742, 39.33529, 39.32295, 39.31041, 39.29767, 39.28472, 39.27157, 
    39.25822, 39.24466, 39.2309, 39.21694, 39.20277, 39.1884, 39.17384, 
    39.15906, 39.14409, 39.12891, 39.11354, 39.09796, 39.08218, 39.0662, 
    39.05002, 39.03363, 39.01706, 39.00027, 38.98329, 38.96611, 38.94873, 
    38.93114, 38.91336, 38.89539, 38.87721, 38.85883, 38.84026, 38.82149, 
    38.80252, 38.78335, 38.76398, 38.74442, 38.72467, 38.70471, 38.68456, 
    38.66421, 38.64367, 38.62292, 38.60199, 38.58086, 38.55954, 38.53801, 
    38.5163, 38.49439, 38.47229, 38.44999, 38.4275, 38.40482, 38.38194, 
    38.35888, 38.33561, 38.31216, 38.28852, 38.26468, 38.24065, 38.21643, 
    38.19202, 38.16742, 38.14263, 38.11765, 38.09248, 38.06712, 38.04158, 
    38.01584, 37.98991, 37.9638, 37.9375, 37.91101, 37.88433, 37.85747, 
    37.83042, 37.80318, 37.77576, 37.74815, 37.72035, 37.69238, 37.66421, 
    37.63586, 37.60733, 37.57861, 37.54971, 37.52062, 37.49136, 37.46191, 
    37.43227, 37.40246, 37.37246, 37.34229, 37.31192, 37.28138, 37.25066, 
    37.21976, 37.18868, 37.15742, 37.12598, 37.09436, 37.06257, 37.03059, 
    36.99844, 36.96611, 36.9336, 36.90092, 36.86806, 36.83502, 36.80181, 
    36.76842, 36.73486,
  33.00328, 33.05161, 33.09979, 33.14783, 33.19574, 33.2435, 33.29111, 
    33.33858, 33.38591, 33.4331, 33.48014, 33.52703, 33.57379, 33.62039, 
    33.66685, 33.71317, 33.75933, 33.80536, 33.85123, 33.89695, 33.94253, 
    33.98796, 34.03324, 34.07837, 34.12336, 34.16819, 34.21287, 34.2574, 
    34.30178, 34.34601, 34.39008, 34.43401, 34.47778, 34.5214, 34.56487, 
    34.60818, 34.65134, 34.69434, 34.73719, 34.77988, 34.82243, 34.86481, 
    34.90703, 34.9491, 34.99102, 35.03277, 35.07437, 35.11581, 35.15709, 
    35.19821, 35.23917, 35.27998, 35.32062, 35.3611, 35.40142, 35.44158, 
    35.48158, 35.52142, 35.5611, 35.60061, 35.63996, 35.67914, 35.71817, 
    35.75702, 35.79572, 35.83425, 35.87261, 35.91081, 35.94884, 35.98671, 
    36.02441, 36.06194, 36.09931, 36.13651, 36.17353, 36.2104, 36.24709, 
    36.28362, 36.31997, 36.35615, 36.39217, 36.42801, 36.46368, 36.49918, 
    36.53451, 36.56967, 36.60466, 36.63947, 36.67411, 36.70857, 36.74287, 
    36.77699, 36.81093, 36.8447, 36.87829, 36.91171, 36.94495, 36.97802, 
    37.01091, 37.04362, 37.07616, 37.10852, 37.1407, 37.1727, 37.20453, 
    37.23618, 37.26764, 37.29893, 37.33004, 37.36096, 37.39171, 37.42228, 
    37.45266, 37.48286, 37.51288, 37.54272, 37.57238, 37.60186, 37.63115, 
    37.66025, 37.68918, 37.71792, 37.74647, 37.77485, 37.80303, 37.83103, 
    37.85885, 37.88648, 37.91392, 37.94118, 37.96825, 37.99513, 38.02183, 
    38.04833, 38.07465, 38.10078, 38.12673, 38.15248, 38.17805, 38.20343, 
    38.22861, 38.25361, 38.27841, 38.30303, 38.32745, 38.35169, 38.37573, 
    38.39958, 38.42324, 38.4467, 38.46998, 38.49306, 38.51595, 38.53864, 
    38.56114, 38.58345, 38.60556, 38.62748, 38.64921, 38.67074, 38.69207, 
    38.71321, 38.73415, 38.7549, 38.77546, 38.79581, 38.81597, 38.83593, 
    38.85569, 38.87526, 38.89463, 38.91381, 38.93278, 38.95156, 38.97013, 
    38.98851, 39.00669, 39.02468, 39.04246, 39.06004, 39.07742, 39.09461, 
    39.11159, 39.12837, 39.14495, 39.16133, 39.17752, 39.19349, 39.20927, 
    39.22485, 39.24022, 39.25539, 39.27037, 39.28513, 39.2997, 39.31406, 
    39.32822, 39.34218, 39.35593, 39.36949, 39.38284, 39.39598, 39.40892, 
    39.42165, 39.43419, 39.44651, 39.45864, 39.47055, 39.48227, 39.49378, 
    39.50508, 39.51618, 39.52707, 39.53776, 39.54824, 39.55852, 39.56859, 
    39.57845, 39.58811, 39.59756, 39.60681, 39.61585, 39.62468, 39.63331, 
    39.64173, 39.64994, 39.65795, 39.66574, 39.67334, 39.68072, 39.6879, 
    39.69487, 39.70163, 39.70818, 39.71453, 39.72066, 39.72659, 39.73232, 
    39.73783, 39.74314, 39.74823, 39.75312, 39.7578, 39.76228, 39.76654, 
    39.7706, 39.77445, 39.77809, 39.78152, 39.78474, 39.78775, 39.79055, 
    39.79315, 39.79554, 39.79771, 39.79968, 39.80145, 39.80299, 39.80434, 
    39.80547, 39.80639, 39.80711, 39.80761, 39.80791, 39.808, 39.80788, 
    39.80755, 39.80701, 39.80626, 39.80531, 39.80414, 39.80276, 39.80118, 
    39.79939, 39.79739, 39.79517, 39.79276, 39.79013, 39.78729, 39.78424, 
    39.78099, 39.77752, 39.77385, 39.76997, 39.76588, 39.76159, 39.75708, 
    39.75237, 39.74744, 39.74231, 39.73697, 39.73143, 39.72567, 39.71971, 
    39.71354, 39.70716, 39.70057, 39.69378, 39.68678, 39.67957, 39.67215, 
    39.66452, 39.65669, 39.64865, 39.64041, 39.63196, 39.6233, 39.61443, 
    39.60536, 39.59608, 39.5866, 39.57691, 39.56701, 39.55691, 39.5466, 
    39.53608, 39.52536, 39.51444, 39.50331, 39.49197, 39.48043, 39.46868, 
    39.45673, 39.44458, 39.43222, 39.41965, 39.40688, 39.39391, 39.38074, 
    39.36736, 39.35378, 39.33999, 39.326, 39.31181, 39.29741, 39.28281, 
    39.26801, 39.25301, 39.2378, 39.2224, 39.20679, 39.19098, 39.17497, 
    39.15876, 39.14235, 39.12573, 39.10892, 39.0919, 39.07469, 39.05727, 
    39.03966, 39.02184, 39.00383, 38.98562, 38.96721, 38.9486, 38.92979, 
    38.91079, 38.89158, 38.87218, 38.85258, 38.83279, 38.81279, 38.7926, 
    38.77222, 38.75163, 38.73085, 38.70988, 38.68871, 38.66734, 38.64578, 
    38.62403, 38.60208, 38.57993, 38.5576, 38.53506, 38.51234, 38.48942, 
    38.46631, 38.443, 38.41951, 38.39582, 38.37194, 38.34787, 38.3236, 
    38.29915, 38.2745, 38.24967, 38.22464, 38.19942, 38.17402, 38.14842, 
    38.12264, 38.09666, 38.0705, 38.04416, 38.01762, 37.99089, 37.96398, 
    37.93688, 37.90959, 37.88212, 37.85446, 37.82661, 37.79858, 37.77037, 
    37.74197, 37.71338, 37.68462, 37.65566, 37.62653, 37.59721, 37.5677, 
    37.53802, 37.50815, 37.4781, 37.44786, 37.41745, 37.38686, 37.35608, 
    37.32513, 37.29399, 37.26268, 37.23118, 37.1995, 37.16765, 37.13562, 
    37.10341, 37.07103, 37.03846, 37.00572, 36.9728, 36.93971, 36.90644, 
    36.87299, 36.83937,
  33.10161, 33.15001, 33.19826, 33.24638, 33.29435, 33.34218, 33.38987, 
    33.43741, 33.48481, 33.53207, 33.57918, 33.62614, 33.67297, 33.71965, 
    33.76617, 33.81256, 33.8588, 33.90489, 33.95083, 33.99663, 34.04228, 
    34.08778, 34.13313, 34.17833, 34.22338, 34.26828, 34.31303, 34.35764, 
    34.40208, 34.44638, 34.49053, 34.53452, 34.57837, 34.62206, 34.66559, 
    34.70897, 34.7522, 34.79527, 34.83818, 34.88095, 34.92355, 34.966, 
    35.0083, 35.05044, 35.09241, 35.13424, 35.1759, 35.21741, 35.25876, 
    35.29995, 35.34098, 35.38184, 35.42255, 35.4631, 35.50349, 35.54372, 
    35.58378, 35.62368, 35.66343, 35.703, 35.74242, 35.78167, 35.82076, 
    35.85968, 35.89844, 35.93703, 35.97546, 36.01372, 36.05182, 36.08975, 
    36.12751, 36.16511, 36.20254, 36.2398, 36.27689, 36.31381, 36.35057, 
    36.38715, 36.42357, 36.45982, 36.49589, 36.5318, 36.56753, 36.60309, 
    36.63848, 36.6737, 36.70874, 36.74362, 36.77832, 36.81284, 36.84719, 
    36.88137, 36.91537, 36.9492, 36.98286, 37.01633, 37.04963, 37.08276, 
    37.11571, 37.14848, 37.18107, 37.21349, 37.24573, 37.27779, 37.30967, 
    37.34137, 37.37289, 37.40423, 37.43539, 37.46638, 37.49718, 37.5278, 
    37.55824, 37.58849, 37.61857, 37.64846, 37.67817, 37.7077, 37.73704, 
    37.7662, 37.79518, 37.82397, 37.85258, 37.881, 37.90924, 37.93729, 
    37.96516, 37.99284, 38.02033, 38.04763, 38.07476, 38.10169, 38.12843, 
    38.15499, 38.18136, 38.20753, 38.23353, 38.25933, 38.28494, 38.31036, 
    38.3356, 38.36064, 38.38549, 38.41015, 38.43462, 38.4589, 38.48299, 
    38.50688, 38.53058, 38.55409, 38.57741, 38.60054, 38.62347, 38.6462, 
    38.66875, 38.6911, 38.71325, 38.73521, 38.75698, 38.77855, 38.79992, 
    38.8211, 38.84208, 38.86287, 38.88346, 38.90385, 38.92405, 38.94405, 
    38.96385, 38.98346, 39.00286, 39.02208, 39.04108, 39.0599, 39.07851, 
    39.09692, 39.11514, 39.13316, 39.15097, 39.16859, 39.186, 39.20322, 
    39.22023, 39.23705, 39.25366, 39.27008, 39.28629, 39.3023, 39.3181, 
    39.33371, 39.34912, 39.36432, 39.37932, 39.39412, 39.40871, 39.4231, 
    39.43729, 39.45127, 39.46505, 39.47863, 39.492, 39.50517, 39.51814, 
    39.5309, 39.54345, 39.55581, 39.56795, 39.57989, 39.59163, 39.60316, 
    39.61449, 39.62561, 39.63652, 39.64723, 39.65773, 39.66803, 39.67812, 
    39.688, 39.69768, 39.70715, 39.71642, 39.72547, 39.73432, 39.74297, 
    39.7514, 39.75963, 39.76765, 39.77546, 39.78307, 39.79047, 39.79766, 
    39.80464, 39.81142, 39.81798, 39.82434, 39.83049, 39.83643, 39.84217, 
    39.84769, 39.85301, 39.85812, 39.86302, 39.86771, 39.87219, 39.87646, 
    39.88053, 39.88438, 39.88803, 39.89146, 39.89469, 39.89771, 39.90052, 
    39.90312, 39.90551, 39.9077, 39.90967, 39.91143, 39.91298, 39.91433, 
    39.91546, 39.91639, 39.91711, 39.91761, 39.91791, 39.918, 39.91788, 
    39.91755, 39.91701, 39.91626, 39.9153, 39.91413, 39.91275, 39.91117, 
    39.90937, 39.90736, 39.90515, 39.90273, 39.90009, 39.89725, 39.8942, 
    39.89093, 39.88747, 39.88379, 39.8799, 39.8758, 39.87149, 39.86698, 
    39.86226, 39.85732, 39.85218, 39.84683, 39.84127, 39.83551, 39.82953, 
    39.82335, 39.81696, 39.81036, 39.80355, 39.79654, 39.78931, 39.78188, 
    39.77424, 39.7664, 39.75834, 39.75008, 39.74161, 39.73294, 39.72405, 
    39.71496, 39.70567, 39.69616, 39.68645, 39.67654, 39.66641, 39.65609, 
    39.64555, 39.63481, 39.62386, 39.61271, 39.60135, 39.58979, 39.57802, 
    39.56604, 39.55386, 39.54148, 39.52889, 39.5161, 39.5031, 39.4899, 
    39.47649, 39.46289, 39.44907, 39.43505, 39.42084, 39.40641, 39.39179, 
    39.37696, 39.36193, 39.34669, 39.33126, 39.31562, 39.29978, 39.28374, 
    39.26749, 39.25105, 39.2344, 39.21756, 39.20051, 39.18326, 39.16581, 
    39.14817, 39.13032, 39.11227, 39.09402, 39.07558, 39.05693, 39.03809, 
    39.01905, 38.99981, 38.98037, 38.96074, 38.9409, 38.92087, 38.90064, 
    38.88021, 38.8596, 38.83878, 38.81776, 38.79655, 38.77515, 38.75355, 
    38.73175, 38.70976, 38.68757, 38.66519, 38.64262, 38.61985, 38.59689, 
    38.57373, 38.55039, 38.52685, 38.50312, 38.47919, 38.45507, 38.43076, 
    38.40627, 38.38157, 38.35669, 38.33162, 38.30635, 38.2809, 38.25526, 
    38.22943, 38.20341, 38.1772, 38.1508, 38.12421, 38.09744, 38.07048, 
    38.04333, 38.01599, 37.98847, 37.96076, 37.93287, 37.90479, 37.87652, 
    37.84806, 37.81943, 37.79061, 37.7616, 37.73241, 37.70304, 37.67348, 
    37.64375, 37.61382, 37.58372, 37.55343, 37.52297, 37.49232, 37.46149, 
    37.43048, 37.39928, 37.36792, 37.33636, 37.30463, 37.27272, 37.24064, 
    37.20837, 37.17593, 37.14331, 37.11051, 37.07753, 37.04438, 37.01105, 
    36.97755, 36.94387,
  33.19991, 33.24837, 33.2967, 33.34489, 33.39293, 33.44083, 33.48859, 
    33.53621, 33.58368, 33.63101, 33.67819, 33.72523, 33.77213, 33.81887, 
    33.86547, 33.91193, 33.95824, 34.0044, 34.05042, 34.09628, 34.142, 
    34.18757, 34.23299, 34.27826, 34.32338, 34.36835, 34.41318, 34.45785, 
    34.50237, 34.54673, 34.59095, 34.63501, 34.67892, 34.72268, 34.76628, 
    34.80973, 34.85303, 34.89617, 34.93916, 34.98199, 35.02466, 35.06718, 
    35.10954, 35.15175, 35.19379, 35.23569, 35.27742, 35.31899, 35.3604, 
    35.40166, 35.44276, 35.48369, 35.52447, 35.56509, 35.60554, 35.64583, 
    35.68596, 35.72593, 35.76574, 35.80538, 35.84486, 35.88417, 35.92333, 
    35.96231, 36.00114, 36.0398, 36.07829, 36.11662, 36.15478, 36.19277, 
    36.2306, 36.26826, 36.30575, 36.34307, 36.38023, 36.41721, 36.45403, 
    36.49068, 36.52716, 36.56346, 36.5996, 36.63557, 36.67136, 36.70699, 
    36.74244, 36.77771, 36.81282, 36.84775, 36.88251, 36.9171, 36.95151, 
    36.98574, 37.01981, 37.0537, 37.08741, 37.12094, 37.1543, 37.18748, 
    37.22049, 37.25332, 37.28597, 37.31844, 37.35073, 37.38285, 37.41479, 
    37.44654, 37.47812, 37.50952, 37.54074, 37.57178, 37.60263, 37.63331, 
    37.6638, 37.69411, 37.72424, 37.75419, 37.78395, 37.81353, 37.84293, 
    37.87214, 37.90117, 37.93001, 37.95867, 37.98714, 38.01543, 38.04354, 
    38.07145, 38.09918, 38.12673, 38.15408, 38.18125, 38.20823, 38.23503, 
    38.26163, 38.28805, 38.31428, 38.34032, 38.36617, 38.39183, 38.41729, 
    38.44257, 38.46766, 38.49256, 38.51727, 38.54178, 38.5661, 38.59024, 
    38.61417, 38.63792, 38.66148, 38.68484, 38.708, 38.73098, 38.75376, 
    38.77634, 38.79873, 38.82093, 38.84293, 38.86474, 38.88635, 38.90776, 
    38.92898, 38.95, 38.97083, 38.99146, 39.01189, 39.03213, 39.05217, 
    39.07201, 39.09165, 39.11109, 39.13034, 39.14938, 39.16823, 39.18688, 
    39.20533, 39.22358, 39.24163, 39.25948, 39.27713, 39.29458, 39.31183, 
    39.32888, 39.34572, 39.36237, 39.37881, 39.39505, 39.41109, 39.42693, 
    39.44257, 39.458, 39.47324, 39.48827, 39.50309, 39.51771, 39.53213, 
    39.54634, 39.56036, 39.57417, 39.58777, 39.60117, 39.61436, 39.62735, 
    39.64014, 39.65272, 39.66509, 39.67727, 39.68923, 39.70099, 39.71254, 
    39.72389, 39.73503, 39.74597, 39.7567, 39.76722, 39.77754, 39.78765, 
    39.79755, 39.80725, 39.81673, 39.82602, 39.83509, 39.84396, 39.85262, 
    39.86107, 39.86932, 39.87735, 39.88519, 39.8928, 39.90022, 39.90742, 
    39.91442, 39.92121, 39.92779, 39.93416, 39.94032, 39.94627, 39.95202, 
    39.95755, 39.96288, 39.968, 39.97291, 39.97761, 39.9821, 39.98638, 
    39.99045, 39.99432, 39.99797, 40.00141, 40.00465, 40.00767, 40.01049, 
    40.01309, 40.01549, 40.01767, 40.01965, 40.02142, 40.02298, 40.02432, 
    40.02546, 40.02639, 40.0271, 40.02761, 40.02791, 40.028, 40.02788, 
    40.02755, 40.027, 40.02625, 40.0253, 40.02412, 40.02274, 40.02115, 
    40.01935, 40.01734, 40.01512, 40.0127, 40.01006, 40.00721, 40.00415, 
    40.00088, 39.99741, 39.99372, 39.98982, 39.98572, 39.9814, 39.97688, 
    39.97215, 39.96721, 39.96205, 39.95669, 39.95112, 39.94535, 39.93936, 
    39.93316, 39.92676, 39.92015, 39.91333, 39.9063, 39.89906, 39.89161, 
    39.88396, 39.8761, 39.86803, 39.85975, 39.85126, 39.84257, 39.83367, 
    39.82456, 39.81525, 39.80573, 39.796, 39.78606, 39.77592, 39.76557, 
    39.75501, 39.74425, 39.73328, 39.72211, 39.71073, 39.69914, 39.68735, 
    39.67535, 39.66315, 39.65074, 39.63813, 39.62531, 39.61229, 39.59906, 
    39.58563, 39.57199, 39.55816, 39.54411, 39.52987, 39.51541, 39.50076, 
    39.4859, 39.47084, 39.45558, 39.44011, 39.42444, 39.40857, 39.3925, 
    39.37622, 39.35975, 39.34307, 39.32619, 39.30911, 39.29183, 39.27435, 
    39.25667, 39.23879, 39.22071, 39.20242, 39.18394, 39.16526, 39.14639, 
    39.1273, 39.10803, 39.08855, 39.06888, 39.04901, 39.02894, 39.00867, 
    38.98821, 38.96755, 38.94669, 38.92564, 38.90439, 38.88294, 38.8613, 
    38.83947, 38.81743, 38.7952, 38.77278, 38.75017, 38.72736, 38.70435, 
    38.68116, 38.65776, 38.63418, 38.6104, 38.58643, 38.56227, 38.53792, 
    38.51337, 38.48864, 38.46371, 38.43859, 38.41328, 38.38778, 38.36209, 
    38.33621, 38.31014, 38.28388, 38.25744, 38.2308, 38.20398, 38.17697, 
    38.14977, 38.12238, 38.09481, 38.06705, 38.0391, 38.01097, 37.98265, 
    37.95415, 37.92546, 37.89659, 37.86753, 37.83829, 37.80886, 37.77925, 
    37.74946, 37.71949, 37.68933, 37.65899, 37.62847, 37.59776, 37.56688, 
    37.53582, 37.50457, 37.47314, 37.44154, 37.40975, 37.37778, 37.34564, 
    37.31332, 37.28082, 37.24813, 37.21528, 37.18225, 37.14904, 37.11565, 
    37.08208, 37.04835,
  33.29817, 33.34671, 33.39511, 33.44337, 33.49149, 33.53946, 33.58729, 
    33.63498, 33.68252, 33.72992, 33.77718, 33.82429, 33.87125, 33.91807, 
    33.96474, 34.01127, 34.05765, 34.10389, 34.14997, 34.19591, 34.2417, 
    34.28734, 34.33283, 34.37817, 34.42336, 34.4684, 34.51329, 34.55804, 
    34.60262, 34.64706, 34.69135, 34.73548, 34.77946, 34.82328, 34.86696, 
    34.91048, 34.95384, 34.99705, 35.0401, 35.083, 35.12575, 35.16833, 
    35.21076, 35.25304, 35.29515, 35.33711, 35.37891, 35.42055, 35.46203, 
    35.50335, 35.54452, 35.58552, 35.62636, 35.66705, 35.70757, 35.74792, 
    35.78812, 35.82816, 35.86803, 35.90773, 35.94728, 35.98666, 36.02588, 
    36.06493, 36.10382, 36.14254, 36.1811, 36.21949, 36.25771, 36.29577, 
    36.33366, 36.37138, 36.40894, 36.44633, 36.48354, 36.52059, 36.55747, 
    36.59418, 36.63072, 36.66709, 36.70329, 36.73932, 36.77517, 36.81086, 
    36.84637, 36.88171, 36.91688, 36.95187, 36.98669, 37.02134, 37.05581, 
    37.0901, 37.12423, 37.15817, 37.19194, 37.22553, 37.25895, 37.29219, 
    37.32526, 37.35814, 37.39085, 37.42338, 37.45573, 37.4879, 37.5199, 
    37.55171, 37.58335, 37.6148, 37.64607, 37.67717, 37.70808, 37.73881, 
    37.76935, 37.79972, 37.8299, 37.8599, 37.88972, 37.91935, 37.9488, 
    37.97807, 38.00715, 38.03605, 38.06475, 38.09328, 38.12162, 38.14977, 
    38.17774, 38.20552, 38.23312, 38.26052, 38.28774, 38.31477, 38.34161, 
    38.36827, 38.39473, 38.42101, 38.44709, 38.47299, 38.4987, 38.52422, 
    38.54954, 38.57468, 38.59962, 38.62437, 38.64893, 38.6733, 38.69748, 
    38.72146, 38.74525, 38.76885, 38.79226, 38.81546, 38.83848, 38.86131, 
    38.88393, 38.90636, 38.9286, 38.95065, 38.97249, 38.99414, 39.0156, 
    39.03686, 39.05792, 39.07878, 39.09945, 39.11993, 39.1402, 39.16027, 
    39.18015, 39.19983, 39.21931, 39.23859, 39.25768, 39.27656, 39.29525, 
    39.31373, 39.33202, 39.3501, 39.36798, 39.38567, 39.40315, 39.42043, 
    39.43752, 39.45439, 39.47107, 39.48755, 39.50382, 39.51989, 39.53576, 
    39.55143, 39.56689, 39.58215, 39.59721, 39.61206, 39.62671, 39.64116, 
    39.6554, 39.66944, 39.68328, 39.69691, 39.71033, 39.72355, 39.73657, 
    39.74938, 39.76198, 39.77438, 39.78658, 39.79856, 39.81034, 39.82192, 
    39.83329, 39.84446, 39.85541, 39.86617, 39.87671, 39.88704, 39.89717, 
    39.9071, 39.91681, 39.92632, 39.93562, 39.94471, 39.9536, 39.96228, 
    39.97075, 39.979, 39.98706, 39.9949, 40.00254, 40.00996, 40.01719, 
    40.02419, 40.03099, 40.03759, 40.04397, 40.05015, 40.05611, 40.06187, 
    40.06741, 40.07275, 40.07788, 40.0828, 40.08751, 40.09201, 40.0963, 
    40.10038, 40.10425, 40.10791, 40.11136, 40.1146, 40.11763, 40.12045, 
    40.12306, 40.12546, 40.12766, 40.12963, 40.1314, 40.13297, 40.13432, 
    40.13546, 40.13638, 40.1371, 40.13761, 40.13791, 40.138, 40.13788, 
    40.13755, 40.137, 40.13625, 40.13529, 40.13411, 40.13273, 40.13114, 
    40.12933, 40.12732, 40.1251, 40.12266, 40.12002, 40.11716, 40.1141, 
    40.11083, 40.10735, 40.10365, 40.09975, 40.09563, 40.09131, 40.08678, 
    40.08204, 40.07708, 40.07192, 40.06655, 40.06097, 40.05518, 40.04918, 
    40.04298, 40.03656, 40.02993, 40.0231, 40.01606, 40.0088, 40.00134, 
    39.99368, 39.9858, 39.97771, 39.96942, 39.96091, 39.95221, 39.94329, 
    39.93416, 39.92483, 39.91529, 39.90554, 39.89558, 39.88542, 39.87505, 
    39.86448, 39.85369, 39.8427, 39.83151, 39.82011, 39.80849, 39.79668, 
    39.78466, 39.77243, 39.76, 39.74736, 39.73452, 39.72147, 39.70822, 
    39.69476, 39.6811, 39.66723, 39.65316, 39.63889, 39.62441, 39.60973, 
    39.59484, 39.57975, 39.56446, 39.54896, 39.53326, 39.51736, 39.50126, 
    39.48495, 39.46844, 39.45174, 39.43483, 39.41771, 39.4004, 39.38288, 
    39.36517, 39.34725, 39.32914, 39.31082, 39.2923, 39.27359, 39.25467, 
    39.23556, 39.21624, 39.19673, 39.17702, 39.15711, 39.137, 39.1167, 
    39.0962, 39.0755, 39.0546, 39.03351, 39.01222, 38.99073, 38.96905, 
    38.94717, 38.9251, 38.90283, 38.88036, 38.85771, 38.83485, 38.81181, 
    38.78857, 38.76513, 38.7415, 38.71768, 38.69366, 38.66946, 38.64506, 
    38.62047, 38.59569, 38.57071, 38.54555, 38.52019, 38.49464, 38.46891, 
    38.44298, 38.41687, 38.39056, 38.36406, 38.33738, 38.31051, 38.28345, 
    38.2562, 38.22876, 38.20114, 38.17333, 38.14533, 38.11715, 38.08878, 
    38.06023, 38.03149, 38.00256, 37.97345, 37.94416, 37.91468, 37.88501, 
    37.85517, 37.82514, 37.79493, 37.76453, 37.73396, 37.7032, 37.67226, 
    37.64114, 37.60984, 37.57835, 37.54669, 37.51485, 37.48283, 37.45063, 
    37.41825, 37.38569, 37.35295, 37.32004, 37.28695, 37.25368, 37.22023, 
    37.18661, 37.15281,
  33.39641, 33.44503, 33.4935, 33.54183, 33.59002, 33.63806, 33.68597, 
    33.73372, 33.78134, 33.82881, 33.87614, 33.92332, 33.97036, 34.01725, 
    34.06399, 34.11059, 34.15704, 34.20334, 34.2495, 34.29551, 34.34137, 
    34.38708, 34.43264, 34.47805, 34.52332, 34.56843, 34.61339, 34.6582, 
    34.70286, 34.74736, 34.79172, 34.83592, 34.87997, 34.92387, 34.96761, 
    35.0112, 35.05463, 35.09791, 35.14103, 35.184, 35.22681, 35.26946, 
    35.31196, 35.3543, 35.39649, 35.43851, 35.48038, 35.52209, 35.56364, 
    35.60503, 35.64626, 35.68732, 35.72823, 35.76898, 35.80957, 35.84999, 
    35.89026, 35.93036, 35.97029, 36.01007, 36.04968, 36.08913, 36.12841, 
    36.16753, 36.20648, 36.24527, 36.28389, 36.32235, 36.36063, 36.39875, 
    36.43671, 36.47449, 36.51211, 36.54956, 36.58685, 36.62395, 36.6609, 
    36.69767, 36.73427, 36.77071, 36.80696, 36.84306, 36.87897, 36.91472, 
    36.95029, 36.98569, 37.02092, 37.05597, 37.09085, 37.12556, 37.16009, 
    37.19444, 37.22862, 37.26263, 37.29646, 37.33011, 37.36359, 37.39688, 
    37.43001, 37.46295, 37.49572, 37.52831, 37.56071, 37.59294, 37.62499, 
    37.65686, 37.68855, 37.72006, 37.75139, 37.78254, 37.81351, 37.84429, 
    37.87489, 37.90531, 37.93555, 37.9656, 37.99547, 38.02516, 38.05466, 
    38.08398, 38.11311, 38.14206, 38.17083, 38.1994, 38.22779, 38.256, 
    38.28402, 38.31185, 38.33949, 38.36695, 38.39422, 38.4213, 38.44819, 
    38.47489, 38.5014, 38.52773, 38.55386, 38.57981, 38.60556, 38.63113, 
    38.6565, 38.68168, 38.70667, 38.73147, 38.75608, 38.78049, 38.80471, 
    38.82874, 38.85257, 38.87622, 38.89967, 38.92292, 38.94598, 38.96884, 
    38.99151, 39.01399, 39.03627, 39.05835, 39.08024, 39.10193, 39.12343, 
    39.14473, 39.16583, 39.18673, 39.20744, 39.22795, 39.24826, 39.26838, 
    39.28829, 39.30801, 39.32753, 39.34685, 39.36597, 39.38489, 39.40361, 
    39.42213, 39.44044, 39.45856, 39.47648, 39.4942, 39.51172, 39.52903, 
    39.54615, 39.56306, 39.57977, 39.59628, 39.61258, 39.62868, 39.64458, 
    39.66028, 39.67577, 39.69106, 39.70615, 39.72103, 39.73571, 39.75019, 
    39.76446, 39.77852, 39.79239, 39.80604, 39.81949, 39.83274, 39.84578, 
    39.85861, 39.87124, 39.88367, 39.89589, 39.90789, 39.9197, 39.9313, 
    39.94269, 39.95388, 39.96486, 39.97563, 39.98619, 39.99655, 40.0067, 
    40.01664, 40.02637, 40.0359, 40.04522, 40.05433, 40.06323, 40.07193, 
    40.08041, 40.08869, 40.09676, 40.10462, 40.11227, 40.11971, 40.12695, 
    40.13397, 40.14079, 40.14739, 40.15379, 40.15997, 40.16595, 40.17172, 
    40.17728, 40.18262, 40.18776, 40.19269, 40.19741, 40.20192, 40.20621, 
    40.2103, 40.21418, 40.21785, 40.22131, 40.22455, 40.22759, 40.23042, 
    40.23303, 40.23544, 40.23763, 40.23962, 40.24139, 40.24295, 40.24431, 
    40.24545, 40.24638, 40.2471, 40.24761, 40.24791, 40.248, 40.24788, 
    40.24754, 40.247, 40.24625, 40.24528, 40.24411, 40.24272, 40.24112, 
    40.23932, 40.2373, 40.23507, 40.23263, 40.22998, 40.22712, 40.22405, 
    40.22078, 40.21728, 40.21358, 40.20967, 40.20555, 40.20122, 40.19667, 
    40.19193, 40.18696, 40.18179, 40.17641, 40.17082, 40.16502, 40.15901, 
    40.15279, 40.14636, 40.13972, 40.13287, 40.12582, 40.11855, 40.11107, 
    40.10339, 40.0955, 40.08739, 40.07909, 40.07057, 40.06184, 40.0529, 
    40.04376, 40.03441, 40.02485, 40.01508, 40.00511, 39.99493, 39.98454, 
    39.97394, 39.96313, 39.95212, 39.9409, 39.92948, 39.91785, 39.90601, 
    39.89397, 39.88171, 39.86926, 39.8566, 39.84373, 39.83065, 39.81738, 
    39.80389, 39.7902, 39.77631, 39.76221, 39.74791, 39.7334, 39.71869, 
    39.70378, 39.68866, 39.67334, 39.65781, 39.64208, 39.62615, 39.61002, 
    39.59368, 39.57714, 39.5604, 39.54345, 39.52631, 39.50896, 39.49141, 
    39.47366, 39.45571, 39.43756, 39.41921, 39.40066, 39.3819, 39.36295, 
    39.3438, 39.32446, 39.3049, 39.28516, 39.26521, 39.24506, 39.22472, 
    39.20418, 39.18344, 39.16251, 39.14137, 39.12004, 39.09851, 39.07679, 
    39.05487, 39.03276, 39.01044, 38.98794, 38.96524, 38.94234, 38.91925, 
    38.89597, 38.87249, 38.84882, 38.82495, 38.80089, 38.77664, 38.7522, 
    38.72756, 38.70273, 38.67771, 38.6525, 38.62709, 38.6015, 38.57572, 
    38.54974, 38.52358, 38.49722, 38.47068, 38.44395, 38.41703, 38.38992, 
    38.36262, 38.33513, 38.30746, 38.2796, 38.25155, 38.22332, 38.1949, 
    38.16629, 38.1375, 38.10852, 38.07936, 38.05001, 38.02048, 37.99076, 
    37.96086, 37.93078, 37.90051, 37.87006, 37.83943, 37.80862, 37.77763, 
    37.74645, 37.71509, 37.68355, 37.65183, 37.61993, 37.58786, 37.5556, 
    37.52316, 37.49055, 37.45775, 37.42478, 37.39163, 37.3583, 37.3248, 
    37.29112, 37.25726,
  33.49463, 33.54331, 33.59185, 33.64026, 33.68852, 33.73664, 33.78461, 
    33.83244, 33.88013, 33.92767, 33.97507, 34.02232, 34.06943, 34.11639, 
    34.16321, 34.20988, 34.2564, 34.30278, 34.349, 34.39508, 34.44101, 
    34.48679, 34.53242, 34.57791, 34.62324, 34.66842, 34.71346, 34.75834, 
    34.80307, 34.84764, 34.89207, 34.93634, 34.98046, 35.02442, 35.06823, 
    35.11189, 35.15539, 35.19874, 35.24193, 35.28497, 35.32785, 35.37057, 
    35.41314, 35.45555, 35.4978, 35.53989, 35.58183, 35.6236, 35.66522, 
    35.70668, 35.74797, 35.78911, 35.83009, 35.8709, 35.91155, 35.95205, 
    35.99237, 36.03254, 36.07254, 36.11238, 36.15206, 36.19157, 36.23092, 
    36.2701, 36.30912, 36.34797, 36.38666, 36.42518, 36.46353, 36.50172, 
    36.53973, 36.57759, 36.61527, 36.65278, 36.69012, 36.7273, 36.76431, 
    36.80114, 36.8378, 36.8743, 36.91062, 36.94677, 36.98275, 37.01856, 
    37.05419, 37.08965, 37.12494, 37.16006, 37.195, 37.22976, 37.26435, 
    37.29877, 37.33301, 37.36707, 37.40096, 37.43467, 37.46821, 37.50156, 
    37.53474, 37.56775, 37.60057, 37.63321, 37.66568, 37.69797, 37.73007, 
    37.762, 37.79375, 37.82531, 37.8567, 37.8879, 37.91892, 37.94976, 
    37.98042, 38.01089, 38.04118, 38.07129, 38.10122, 38.13095, 38.16051, 
    38.18988, 38.21907, 38.24807, 38.27689, 38.30552, 38.33396, 38.36221, 
    38.39028, 38.41816, 38.44586, 38.47337, 38.50068, 38.52781, 38.55475, 
    38.5815, 38.60807, 38.63444, 38.66063, 38.68661, 38.71242, 38.73803, 
    38.76345, 38.78868, 38.81371, 38.83856, 38.86321, 38.88767, 38.91193, 
    38.93601, 38.95989, 38.98357, 39.00706, 39.03036, 39.05347, 39.07637, 
    39.09909, 39.1216, 39.14392, 39.16605, 39.18798, 39.20971, 39.23125, 
    39.25259, 39.27373, 39.29468, 39.31542, 39.33597, 39.35632, 39.37648, 
    39.39643, 39.41618, 39.43574, 39.45509, 39.47425, 39.49321, 39.51196, 
    39.53052, 39.54887, 39.56702, 39.58498, 39.60273, 39.62028, 39.63763, 
    39.65477, 39.67172, 39.68846, 39.705, 39.72134, 39.73747, 39.7534, 
    39.76913, 39.78465, 39.79997, 39.81509, 39.83, 39.84471, 39.85921, 
    39.87351, 39.8876, 39.90149, 39.91517, 39.92865, 39.94192, 39.95499, 
    39.96785, 39.9805, 39.99295, 40.00519, 40.01723, 40.02905, 40.04068, 
    40.05209, 40.0633, 40.0743, 40.08509, 40.09568, 40.10605, 40.11622, 
    40.12618, 40.13594, 40.14548, 40.15482, 40.16395, 40.17287, 40.18158, 
    40.19008, 40.19838, 40.20646, 40.21434, 40.222, 40.22946, 40.23671, 
    40.24374, 40.25057, 40.25719, 40.2636, 40.2698, 40.27579, 40.28157, 
    40.28714, 40.29249, 40.29764, 40.30258, 40.30731, 40.31182, 40.31613, 
    40.32023, 40.32412, 40.32779, 40.33125, 40.33451, 40.33755, 40.34038, 
    40.343, 40.34541, 40.34761, 40.3496, 40.35138, 40.35294, 40.3543, 
    40.35545, 40.35638, 40.3571, 40.35761, 40.35791, 40.358, 40.35788, 
    40.35754, 40.357, 40.35624, 40.35528, 40.3541, 40.35271, 40.35111, 
    40.3493, 40.34728, 40.34505, 40.3426, 40.33995, 40.33708, 40.33401, 
    40.33072, 40.32722, 40.32351, 40.3196, 40.31546, 40.31113, 40.30658, 
    40.30182, 40.29684, 40.29166, 40.28627, 40.28067, 40.27485, 40.26883, 
    40.2626, 40.25616, 40.2495, 40.24265, 40.23557, 40.22829, 40.2208, 
    40.2131, 40.2052, 40.19708, 40.18875, 40.18021, 40.17147, 40.16252, 
    40.15336, 40.14399, 40.13441, 40.12462, 40.11463, 40.10443, 40.09402, 
    40.0834, 40.07257, 40.06154, 40.0503, 40.03885, 40.0272, 40.01534, 
    40.00327, 39.99099, 39.97851, 39.96583, 39.95293, 39.93983, 39.92653, 
    39.91302, 39.8993, 39.88538, 39.87126, 39.85693, 39.84239, 39.82765, 
    39.81271, 39.79756, 39.78221, 39.76665, 39.7509, 39.73493, 39.71877, 
    39.7024, 39.68583, 39.66905, 39.65208, 39.6349, 39.61752, 39.59993, 
    39.58215, 39.56417, 39.54598, 39.5276, 39.50901, 39.49022, 39.47123, 
    39.45205, 39.43266, 39.41307, 39.39328, 39.3733, 39.35312, 39.33273, 
    39.31216, 39.29138, 39.2704, 39.24923, 39.22786, 39.20629, 39.18452, 
    39.16256, 39.14041, 39.11806, 39.09551, 39.07276, 39.04982, 39.02669, 
    39.00336, 38.97984, 38.95612, 38.93221, 38.90811, 38.88381, 38.85932, 
    38.83464, 38.80976, 38.7847, 38.75944, 38.73399, 38.70835, 38.68252, 
    38.65649, 38.63028, 38.60388, 38.57729, 38.55051, 38.52353, 38.49638, 
    38.46902, 38.44149, 38.41376, 38.38585, 38.35775, 38.32947, 38.301, 
    38.27234, 38.2435, 38.21447, 38.18525, 38.15585, 38.12626, 38.0965, 
    38.06654, 38.0364, 38.00608, 37.97558, 37.9449, 37.91403, 37.88298, 
    37.85175, 37.82033, 37.78874, 37.75696, 37.72501, 37.69287, 37.66056, 
    37.62806, 37.59539, 37.56254, 37.52951, 37.4963, 37.46291, 37.42935, 
    37.39561, 37.36169,
  33.59281, 33.64157, 33.69019, 33.73866, 33.78699, 33.83518, 33.88323, 
    33.93113, 33.97889, 34.0265, 34.07397, 34.1213, 34.16848, 34.21551, 
    34.2624, 34.30914, 34.35574, 34.40218, 34.44848, 34.49463, 34.54063, 
    34.58648, 34.63219, 34.67774, 34.72314, 34.76839, 34.8135, 34.85845, 
    34.90325, 34.9479, 34.99239, 35.03673, 35.08092, 35.12495, 35.16883, 
    35.21256, 35.25613, 35.29955, 35.34281, 35.38591, 35.42886, 35.47165, 
    35.51429, 35.55677, 35.59909, 35.64125, 35.68325, 35.72509, 35.76678, 
    35.8083, 35.84967, 35.89087, 35.93192, 35.9728, 36.01352, 36.05407, 
    36.09447, 36.1347, 36.17477, 36.21468, 36.25442, 36.294, 36.33341, 
    36.37266, 36.41174, 36.45066, 36.48941, 36.52799, 36.56641, 36.60466, 
    36.64274, 36.68066, 36.7184, 36.75598, 36.79339, 36.83062, 36.86769, 
    36.90459, 36.94132, 36.97787, 37.01426, 37.05047, 37.08651, 37.12238, 
    37.15808, 37.1936, 37.22895, 37.26412, 37.29913, 37.33395, 37.3686, 
    37.40308, 37.43738, 37.4715, 37.50545, 37.53922, 37.57281, 37.60623, 
    37.63947, 37.67252, 37.70541, 37.73811, 37.77063, 37.80297, 37.83514, 
    37.86712, 37.89893, 37.93055, 37.96199, 37.99325, 38.02432, 38.05522, 
    38.08593, 38.11646, 38.1468, 38.17697, 38.20695, 38.23674, 38.26635, 
    38.29577, 38.32501, 38.35406, 38.38293, 38.41161, 38.44011, 38.46841, 
    38.49654, 38.52447, 38.55221, 38.57977, 38.60714, 38.63432, 38.66131, 
    38.68811, 38.71472, 38.74114, 38.76737, 38.79342, 38.81926, 38.84492, 
    38.87039, 38.89566, 38.92075, 38.94564, 38.97033, 38.99484, 39.01915, 
    39.04327, 39.06719, 39.09092, 39.11446, 39.1378, 39.16095, 39.1839, 
    39.20665, 39.22921, 39.25158, 39.27374, 39.29572, 39.31749, 39.33907, 
    39.36045, 39.38163, 39.40261, 39.4234, 39.44398, 39.46437, 39.48457, 
    39.50456, 39.52435, 39.54394, 39.56334, 39.58253, 39.60152, 39.62031, 
    39.6389, 39.65729, 39.67548, 39.69347, 39.71125, 39.72884, 39.74622, 
    39.7634, 39.78038, 39.79715, 39.81372, 39.83009, 39.84625, 39.86222, 
    39.87797, 39.89353, 39.90887, 39.92402, 39.93896, 39.9537, 39.96823, 
    39.98256, 39.99667, 40.01059, 40.0243, 40.0378, 40.0511, 40.06419, 
    40.07708, 40.08976, 40.10223, 40.11449, 40.12655, 40.1384, 40.15005, 
    40.16149, 40.17272, 40.18374, 40.19455, 40.20516, 40.21556, 40.22575, 
    40.23573, 40.2455, 40.25506, 40.26442, 40.27356, 40.2825, 40.29123, 
    40.29975, 40.30806, 40.31616, 40.32405, 40.33173, 40.3392, 40.34647, 
    40.35352, 40.36036, 40.36699, 40.37341, 40.37962, 40.38562, 40.39141, 
    40.397, 40.40236, 40.40752, 40.41247, 40.41721, 40.42173, 40.42605, 
    40.43015, 40.43405, 40.43773, 40.4412, 40.44446, 40.44751, 40.45035, 
    40.45297, 40.45539, 40.45759, 40.45958, 40.46136, 40.46294, 40.46429, 
    40.46544, 40.46637, 40.4671, 40.46761, 40.46791, 40.468, 40.46788, 
    40.46754, 40.467, 40.46624, 40.46527, 40.46409, 40.4627, 40.4611, 
    40.45928, 40.45726, 40.45502, 40.45257, 40.44991, 40.44704, 40.44396, 
    40.44067, 40.43716, 40.43344, 40.42952, 40.42538, 40.42103, 40.41647, 
    40.4117, 40.40672, 40.40153, 40.39613, 40.39051, 40.38469, 40.37865, 
    40.37241, 40.36596, 40.35929, 40.35242, 40.34533, 40.33804, 40.33053, 
    40.32281, 40.31489, 40.30676, 40.29842, 40.28986, 40.2811, 40.27213, 
    40.26295, 40.25356, 40.24397, 40.23416, 40.22415, 40.21392, 40.2035, 
    40.19286, 40.18201, 40.17095, 40.15969, 40.14822, 40.13654, 40.12466, 
    40.11257, 40.10027, 40.08776, 40.07505, 40.06214, 40.04901, 40.03568, 
    40.02214, 40.0084, 39.99445, 39.9803, 39.96594, 39.95138, 39.93661, 
    39.92164, 39.90646, 39.89108, 39.8755, 39.8597, 39.84371, 39.82751, 
    39.81112, 39.79451, 39.7777, 39.7607, 39.74348, 39.72607, 39.70845, 
    39.69064, 39.67262, 39.6544, 39.63597, 39.61735, 39.59853, 39.57951, 
    39.56028, 39.54086, 39.52123, 39.50141, 39.48138, 39.46116, 39.44074, 
    39.42012, 39.39931, 39.37829, 39.35708, 39.33567, 39.31406, 39.29225, 
    39.27025, 39.24805, 39.22566, 39.20307, 39.18028, 39.1573, 39.13412, 
    39.11075, 39.08718, 39.06342, 39.03947, 39.01532, 38.99097, 38.96644, 
    38.94171, 38.91679, 38.89168, 38.86637, 38.84088, 38.81519, 38.78931, 
    38.76324, 38.73698, 38.71053, 38.68388, 38.65705, 38.63003, 38.60282, 
    38.57542, 38.54784, 38.52006, 38.4921, 38.46395, 38.43561, 38.40709, 
    38.37838, 38.34948, 38.3204, 38.29113, 38.26168, 38.23204, 38.20222, 
    38.17221, 38.14202, 38.11164, 38.08109, 38.05034, 38.01942, 37.98832, 
    37.95703, 37.92556, 37.89391, 37.86208, 37.83006, 37.79787, 37.7655, 
    37.73295, 37.70022, 37.66731, 37.63422, 37.60095, 37.56751, 37.53389, 
    37.50009, 37.46611,
  33.69096, 33.7398, 33.78848, 33.83703, 33.88544, 33.9337, 33.98182, 
    34.02979, 34.07763, 34.12531, 34.17285, 34.22025, 34.2675, 34.31461, 
    34.36156, 34.40838, 34.45504, 34.50156, 34.54793, 34.59415, 34.64022, 
    34.68615, 34.73192, 34.77755, 34.82302, 34.86834, 34.91351, 34.95853, 
    35.00341, 35.04812, 35.09269, 35.1371, 35.18135, 35.22546, 35.26941, 
    35.31321, 35.35685, 35.40033, 35.44366, 35.48684, 35.52985, 35.57272, 
    35.61542, 35.65796, 35.70035, 35.74258, 35.78465, 35.82656, 35.86832, 
    35.90991, 35.95134, 35.99261, 36.03372, 36.07467, 36.11546, 36.15608, 
    36.19654, 36.23684, 36.27698, 36.31695, 36.35676, 36.3964, 36.43588, 
    36.4752, 36.51434, 36.55333, 36.59214, 36.63079, 36.66927, 36.70758, 
    36.74573, 36.78371, 36.82152, 36.85916, 36.89663, 36.93393, 36.97106, 
    37.00802, 37.04482, 37.08143, 37.11788, 37.15416, 37.19026, 37.22619, 
    37.26194, 37.29753, 37.33294, 37.36818, 37.40324, 37.43812, 37.47283, 
    37.50737, 37.54173, 37.57591, 37.60992, 37.64375, 37.6774, 37.71088, 
    37.74417, 37.77729, 37.81023, 37.84299, 37.87557, 37.90797, 37.94019, 
    37.97223, 38.00409, 38.03577, 38.06726, 38.09858, 38.12971, 38.16066, 
    38.19143, 38.22202, 38.25241, 38.28263, 38.31266, 38.34251, 38.37217, 
    38.40165, 38.43094, 38.46005, 38.48897, 38.5177, 38.54625, 38.57461, 
    38.60278, 38.63076, 38.65856, 38.68616, 38.71358, 38.74081, 38.76785, 
    38.7947, 38.82137, 38.84784, 38.87411, 38.9002, 38.9261, 38.95181, 
    38.97732, 39.00264, 39.02777, 39.05271, 39.07745, 39.102, 39.12636, 
    39.15052, 39.17449, 39.19827, 39.22184, 39.24523, 39.26842, 39.29141, 
    39.31421, 39.33681, 39.35922, 39.38143, 39.40344, 39.42526, 39.44688, 
    39.4683, 39.48952, 39.51054, 39.53137, 39.55199, 39.57242, 39.59265, 
    39.61268, 39.63251, 39.65214, 39.67157, 39.6908, 39.70983, 39.72866, 
    39.74728, 39.76571, 39.78393, 39.80195, 39.81977, 39.83739, 39.8548, 
    39.87202, 39.88903, 39.90583, 39.92244, 39.93884, 39.95503, 39.97103, 
    39.98681, 40.0024, 40.01778, 40.03295, 40.04792, 40.06269, 40.07724, 
    40.0916, 40.10575, 40.11969, 40.13343, 40.14696, 40.16028, 40.1734, 
    40.18631, 40.19901, 40.21151, 40.2238, 40.23588, 40.24775, 40.25942, 
    40.27088, 40.28213, 40.29317, 40.30401, 40.31464, 40.32505, 40.33527, 
    40.34527, 40.35506, 40.36464, 40.37402, 40.38318, 40.39214, 40.40088, 
    40.40942, 40.41774, 40.42586, 40.43377, 40.44146, 40.44895, 40.45622, 
    40.46329, 40.47015, 40.47679, 40.48322, 40.48945, 40.49546, 40.50126, 
    40.50686, 40.51223, 40.5174, 40.52236, 40.52711, 40.53164, 40.53596, 
    40.54008, 40.54398, 40.54767, 40.55115, 40.55441, 40.55747, 40.56031, 
    40.56294, 40.56536, 40.56757, 40.56957, 40.57135, 40.57293, 40.57428, 
    40.57544, 40.57637, 40.5771, 40.57761, 40.57791, 40.578, 40.57788, 
    40.57754, 40.577, 40.57624, 40.57527, 40.57409, 40.57269, 40.57108, 
    40.56927, 40.56724, 40.56499, 40.56254, 40.55988, 40.557, 40.55391, 
    40.55061, 40.5471, 40.54338, 40.53944, 40.5353, 40.53094, 40.52637, 
    40.52159, 40.5166, 40.5114, 40.50598, 40.50036, 40.49452, 40.48848, 
    40.48222, 40.47575, 40.46907, 40.46218, 40.45509, 40.44778, 40.44026, 
    40.43253, 40.42459, 40.41644, 40.40808, 40.39951, 40.39073, 40.38174, 
    40.37255, 40.36314, 40.35352, 40.3437, 40.33366, 40.32342, 40.31297, 
    40.30231, 40.29144, 40.28036, 40.26908, 40.25759, 40.24589, 40.23398, 
    40.22187, 40.20955, 40.19701, 40.18428, 40.17134, 40.15818, 40.14483, 
    40.13127, 40.1175, 40.10352, 40.08934, 40.07495, 40.06036, 40.04557, 
    40.03056, 40.01536, 39.99995, 39.98433, 39.96851, 39.95248, 39.93626, 
    39.91983, 39.90319, 39.88635, 39.86931, 39.85207, 39.83462, 39.81697, 
    39.79911, 39.78106, 39.76281, 39.74435, 39.72569, 39.70683, 39.68777, 
    39.66851, 39.64905, 39.62939, 39.60953, 39.58947, 39.56921, 39.54874, 
    39.52809, 39.50723, 39.48618, 39.46492, 39.44347, 39.42182, 39.39997, 
    39.37793, 39.35569, 39.33325, 39.31062, 39.28779, 39.26476, 39.24154, 
    39.21813, 39.19452, 39.17071, 39.14671, 39.12252, 39.09813, 39.07355, 
    39.04877, 39.02381, 38.99865, 38.9733, 38.94775, 38.92202, 38.89609, 
    38.86997, 38.84366, 38.81716, 38.79047, 38.76359, 38.73652, 38.70926, 
    38.68181, 38.65417, 38.62635, 38.59834, 38.57013, 38.54174, 38.51317, 
    38.48441, 38.45546, 38.42632, 38.397, 38.36749, 38.3378, 38.30793, 
    38.27786, 38.24762, 38.21719, 38.18658, 38.15578, 38.1248, 38.09364, 
    38.0623, 38.03077, 37.99907, 37.96717, 37.93511, 37.90286, 37.87043, 
    37.83782, 37.80503, 37.77206, 37.73892, 37.70559, 37.67209, 37.63841, 
    37.60455, 37.57051,
  33.78909, 33.83799, 33.88676, 33.93538, 33.98385, 34.03219, 34.08038, 
    34.12843, 34.17633, 34.22409, 34.2717, 34.31917, 34.36649, 34.41367, 
    34.4607, 34.50759, 34.55432, 34.60091, 34.64735, 34.69365, 34.73979, 
    34.78579, 34.83163, 34.87732, 34.92287, 34.96826, 35.0135, 35.0586, 
    35.10354, 35.14832, 35.19296, 35.23744, 35.28177, 35.32594, 35.36996, 
    35.41383, 35.45754, 35.50109, 35.54449, 35.58773, 35.63082, 35.67375, 
    35.71652, 35.75914, 35.80159, 35.84389, 35.88603, 35.92801, 35.96983, 
    36.01149, 36.05299, 36.09433, 36.13551, 36.17652, 36.21738, 36.25807, 
    36.2986, 36.33896, 36.37917, 36.4192, 36.45908, 36.49879, 36.53833, 
    36.57771, 36.61692, 36.65597, 36.69485, 36.73357, 36.77211, 36.81049, 
    36.8487, 36.88674, 36.92462, 36.96232, 36.99986, 37.03722, 37.07441, 
    37.11144, 37.14829, 37.18497, 37.22148, 37.25782, 37.29398, 37.32998, 
    37.3658, 37.40144, 37.43691, 37.47221, 37.50733, 37.54228, 37.57705, 
    37.61164, 37.64606, 37.68031, 37.71437, 37.74826, 37.78197, 37.81551, 
    37.84886, 37.88204, 37.91504, 37.94785, 37.98049, 38.01295, 38.04523, 
    38.07733, 38.10924, 38.14098, 38.17253, 38.2039, 38.23509, 38.26609, 
    38.29692, 38.32756, 38.35801, 38.38828, 38.41837, 38.44827, 38.47799, 
    38.50751, 38.53686, 38.56602, 38.59499, 38.62378, 38.65237, 38.68079, 
    38.70901, 38.73705, 38.76489, 38.79255, 38.82002, 38.8473, 38.87439, 
    38.90129, 38.928, 38.95451, 38.98084, 39.00698, 39.03292, 39.05868, 
    39.08424, 39.10961, 39.13478, 39.15977, 39.18456, 39.20916, 39.23356, 
    39.25777, 39.28178, 39.3056, 39.32922, 39.35265, 39.37589, 39.39892, 
    39.42176, 39.44441, 39.46686, 39.48911, 39.51116, 39.53302, 39.55468, 
    39.57614, 39.5974, 39.61847, 39.63933, 39.66, 39.68046, 39.70073, 
    39.7208, 39.74067, 39.76033, 39.7798, 39.79906, 39.81813, 39.83699, 
    39.85566, 39.87412, 39.89238, 39.91043, 39.92829, 39.94594, 39.96339, 
    39.98063, 39.99768, 40.01451, 40.03115, 40.04758, 40.06381, 40.07983, 
    40.09565, 40.11127, 40.12667, 40.14188, 40.15688, 40.17167, 40.18626, 
    40.20064, 40.21482, 40.22879, 40.24255, 40.25611, 40.26945, 40.2826, 
    40.29553, 40.30826, 40.32079, 40.3331, 40.3452, 40.3571, 40.36879, 
    40.38027, 40.39155, 40.40261, 40.41347, 40.42411, 40.43456, 40.44479, 
    40.4548, 40.46461, 40.47422, 40.48361, 40.49279, 40.50177, 40.51053, 
    40.51908, 40.52742, 40.53556, 40.54348, 40.55119, 40.55869, 40.56598, 
    40.57306, 40.57993, 40.58659, 40.59304, 40.59927, 40.6053, 40.61111, 
    40.61671, 40.6221, 40.62728, 40.63225, 40.637, 40.64155, 40.64588, 40.65, 
    40.65391, 40.65761, 40.66109, 40.66437, 40.66743, 40.67028, 40.67291, 
    40.67534, 40.67755, 40.67955, 40.68134, 40.68291, 40.68428, 40.68543, 
    40.68637, 40.6871, 40.68761, 40.68791, 40.688, 40.68788, 40.68754, 
    40.68699, 40.68623, 40.68526, 40.68408, 40.68268, 40.68107, 40.67925, 
    40.67722, 40.67497, 40.67251, 40.66984, 40.66696, 40.66386, 40.66056, 
    40.65704, 40.65331, 40.64936, 40.64521, 40.64085, 40.63627, 40.63148, 
    40.62648, 40.62127, 40.61584, 40.6102, 40.60436, 40.5983, 40.59203, 
    40.58555, 40.57886, 40.57196, 40.56484, 40.55752, 40.54998, 40.54224, 
    40.53428, 40.52612, 40.51774, 40.50916, 40.50036, 40.49136, 40.48214, 
    40.47271, 40.46308, 40.45324, 40.44318, 40.43292, 40.42245, 40.41177, 
    40.40088, 40.38978, 40.37847, 40.36695, 40.35523, 40.3433, 40.33117, 
    40.31882, 40.30626, 40.2935, 40.28053, 40.26736, 40.25397, 40.24039, 
    40.22659, 40.21259, 40.19838, 40.18396, 40.16935, 40.15452, 40.13949, 
    40.12425, 40.10881, 40.09316, 40.07731, 40.06126, 40.045, 40.02853, 
    40.01187, 39.995, 39.97792, 39.96064, 39.94316, 39.92548, 39.90759, 
    39.8895, 39.87121, 39.85272, 39.83403, 39.81513, 39.79603, 39.77673, 
    39.75724, 39.73754, 39.71764, 39.69754, 39.67724, 39.65674, 39.63604, 
    39.61515, 39.59405, 39.57276, 39.55127, 39.52958, 39.50769, 39.4856, 
    39.46332, 39.44084, 39.41816, 39.39529, 39.37222, 39.34896, 39.3255, 
    39.30185, 39.27799, 39.25395, 39.22971, 39.20528, 39.18065, 39.15583, 
    39.13082, 39.10561, 39.08021, 39.05462, 39.02884, 39.00286, 38.97669, 
    38.95033, 38.92378, 38.89705, 38.87011, 38.84299, 38.81569, 38.78819, 
    38.7605, 38.73262, 38.70456, 38.6763, 38.64787, 38.61924, 38.59042, 
    38.56142, 38.53223, 38.50286, 38.4733, 38.44355, 38.41362, 38.3835, 
    38.35321, 38.32272, 38.29205, 38.2612, 38.23017, 38.19895, 38.16755, 
    38.13597, 38.10421, 38.07226, 38.04013, 38.00783, 37.97534, 37.94268, 
    37.90983, 37.8768, 37.8436, 37.81021, 37.77665, 37.74291, 37.709, 37.6749,
  33.88719, 33.93616, 33.985, 34.03369, 34.08224, 34.13065, 34.17891, 
    34.22703, 34.27501, 34.32284, 34.37053, 34.41807, 34.46546, 34.51271, 
    34.55981, 34.60677, 34.65358, 34.70024, 34.74675, 34.79311, 34.83933, 
    34.8854, 34.93131, 34.97708, 35.02269, 35.06816, 35.11347, 35.15863, 
    35.20364, 35.2485, 35.29321, 35.33776, 35.38216, 35.4264, 35.47049, 
    35.51442, 35.5582, 35.60183, 35.6453, 35.68861, 35.73177, 35.77477, 
    35.8176, 35.86029, 35.90281, 35.94518, 35.98738, 36.02943, 36.07132, 
    36.11305, 36.15462, 36.19602, 36.23727, 36.27835, 36.31927, 36.36003, 
    36.40063, 36.44106, 36.48133, 36.52143, 36.56137, 36.60115, 36.64076, 
    36.6802, 36.71948, 36.75859, 36.79754, 36.83632, 36.87493, 36.91338, 
    36.95165, 36.98976, 37.02769, 37.06546, 37.10306, 37.14049, 37.17775, 
    37.21483, 37.25175, 37.28849, 37.32507, 37.36147, 37.39769, 37.43375, 
    37.46963, 37.50533, 37.54087, 37.57623, 37.61141, 37.64642, 37.68125, 
    37.7159, 37.75039, 37.78469, 37.81881, 37.85276, 37.88653, 37.92012, 
    37.95354, 37.98677, 38.01983, 38.0527, 38.0854, 38.11792, 38.15025, 
    38.18241, 38.21438, 38.24617, 38.27778, 38.30921, 38.34045, 38.37151, 
    38.40239, 38.43308, 38.46359, 38.49392, 38.52406, 38.55401, 38.58378, 
    38.61337, 38.64277, 38.67198, 38.701, 38.72984, 38.75849, 38.78695, 
    38.81523, 38.84332, 38.87121, 38.89892, 38.92644, 38.95377, 38.98091, 
    39.00786, 39.03462, 39.06119, 39.08756, 39.11375, 39.13974, 39.16554, 
    39.19115, 39.21657, 39.24179, 39.26682, 39.29166, 39.3163, 39.34075, 
    39.365, 39.38906, 39.41292, 39.43659, 39.46006, 39.48334, 39.50642, 
    39.52931, 39.55199, 39.57449, 39.59678, 39.61887, 39.64077, 39.66247, 
    39.68398, 39.70528, 39.72638, 39.74729, 39.76799, 39.7885, 39.8088, 
    39.82891, 39.84882, 39.86852, 39.88802, 39.90733, 39.92643, 39.94533, 
    39.96403, 39.98252, 40.00082, 40.01891, 40.0368, 40.05448, 40.07196, 
    40.08924, 40.10632, 40.12319, 40.13986, 40.15632, 40.17258, 40.18864, 
    40.20449, 40.22013, 40.23557, 40.2508, 40.26583, 40.28065, 40.29527, 
    40.30968, 40.32388, 40.33788, 40.35167, 40.36525, 40.37863, 40.3918, 
    40.40476, 40.41751, 40.43006, 40.44239, 40.45452, 40.46645, 40.47816, 
    40.48966, 40.50096, 40.51205, 40.52292, 40.53359, 40.54405, 40.5543, 
    40.56434, 40.57417, 40.58379, 40.5932, 40.60241, 40.6114, 40.62017, 
    40.62875, 40.6371, 40.64525, 40.65319, 40.66092, 40.66843, 40.67574, 
    40.68283, 40.68972, 40.69639, 40.70285, 40.7091, 40.71513, 40.72096, 
    40.72657, 40.73197, 40.73716, 40.74214, 40.7469, 40.75146, 40.7558, 
    40.75993, 40.76384, 40.76755, 40.77104, 40.77432, 40.77739, 40.78024, 
    40.78288, 40.78531, 40.78753, 40.78954, 40.79132, 40.7929, 40.79427, 
    40.79543, 40.79636, 40.79709, 40.79761, 40.79791, 40.798, 40.79787, 
    40.79754, 40.79699, 40.79623, 40.79525, 40.79407, 40.79267, 40.79106, 
    40.78923, 40.78719, 40.78494, 40.78248, 40.7798, 40.77692, 40.77382, 
    40.7705, 40.76698, 40.76324, 40.75929, 40.75513, 40.75075, 40.74616, 
    40.74136, 40.73635, 40.73113, 40.7257, 40.72005, 40.71419, 40.70812, 
    40.70184, 40.69535, 40.68864, 40.68172, 40.6746, 40.66726, 40.65971, 
    40.65195, 40.64398, 40.6358, 40.6274, 40.6188, 40.60999, 40.60096, 
    40.59173, 40.58229, 40.57263, 40.56277, 40.5527, 40.54241, 40.53192, 
    40.52122, 40.51031, 40.49919, 40.48786, 40.47632, 40.46457, 40.45262, 
    40.44046, 40.42809, 40.41551, 40.40272, 40.38973, 40.37653, 40.36312, 
    40.3495, 40.33568, 40.32165, 40.30742, 40.29297, 40.27832, 40.26347, 
    40.24841, 40.23314, 40.21767, 40.20199, 40.18611, 40.17002, 40.15373, 
    40.13724, 40.12054, 40.10363, 40.08652, 40.06921, 40.0517, 40.03398, 
    40.01606, 39.99794, 39.97961, 39.96108, 39.94235, 39.92342, 39.90429, 
    39.88495, 39.86542, 39.84568, 39.82574, 39.80561, 39.78527, 39.76473, 
    39.74399, 39.72306, 39.70192, 39.68059, 39.65905, 39.63732, 39.61539, 
    39.59327, 39.57094, 39.54842, 39.5257, 39.50278, 39.47967, 39.45636, 
    39.43286, 39.40916, 39.38527, 39.36118, 39.33689, 39.31242, 39.28774, 
    39.26287, 39.23781, 39.21256, 39.18711, 39.16148, 39.13564, 39.10962, 
    39.0834, 39.057, 39.0304, 39.00361, 38.97663, 38.94946, 38.9221, 
    38.89455, 38.86681, 38.83889, 38.81077, 38.78246, 38.75397, 38.72529, 
    38.69642, 38.66737, 38.63813, 38.6087, 38.57909, 38.54929, 38.5193, 
    38.48913, 38.45878, 38.42824, 38.39752, 38.36661, 38.33552, 38.30425, 
    38.27279, 38.24115, 38.20934, 38.17733, 38.14515, 38.11279, 38.08024, 
    38.04752, 38.01461, 37.98153, 37.94827, 37.91482, 37.8812, 37.8474, 
    37.81343, 37.77927,
  33.98526, 34.03431, 34.08321, 34.13198, 34.1806, 34.22908, 34.27742, 
    34.32561, 34.37366, 34.42156, 34.46932, 34.51693, 34.5644, 34.61172, 
    34.6589, 34.70592, 34.7528, 34.79954, 34.84612, 34.89256, 34.93884, 
    34.98498, 35.03097, 35.07681, 35.12249, 35.16803, 35.21341, 35.25864, 
    35.30373, 35.34865, 35.39343, 35.43805, 35.48252, 35.52683, 35.57099, 
    35.615, 35.65885, 35.70254, 35.74608, 35.78946, 35.83268, 35.87575, 
    35.91866, 35.96141, 36.00401, 36.04644, 36.08872, 36.13084, 36.17279, 
    36.21459, 36.25622, 36.2977, 36.33901, 36.38016, 36.42115, 36.46198, 
    36.50264, 36.54314, 36.58347, 36.62364, 36.66365, 36.70349, 36.74317, 
    36.78268, 36.82202, 36.8612, 36.90021, 36.93906, 36.97773, 37.01624, 
    37.05458, 37.09275, 37.13075, 37.16858, 37.20625, 37.24374, 37.28106, 
    37.31821, 37.35519, 37.392, 37.42863, 37.4651, 37.50138, 37.5375, 
    37.57344, 37.60921, 37.64481, 37.68023, 37.71547, 37.75054, 37.78543, 
    37.82014, 37.85469, 37.88905, 37.92324, 37.95724, 37.99107, 38.02472, 
    38.0582, 38.09149, 38.12461, 38.15754, 38.19029, 38.22287, 38.25526, 
    38.28747, 38.3195, 38.35135, 38.38301, 38.4145, 38.4458, 38.47691, 
    38.50785, 38.5386, 38.56916, 38.59954, 38.62974, 38.65975, 38.68957, 
    38.71921, 38.74866, 38.77792, 38.807, 38.83589, 38.8646, 38.89311, 
    38.92144, 38.94957, 38.97752, 39.00528, 39.03285, 39.06023, 39.08742, 
    39.11442, 39.14123, 39.16785, 39.19427, 39.2205, 39.24655, 39.2724, 
    39.29805, 39.32352, 39.34879, 39.37386, 39.39875, 39.42344, 39.44793, 
    39.47223, 39.49633, 39.52024, 39.54395, 39.56747, 39.59079, 39.61391, 
    39.63684, 39.65957, 39.68211, 39.70444, 39.72658, 39.74852, 39.77026, 
    39.7918, 39.81314, 39.83429, 39.85524, 39.87598, 39.89653, 39.91687, 
    39.93702, 39.95696, 39.9767, 39.99624, 40.01558, 40.03472, 40.05366, 
    40.07239, 40.09092, 40.10925, 40.12738, 40.1453, 40.16302, 40.18054, 
    40.19785, 40.21496, 40.23186, 40.24857, 40.26506, 40.28135, 40.29744, 
    40.31332, 40.32899, 40.34446, 40.35972, 40.37478, 40.38963, 40.40428, 
    40.41871, 40.43295, 40.44697, 40.46078, 40.4744, 40.4878, 40.50099, 
    40.51398, 40.52676, 40.53933, 40.55169, 40.56384, 40.57579, 40.58752, 
    40.59905, 40.61037, 40.62148, 40.63238, 40.64307, 40.65355, 40.66382, 
    40.67388, 40.68373, 40.69337, 40.7028, 40.71202, 40.72102, 40.72982, 
    40.73841, 40.74678, 40.75495, 40.76291, 40.77065, 40.77818, 40.7855, 
    40.7926, 40.7995, 40.80619, 40.81266, 40.81892, 40.82497, 40.8308, 
    40.83643, 40.84184, 40.84704, 40.85203, 40.8568, 40.86136, 40.86572, 
    40.86985, 40.87378, 40.87749, 40.88099, 40.88427, 40.88734, 40.89021, 
    40.89285, 40.89529, 40.89751, 40.89952, 40.90131, 40.90289, 40.90426, 
    40.90542, 40.90636, 40.90709, 40.90761, 40.90791, 40.908, 40.90788, 
    40.90754, 40.90699, 40.90623, 40.90525, 40.90406, 40.90266, 40.90104, 
    40.89921, 40.89717, 40.89492, 40.89245, 40.88977, 40.88688, 40.88377, 
    40.88045, 40.87691, 40.87317, 40.86921, 40.86504, 40.86066, 40.85606, 
    40.85125, 40.84623, 40.841, 40.83555, 40.8299, 40.82402, 40.81794, 
    40.81165, 40.80514, 40.79842, 40.79149, 40.78435, 40.777, 40.76944, 
    40.76166, 40.75367, 40.74548, 40.73706, 40.72844, 40.71961, 40.71057, 
    40.70132, 40.69186, 40.68218, 40.6723, 40.66221, 40.65191, 40.64139, 
    40.63067, 40.61974, 40.60859, 40.59724, 40.58568, 40.57391, 40.56194, 
    40.54975, 40.53735, 40.52475, 40.51194, 40.49892, 40.48569, 40.47226, 
    40.45861, 40.44476, 40.43071, 40.41644, 40.40197, 40.38729, 40.37241, 
    40.35732, 40.34203, 40.32653, 40.31082, 40.29491, 40.27879, 40.26246, 
    40.24594, 40.2292, 40.21227, 40.19513, 40.17778, 40.16023, 40.14248, 
    40.12453, 40.10637, 40.08801, 40.06944, 40.05067, 40.03171, 40.01254, 
    39.99316, 39.97359, 39.95382, 39.93384, 39.91367, 39.89329, 39.87271, 
    39.85194, 39.83096, 39.80978, 39.78841, 39.76683, 39.74506, 39.72309, 
    39.70092, 39.67855, 39.65599, 39.63323, 39.61027, 39.58712, 39.56376, 
    39.54021, 39.51647, 39.49253, 39.4684, 39.44407, 39.41954, 39.39482, 
    39.36991, 39.3448, 39.3195, 39.29401, 39.26832, 39.24244, 39.21637, 
    39.19011, 39.16365, 39.137, 39.11016, 39.08313, 39.05592, 39.0285, 
    39.0009, 38.97311, 38.94514, 38.91697, 38.88861, 38.86007, 38.83134, 
    38.80241, 38.77331, 38.74401, 38.71453, 38.68486, 38.65501, 38.62497, 
    38.59475, 38.56434, 38.53374, 38.50297, 38.472, 38.44086, 38.40953, 
    38.37802, 38.34632, 38.31445, 38.28239, 38.25015, 38.21773, 38.18512, 
    38.15234, 38.11938, 38.08624, 38.05291, 38.01941, 37.98573, 37.95187, 
    37.91784, 37.88363,
  34.08329, 34.13242, 34.1814, 34.23024, 34.27893, 34.32748, 34.37589, 
    34.42416, 34.47228, 34.52026, 34.56809, 34.61577, 34.66331, 34.7107, 
    34.75795, 34.80505, 34.85201, 34.89881, 34.94546, 34.99197, 35.03833, 
    35.08454, 35.1306, 35.17651, 35.22226, 35.26787, 35.31332, 35.35863, 
    35.40378, 35.44878, 35.49363, 35.53832, 35.58286, 35.62724, 35.67147, 
    35.71555, 35.75946, 35.80323, 35.84684, 35.89029, 35.93358, 35.97672, 
    36.0197, 36.06252, 36.10518, 36.14768, 36.19003, 36.23221, 36.27424, 
    36.3161, 36.3578, 36.39935, 36.44073, 36.48195, 36.523, 36.56389, 
    36.60462, 36.64519, 36.68559, 36.72583, 36.7659, 36.80581, 36.84555, 
    36.88513, 36.92454, 36.96378, 37.00286, 37.04177, 37.08051, 37.11908, 
    37.15749, 37.19572, 37.23379, 37.27169, 37.30941, 37.34697, 37.38435, 
    37.42157, 37.45861, 37.49548, 37.53218, 37.5687, 37.60506, 37.64124, 
    37.67724, 37.71307, 37.74873, 37.78421, 37.81951, 37.85464, 37.8896, 
    37.92437, 37.95897, 37.9934, 38.02764, 38.06171, 38.0956, 38.12931, 
    38.16284, 38.19619, 38.22937, 38.26236, 38.29517, 38.3278, 38.36025, 
    38.39252, 38.42461, 38.45651, 38.48824, 38.51978, 38.55113, 38.58231, 
    38.61329, 38.6441, 38.67472, 38.70515, 38.7354, 38.76546, 38.79535, 
    38.82504, 38.85454, 38.88386, 38.91299, 38.94193, 38.97069, 38.99926, 
    39.02763, 39.05582, 39.08382, 39.11163, 39.13926, 39.16668, 39.19392, 
    39.22097, 39.24783, 39.2745, 39.30097, 39.32726, 39.35334, 39.37924, 
    39.40495, 39.43046, 39.45577, 39.4809, 39.50583, 39.53056, 39.5551, 
    39.57944, 39.6036, 39.62755, 39.65131, 39.67487, 39.69823, 39.7214, 
    39.74437, 39.76714, 39.78972, 39.8121, 39.83428, 39.85626, 39.87804, 
    39.89962, 39.92101, 39.94219, 39.96318, 39.98396, 40.00455, 40.02493, 
    40.04512, 40.0651, 40.08488, 40.10446, 40.12383, 40.14301, 40.16198, 
    40.18075, 40.19932, 40.21768, 40.23584, 40.2538, 40.27156, 40.28911, 
    40.30645, 40.3236, 40.34053, 40.35727, 40.37379, 40.39011, 40.40623, 
    40.42214, 40.43785, 40.45335, 40.46864, 40.48373, 40.49861, 40.51328, 
    40.52774, 40.542, 40.55606, 40.5699, 40.58354, 40.59697, 40.61019, 
    40.6232, 40.636, 40.6486, 40.66098, 40.67316, 40.68513, 40.69689, 
    40.70844, 40.71978, 40.73091, 40.74183, 40.75254, 40.76304, 40.77333, 
    40.78341, 40.79328, 40.80294, 40.81239, 40.82162, 40.83065, 40.83947, 
    40.84807, 40.85646, 40.86464, 40.87262, 40.88037, 40.88792, 40.89525, 
    40.90237, 40.90928, 40.91598, 40.92247, 40.92874, 40.9348, 40.94065, 
    40.94629, 40.95171, 40.95692, 40.96191, 40.9667, 40.97127, 40.97563, 
    40.97977, 40.98371, 40.98743, 40.99093, 40.99422, 40.9973, 41.00017, 
    41.00282, 41.00526, 41.00749, 41.0095, 41.0113, 41.01288, 41.01426, 
    41.01542, 41.01636, 41.01709, 41.0176, 41.01791, 41.018, 41.01788, 
    41.01754, 41.01699, 41.01622, 41.01524, 41.01405, 41.01265, 41.01103, 
    41.0092, 41.00715, 41.00489, 41.00242, 40.99973, 40.99683, 40.99372, 
    40.99039, 40.98685, 40.9831, 40.97913, 40.97495, 40.97056, 40.96596, 
    40.96114, 40.95611, 40.95086, 40.94541, 40.93974, 40.93386, 40.92776, 
    40.92146, 40.91494, 40.9082, 40.90126, 40.89411, 40.88674, 40.87916, 
    40.87137, 40.86337, 40.85515, 40.84673, 40.83809, 40.82924, 40.82018, 
    40.81091, 40.80143, 40.79174, 40.78183, 40.77172, 40.76139, 40.75086, 
    40.74012, 40.72916, 40.718, 40.70663, 40.69504, 40.68325, 40.67125, 
    40.65904, 40.64662, 40.63399, 40.62115, 40.60811, 40.59486, 40.58139, 
    40.56773, 40.55385, 40.53976, 40.52547, 40.51097, 40.49627, 40.48135, 
    40.46624, 40.45091, 40.43538, 40.41964, 40.40369, 40.38755, 40.37119, 
    40.35463, 40.33787, 40.3209, 40.30372, 40.28635, 40.26876, 40.25098, 
    40.23299, 40.21479, 40.1964, 40.1778, 40.15899, 40.13999, 40.12078, 
    40.10137, 40.08176, 40.06195, 40.04193, 40.02172, 40.0013, 39.98069, 
    39.95987, 39.93886, 39.91764, 39.89622, 39.87461, 39.85279, 39.83078, 
    39.80857, 39.78616, 39.76356, 39.74075, 39.71775, 39.69455, 39.67115, 
    39.64756, 39.62377, 39.59979, 39.57561, 39.55123, 39.52666, 39.5019, 
    39.47694, 39.45178, 39.42643, 39.40089, 39.37516, 39.34923, 39.32311, 
    39.2968, 39.27029, 39.2436, 39.21671, 39.18963, 39.16236, 39.1349, 
    39.10725, 39.07941, 39.05138, 39.02316, 38.99475, 38.96615, 38.93737, 
    38.90839, 38.87923, 38.84989, 38.82035, 38.79063, 38.76072, 38.73063, 
    38.70035, 38.66989, 38.63924, 38.6084, 38.57738, 38.54618, 38.5148, 
    38.48323, 38.45148, 38.41954, 38.38743, 38.35513, 38.32265, 38.28999, 
    38.25715, 38.22413, 38.19093, 38.15755, 38.12399, 38.09025, 38.05633, 
    38.02224, 37.98796,
  34.1813, 34.2305, 34.27955, 34.32846, 34.37724, 34.42586, 34.47434, 
    34.52268, 34.57087, 34.61892, 34.66682, 34.71458, 34.7622, 34.80966, 
    34.85698, 34.90415, 34.95118, 34.99805, 35.04478, 35.09136, 35.13779, 
    35.18407, 35.2302, 35.27618, 35.32201, 35.36769, 35.41321, 35.45859, 
    35.50381, 35.54888, 35.5938, 35.63856, 35.68317, 35.72762, 35.77192, 
    35.81607, 35.86006, 35.90389, 35.94757, 35.99109, 36.03445, 36.07766, 
    36.12071, 36.1636, 36.20633, 36.2489, 36.29131, 36.33357, 36.37566, 
    36.41759, 36.45936, 36.50097, 36.54242, 36.58371, 36.62483, 36.66579, 
    36.70659, 36.74722, 36.78769, 36.828, 36.86814, 36.90811, 36.94792, 
    36.98756, 37.02704, 37.06635, 37.10549, 37.14447, 37.18327, 37.22191, 
    37.26038, 37.29868, 37.33681, 37.37477, 37.41256, 37.45018, 37.48763, 
    37.52491, 37.56202, 37.59895, 37.63571, 37.67229, 37.70871, 37.74495, 
    37.78102, 37.81691, 37.85263, 37.88817, 37.92354, 37.95873, 37.99374, 
    38.02858, 38.06324, 38.09772, 38.13203, 38.16616, 38.20011, 38.23388, 
    38.26747, 38.30088, 38.33411, 38.36716, 38.40004, 38.43272, 38.46523, 
    38.49756, 38.5297, 38.56166, 38.59344, 38.62504, 38.65645, 38.68768, 
    38.71873, 38.74958, 38.78026, 38.81075, 38.84105, 38.87117, 38.9011, 
    38.93085, 38.96041, 38.98978, 39.01897, 39.04796, 39.07677, 39.10539, 
    39.13382, 39.16206, 39.19011, 39.21797, 39.24564, 39.27312, 39.30042, 
    39.32751, 39.35442, 39.38114, 39.40766, 39.43399, 39.46013, 39.48608, 
    39.51183, 39.53739, 39.56275, 39.58792, 39.6129, 39.63768, 39.66227, 
    39.68666, 39.71085, 39.73485, 39.75865, 39.78226, 39.80566, 39.82888, 
    39.85189, 39.87471, 39.89733, 39.91975, 39.94197, 39.96399, 39.98582, 
    40.00744, 40.02887, 40.05009, 40.07111, 40.09194, 40.11256, 40.13299, 
    40.15321, 40.17323, 40.19305, 40.21266, 40.23208, 40.25129, 40.2703, 
    40.2891, 40.30771, 40.32611, 40.34431, 40.3623, 40.38008, 40.39767, 
    40.41505, 40.43222, 40.4492, 40.46596, 40.48252, 40.49887, 40.51502, 
    40.53096, 40.5467, 40.56223, 40.57755, 40.59267, 40.60758, 40.62228, 
    40.63678, 40.65106, 40.66514, 40.67901, 40.69268, 40.70613, 40.71938, 
    40.73241, 40.74524, 40.75786, 40.77028, 40.78247, 40.79447, 40.80625, 
    40.81782, 40.82919, 40.84034, 40.85128, 40.86201, 40.87254, 40.88285, 
    40.89294, 40.90284, 40.91251, 40.92198, 40.93124, 40.94028, 40.94911, 
    40.95773, 40.96614, 40.97434, 40.98232, 40.9901, 40.99766, 41.00501, 
    41.01214, 41.01907, 41.02578, 41.03228, 41.03856, 41.04464, 41.0505, 
    41.05614, 41.06158, 41.0668, 41.0718, 41.0766, 41.08118, 41.08554, 
    41.0897, 41.09364, 41.09737, 41.10088, 41.10418, 41.10726, 41.11013, 
    41.11279, 41.11524, 41.11747, 41.11948, 41.12128, 41.12288, 41.12425, 
    41.12541, 41.12635, 41.12709, 41.12761, 41.12791, 41.128, 41.12788, 
    41.12754, 41.12698, 41.12622, 41.12524, 41.12405, 41.12263, 41.12101, 
    41.11918, 41.11713, 41.11486, 41.11238, 41.1097, 41.10679, 41.10367, 
    41.10034, 41.09679, 41.09303, 41.08905, 41.08487, 41.08047, 41.07585, 
    41.07103, 41.06598, 41.06073, 41.05526, 41.04958, 41.04369, 41.03758, 
    41.03126, 41.02473, 41.01799, 41.01103, 41.00386, 40.99648, 40.98888, 
    40.98108, 40.97306, 40.96482, 40.95638, 40.94773, 40.93886, 40.92978, 
    40.92049, 40.911, 40.90128, 40.89136, 40.88123, 40.87088, 40.86033, 
    40.84956, 40.83859, 40.8274, 40.81601, 40.8044, 40.79258, 40.78056, 
    40.76833, 40.75588, 40.74323, 40.73037, 40.7173, 40.70402, 40.69053, 
    40.67683, 40.66293, 40.64882, 40.63449, 40.61997, 40.60523, 40.59029, 
    40.57514, 40.55979, 40.54422, 40.52846, 40.51248, 40.4963, 40.47992, 
    40.46332, 40.44653, 40.42952, 40.41232, 40.39491, 40.37729, 40.35947, 
    40.34144, 40.32321, 40.30478, 40.28614, 40.26731, 40.24826, 40.22902, 
    40.20958, 40.18993, 40.17007, 40.15002, 40.12977, 40.10931, 40.08866, 
    40.0678, 40.04675, 40.02549, 40.00403, 39.98238, 39.96052, 39.93847, 
    39.91621, 39.89376, 39.87111, 39.84826, 39.82522, 39.80198, 39.77854, 
    39.7549, 39.73106, 39.70704, 39.68281, 39.65839, 39.63377, 39.60896, 
    39.58395, 39.55875, 39.53336, 39.50777, 39.48199, 39.45601, 39.42984, 
    39.40348, 39.37693, 39.35018, 39.32324, 39.29611, 39.26879, 39.24128, 
    39.21358, 39.18569, 39.1576, 39.12933, 39.10087, 39.07222, 39.04339, 
    39.01436, 38.98515, 38.95575, 38.92616, 38.89638, 38.86642, 38.83627, 
    38.80594, 38.77542, 38.74472, 38.71383, 38.68275, 38.6515, 38.62005, 
    38.58843, 38.55662, 38.52463, 38.49246, 38.4601, 38.42757, 38.39485, 
    38.36195, 38.32887, 38.29561, 38.26217, 38.22855, 38.19475, 38.16077, 
    38.12662, 38.09228,
  34.27929, 34.32855, 34.37768, 34.42667, 34.47551, 34.5242, 34.57276, 
    34.62117, 34.66944, 34.71756, 34.76553, 34.81337, 34.86105, 34.90859, 
    34.95598, 35.00322, 35.05032, 35.09727, 35.14407, 35.19072, 35.23722, 
    35.28357, 35.32977, 35.37582, 35.42173, 35.46748, 35.51307, 35.55852, 
    35.60381, 35.64895, 35.69394, 35.73877, 35.78345, 35.82798, 35.87235, 
    35.91656, 35.96062, 36.00453, 36.04827, 36.09187, 36.1353, 36.17857, 
    36.22169, 36.26465, 36.30745, 36.35009, 36.39257, 36.4349, 36.47706, 
    36.51906, 36.5609, 36.60258, 36.64409, 36.68545, 36.72664, 36.76767, 
    36.80853, 36.84923, 36.88977, 36.93014, 36.97035, 37.01039, 37.05026, 
    37.08997, 37.12951, 37.16889, 37.2081, 37.24714, 37.28601, 37.32471, 
    37.36325, 37.40162, 37.43981, 37.47784, 37.51569, 37.55338, 37.59089, 
    37.62823, 37.6654, 37.70239, 37.73922, 37.77587, 37.81235, 37.84865, 
    37.88478, 37.92073, 37.95651, 37.99212, 38.02755, 38.0628, 38.09787, 
    38.13277, 38.1675, 38.20204, 38.2364, 38.27059, 38.3046, 38.33843, 
    38.37208, 38.40555, 38.43884, 38.47195, 38.50488, 38.53763, 38.57019, 
    38.60258, 38.63478, 38.6668, 38.69864, 38.73029, 38.76176, 38.79304, 
    38.82414, 38.85506, 38.88579, 38.91634, 38.94669, 38.97687, 39.00686, 
    39.03665, 39.06627, 39.09569, 39.12493, 39.15398, 39.18284, 39.21151, 
    39.23999, 39.26828, 39.29639, 39.3243, 39.35202, 39.37955, 39.40689, 
    39.43404, 39.461, 39.48777, 39.51434, 39.54072, 39.56691, 39.5929, 
    39.6187, 39.64431, 39.66972, 39.69494, 39.71996, 39.74479, 39.76942, 
    39.79386, 39.8181, 39.84214, 39.86599, 39.88964, 39.91309, 39.93635, 
    39.9594, 39.98227, 40.00492, 40.02739, 40.04965, 40.07172, 40.09358, 
    40.11525, 40.13671, 40.15798, 40.17905, 40.19991, 40.22057, 40.24104, 
    40.2613, 40.28135, 40.30121, 40.32087, 40.34032, 40.35957, 40.37861, 
    40.39745, 40.4161, 40.43453, 40.45276, 40.47079, 40.48861, 40.50623, 
    40.52364, 40.54085, 40.55785, 40.57465, 40.59124, 40.60763, 40.62381, 
    40.63978, 40.65555, 40.67111, 40.68646, 40.70161, 40.71655, 40.73128, 
    40.7458, 40.76012, 40.77422, 40.78812, 40.80181, 40.81529, 40.82856, 
    40.84163, 40.85448, 40.86713, 40.87956, 40.89179, 40.9038, 40.91561, 
    40.9272, 40.93859, 40.94976, 40.96073, 40.97148, 40.98203, 40.99236, 
    41.00248, 41.01239, 41.02208, 41.03157, 41.04084, 41.0499, 41.05875, 
    41.06739, 41.07582, 41.08403, 41.09203, 41.09982, 41.1074, 41.11476, 
    41.12191, 41.12885, 41.13557, 41.14209, 41.14838, 41.15447, 41.16034, 
    41.166, 41.17144, 41.17667, 41.18169, 41.18649, 41.19108, 41.19546, 
    41.19962, 41.20357, 41.2073, 41.21082, 41.21413, 41.21722, 41.2201, 
    41.22276, 41.22521, 41.22745, 41.22947, 41.23127, 41.23286, 41.23424, 
    41.2354, 41.23635, 41.23708, 41.23761, 41.23791, 41.238, 41.23788, 
    41.23754, 41.23698, 41.23622, 41.23523, 41.23404, 41.23262, 41.231, 
    41.22916, 41.22711, 41.22484, 41.22235, 41.21966, 41.21675, 41.21362, 
    41.21028, 41.20673, 41.20296, 41.19898, 41.19478, 41.19037, 41.18575, 
    41.18091, 41.17586, 41.17059, 41.16512, 41.15942, 41.15352, 41.1474, 
    41.14107, 41.13453, 41.12777, 41.1208, 41.11361, 41.10621, 41.0986, 
    41.09078, 41.08275, 41.0745, 41.06604, 41.05737, 41.04848, 41.03939, 
    41.03008, 41.02056, 41.01083, 41.00089, 40.99073, 40.98037, 40.9698, 
    40.95901, 40.94801, 40.9368, 40.92538, 40.91376, 40.90192, 40.88987, 
    40.87761, 40.86514, 40.85246, 40.83958, 40.82648, 40.81318, 40.79966, 
    40.78594, 40.772, 40.75787, 40.74352, 40.72896, 40.7142, 40.69923, 
    40.68405, 40.66866, 40.65307, 40.63727, 40.62127, 40.60505, 40.58863, 
    40.57201, 40.55518, 40.53814, 40.5209, 40.50346, 40.48581, 40.46795, 
    40.44989, 40.43163, 40.41316, 40.39449, 40.37561, 40.35653, 40.33725, 
    40.31777, 40.29808, 40.27819, 40.2581, 40.23781, 40.21732, 40.19662, 
    40.17573, 40.15463, 40.13333, 40.11184, 40.09014, 40.06824, 40.04614, 
    40.02385, 40.00135, 39.97866, 39.95577, 39.93268, 39.90939, 39.88591, 
    39.86223, 39.83835, 39.81427, 39.79, 39.76554, 39.74088, 39.71601, 
    39.69096, 39.66571, 39.64027, 39.61464, 39.5888, 39.56278, 39.53656, 
    39.51015, 39.48355, 39.45675, 39.42976, 39.40258, 39.37521, 39.34765, 
    39.3199, 39.29195, 39.26382, 39.2355, 39.20699, 39.17828, 39.14939, 
    39.12032, 39.09105, 39.0616, 39.03195, 39.00212, 38.97211, 38.94191, 
    38.91151, 38.88094, 38.85018, 38.81924, 38.78811, 38.75679, 38.7253, 
    38.69361, 38.66175, 38.6297, 38.59747, 38.56506, 38.53246, 38.49968, 
    38.46673, 38.43359, 38.40027, 38.36677, 38.33309, 38.29923, 38.2652, 
    38.23098, 38.19659,
  34.37724, 34.42658, 34.47578, 34.52483, 34.57375, 34.62252, 34.67115, 
    34.71964, 34.76797, 34.81617, 34.86422, 34.91212, 34.95988, 35.00749, 
    35.05495, 35.10227, 35.14944, 35.19646, 35.24333, 35.29005, 35.33662, 
    35.38305, 35.42932, 35.47544, 35.52142, 35.56724, 35.61291, 35.65842, 
    35.70379, 35.749, 35.79406, 35.83896, 35.88371, 35.92831, 35.97275, 
    36.01704, 36.06116, 36.10514, 36.14896, 36.19262, 36.23612, 36.27946, 
    36.32265, 36.36568, 36.40855, 36.45126, 36.49381, 36.53621, 36.57843, 
    36.6205, 36.66241, 36.70416, 36.74574, 36.78717, 36.82842, 36.86952, 
    36.91045, 36.95122, 36.99183, 37.03226, 37.07254, 37.11264, 37.15258, 
    37.19236, 37.23197, 37.27141, 37.31068, 37.34979, 37.38873, 37.4275, 
    37.4661, 37.50453, 37.54279, 37.58088, 37.6188, 37.65655, 37.69412, 
    37.73153, 37.76876, 37.80582, 37.84271, 37.87943, 37.91597, 37.95233, 
    37.98852, 38.02454, 38.06038, 38.09605, 38.13154, 38.16685, 38.20199, 
    38.23695, 38.27173, 38.30634, 38.34076, 38.37501, 38.40908, 38.44297, 
    38.47668, 38.51021, 38.54356, 38.57673, 38.60971, 38.64252, 38.67514, 
    38.70758, 38.73985, 38.77192, 38.80381, 38.83553, 38.86705, 38.89839, 
    38.92955, 38.96052, 38.99131, 39.0219, 39.05232, 39.08255, 39.11259, 
    39.14244, 39.17211, 39.20159, 39.23088, 39.25998, 39.28889, 39.31762, 
    39.34615, 39.3745, 39.40265, 39.43062, 39.45839, 39.48597, 39.51337, 
    39.54057, 39.56757, 39.59439, 39.62101, 39.64744, 39.67368, 39.69972, 
    39.72557, 39.75122, 39.77668, 39.80194, 39.82701, 39.85189, 39.87656, 
    39.90105, 39.92533, 39.94942, 39.97332, 39.99701, 40.02051, 40.04381, 
    40.06691, 40.08981, 40.11252, 40.13502, 40.15733, 40.17944, 40.20134, 
    40.22305, 40.24456, 40.26586, 40.28697, 40.30787, 40.32858, 40.34908, 
    40.36938, 40.38947, 40.40937, 40.42906, 40.44855, 40.46783, 40.48692, 
    40.5058, 40.52448, 40.54295, 40.56121, 40.57927, 40.59713, 40.61478, 
    40.63223, 40.64948, 40.66651, 40.68334, 40.69997, 40.71638, 40.73259, 
    40.7486, 40.7644, 40.77999, 40.79537, 40.81054, 40.82551, 40.84027, 
    40.85482, 40.86917, 40.8833, 40.89723, 40.91094, 40.92445, 40.93775, 
    40.95084, 40.96372, 40.97639, 40.98885, 41.0011, 41.01314, 41.02497, 
    41.03659, 41.04799, 41.05919, 41.07018, 41.08095, 41.09151, 41.10186, 
    41.11201, 41.12193, 41.13165, 41.14116, 41.15045, 41.15953, 41.1684, 
    41.17705, 41.18549, 41.19372, 41.20174, 41.20955, 41.21714, 41.22451, 
    41.23168, 41.23863, 41.24537, 41.25189, 41.2582, 41.2643, 41.27018, 
    41.27585, 41.28131, 41.28655, 41.29158, 41.29639, 41.30099, 41.30537, 
    41.30954, 41.3135, 41.31724, 41.32077, 41.32408, 41.32718, 41.33006, 
    41.33273, 41.33519, 41.33743, 41.33945, 41.34126, 41.34285, 41.34423, 
    41.3454, 41.34635, 41.34708, 41.3476, 41.34791, 41.348, 41.34787, 
    41.34753, 41.34698, 41.34621, 41.34523, 41.34403, 41.34262, 41.34099, 
    41.33914, 41.33709, 41.33481, 41.33232, 41.32962, 41.3267, 41.32357, 
    41.32022, 41.31667, 41.31289, 41.3089, 41.3047, 41.30028, 41.29564, 
    41.2908, 41.28574, 41.28046, 41.27497, 41.26927, 41.26335, 41.25722, 
    41.25087, 41.24432, 41.23755, 41.23056, 41.22336, 41.21595, 41.20832, 
    41.20049, 41.19244, 41.18417, 41.1757, 41.16701, 41.1581, 41.14899, 
    41.13967, 41.13013, 41.12038, 41.11042, 41.10024, 41.08986, 41.07926, 
    41.06845, 41.05743, 41.0462, 41.03476, 41.02311, 41.01125, 40.99918, 
    40.98689, 40.9744, 40.9617, 40.94878, 40.93566, 40.92233, 40.90879, 
    40.89504, 40.88108, 40.86691, 40.85254, 40.83795, 40.82316, 40.80816, 
    40.79295, 40.77753, 40.76191, 40.74608, 40.73004, 40.7138, 40.69735, 
    40.68069, 40.66383, 40.64676, 40.62949, 40.61201, 40.59432, 40.57643, 
    40.55833, 40.54004, 40.52153, 40.50283, 40.48391, 40.4648, 40.44548, 
    40.42596, 40.40623, 40.38631, 40.36618, 40.34585, 40.32531, 40.30458, 
    40.28364, 40.2625, 40.24117, 40.21963, 40.19789, 40.17595, 40.15381, 
    40.13148, 40.10894, 40.0862, 40.06327, 40.04013, 40.0168, 39.99327, 
    39.96955, 39.94563, 39.9215, 39.89719, 39.87267, 39.84797, 39.82306, 
    39.79796, 39.77266, 39.74717, 39.72149, 39.69561, 39.66954, 39.64327, 
    39.61681, 39.59016, 39.56331, 39.53627, 39.50904, 39.48162, 39.45401, 
    39.42621, 39.39821, 39.37003, 39.34165, 39.31309, 39.28433, 39.25539, 
    39.22626, 39.19694, 39.16743, 39.13773, 39.10785, 39.07778, 39.04752, 
    39.01708, 38.98645, 38.95563, 38.92463, 38.89344, 38.86208, 38.83052, 
    38.79878, 38.76686, 38.73475, 38.70247, 38.66999, 38.63734, 38.60451, 
    38.57149, 38.5383, 38.50492, 38.47136, 38.43762, 38.4037, 38.36961, 
    38.33533, 38.30087,
  34.47515, 34.52457, 34.57384, 34.62297, 34.67197, 34.72081, 34.76951, 
    34.81807, 34.86648, 34.91475, 34.96287, 35.01085, 35.05867, 35.10636, 
    35.1539, 35.20128, 35.24852, 35.29562, 35.34256, 35.38935, 35.436, 
    35.4825, 35.52884, 35.57504, 35.62108, 35.66697, 35.71272, 35.7583, 
    35.80374, 35.84902, 35.89415, 35.93913, 35.98395, 36.02861, 36.07313, 
    36.11749, 36.16168, 36.20573, 36.24961, 36.29335, 36.33692, 36.38033, 
    36.42359, 36.46669, 36.50963, 36.55241, 36.59503, 36.63749, 36.67979, 
    36.72192, 36.7639, 36.80572, 36.84737, 36.88886, 36.93019, 36.97135, 
    37.01235, 37.05318, 37.09386, 37.13436, 37.1747, 37.21488, 37.25489, 
    37.29473, 37.3344, 37.37391, 37.41325, 37.45242, 37.49143, 37.53026, 
    37.56893, 37.60742, 37.64575, 37.6839, 37.72189, 37.7597, 37.79734, 
    37.83481, 37.87211, 37.90923, 37.94618, 37.98296, 38.01957, 38.05599, 
    38.09225, 38.12833, 38.16423, 38.19996, 38.23551, 38.27089, 38.30608, 
    38.34111, 38.37595, 38.41061, 38.4451, 38.47941, 38.51354, 38.54749, 
    38.58126, 38.61485, 38.64826, 38.68148, 38.71453, 38.74739, 38.78008, 
    38.81258, 38.84489, 38.87703, 38.90898, 38.94075, 38.97233, 39.00373, 
    39.03494, 39.06596, 39.09681, 39.12746, 39.15793, 39.18821, 39.21831, 
    39.24822, 39.27794, 39.30747, 39.33682, 39.36597, 39.39494, 39.42372, 
    39.4523, 39.4807, 39.50891, 39.53692, 39.56475, 39.59238, 39.61982, 
    39.64707, 39.67413, 39.701, 39.72767, 39.75415, 39.78043, 39.80652, 
    39.83242, 39.85812, 39.88363, 39.90894, 39.93406, 39.95898, 39.9837, 
    40.00823, 40.03256, 40.0567, 40.08064, 40.10437, 40.12791, 40.15126, 
    40.1744, 40.19735, 40.2201, 40.24265, 40.265, 40.28715, 40.30909, 
    40.33084, 40.35239, 40.37374, 40.39489, 40.41583, 40.43657, 40.45711, 
    40.47745, 40.49759, 40.51752, 40.53725, 40.55678, 40.5761, 40.59522, 
    40.61414, 40.63285, 40.65136, 40.66966, 40.68776, 40.70565, 40.72334, 
    40.74081, 40.75809, 40.77516, 40.79202, 40.80868, 40.82513, 40.84137, 
    40.85741, 40.87324, 40.88886, 40.90427, 40.91948, 40.93447, 40.94926, 
    40.96384, 40.97821, 40.99237, 41.00633, 41.02007, 41.03361, 41.04693, 
    41.06005, 41.07295, 41.08565, 41.09813, 41.1104, 41.12247, 41.13432, 
    41.14597, 41.15739, 41.16861, 41.17962, 41.19042, 41.201, 41.21137, 
    41.22153, 41.23148, 41.24122, 41.25074, 41.26005, 41.26915, 41.27803, 
    41.28671, 41.29517, 41.30341, 41.31145, 41.31927, 41.32687, 41.33427, 
    41.34145, 41.34841, 41.35516, 41.3617, 41.36802, 41.37413, 41.38003, 
    41.38571, 41.39117, 41.39643, 41.40146, 41.40629, 41.4109, 41.41529, 
    41.41947, 41.42343, 41.42718, 41.43071, 41.43403, 41.43714, 41.44003, 
    41.4427, 41.44516, 41.4474, 41.44943, 41.45124, 41.45284, 41.45422, 
    41.45539, 41.45634, 41.45708, 41.4576, 41.45791, 41.458, 41.45787, 
    41.45753, 41.45698, 41.45621, 41.45522, 41.45402, 41.45261, 41.45097, 
    41.44912, 41.44706, 41.44479, 41.44229, 41.43958, 41.43666, 41.43352, 
    41.43017, 41.4266, 41.42282, 41.41882, 41.41461, 41.41018, 41.40554, 
    41.40068, 41.39561, 41.39032, 41.38482, 41.37911, 41.37318, 41.36704, 
    41.36068, 41.35411, 41.34732, 41.34032, 41.33311, 41.32568, 41.31805, 
    41.31019, 41.30212, 41.29384, 41.28535, 41.27665, 41.26773, 41.25859, 
    41.24925, 41.23969, 41.22992, 41.21994, 41.20975, 41.19934, 41.18872, 
    41.17789, 41.16685, 41.1556, 41.14413, 41.13246, 41.12057, 41.10848, 
    41.09617, 41.08365, 41.07093, 41.05799, 41.04484, 41.03148, 41.01791, 
    41.00414, 40.99015, 40.97596, 40.96155, 40.94694, 40.93211, 40.91708, 
    40.90185, 40.8864, 40.87075, 40.85489, 40.83882, 40.82254, 40.80606, 
    40.78937, 40.77247, 40.75537, 40.73806, 40.72055, 40.70283, 40.68491, 
    40.66677, 40.64844, 40.6299, 40.61116, 40.59221, 40.57306, 40.5537, 
    40.53414, 40.51438, 40.49442, 40.47425, 40.45388, 40.4333, 40.41253, 
    40.39155, 40.37038, 40.349, 40.32742, 40.30564, 40.28366, 40.26147, 
    40.23909, 40.21651, 40.19374, 40.17076, 40.14758, 40.12421, 40.10063, 
    40.07686, 40.05289, 40.02872, 40.00436, 39.9798, 39.95505, 39.9301, 
    39.90495, 39.8796, 39.85407, 39.82833, 39.80241, 39.77629, 39.74997, 
    39.72346, 39.69676, 39.66986, 39.64278, 39.61549, 39.58802, 39.56036, 
    39.53251, 39.50446, 39.47622, 39.44779, 39.41918, 39.39037, 39.36137, 
    39.33219, 39.30281, 39.27325, 39.2435, 39.21356, 39.18344, 39.15313, 
    39.12263, 39.09194, 39.06107, 39.03001, 38.99877, 38.96734, 38.93573, 
    38.90394, 38.87196, 38.83979, 38.80745, 38.77492, 38.74221, 38.70932, 
    38.67624, 38.64298, 38.60955, 38.57593, 38.54213, 38.50815, 38.474, 
    38.43966, 38.40514,
  34.57304, 34.62254, 34.67188, 34.72109, 34.77015, 34.81907, 34.86784, 
    34.91647, 34.96496, 35.0133, 35.06149, 35.10954, 35.15744, 35.2052, 
    35.25281, 35.30027, 35.34758, 35.39475, 35.44176, 35.48863, 35.53535, 
    35.58192, 35.62834, 35.6746, 35.72072, 35.76669, 35.8125, 35.85816, 
    35.90366, 35.94902, 35.99422, 36.03926, 36.08416, 36.12889, 36.17348, 
    36.2179, 36.26218, 36.30629, 36.35025, 36.39405, 36.43769, 36.48117, 
    36.5245, 36.56767, 36.61068, 36.65353, 36.69622, 36.73875, 36.78112, 
    36.82332, 36.86537, 36.90725, 36.94897, 36.99053, 37.03193, 37.07316, 
    37.11422, 37.15513, 37.19587, 37.23644, 37.27685, 37.31709, 37.35717, 
    37.39708, 37.43682, 37.47639, 37.5158, 37.55503, 37.5941, 37.633, 
    37.67173, 37.7103, 37.74869, 37.78691, 37.82495, 37.86283, 37.90054, 
    37.93807, 37.97543, 38.01262, 38.04964, 38.08648, 38.12315, 38.15964, 
    38.19595, 38.2321, 38.26806, 38.30385, 38.33947, 38.3749, 38.41016, 
    38.44525, 38.48015, 38.51488, 38.54943, 38.58379, 38.61798, 38.65199, 
    38.68582, 38.71947, 38.75294, 38.78622, 38.81933, 38.85225, 38.88499, 
    38.91755, 38.94993, 38.98212, 39.01413, 39.04595, 39.07759, 39.10904, 
    39.14031, 39.1714, 39.20229, 39.23301, 39.26353, 39.29387, 39.32402, 
    39.35398, 39.38376, 39.41335, 39.44274, 39.47195, 39.50097, 39.5298, 
    39.55844, 39.58689, 39.61515, 39.64322, 39.67109, 39.69878, 39.72627, 
    39.75357, 39.78068, 39.80759, 39.83432, 39.86084, 39.88718, 39.91331, 
    39.93926, 39.96501, 39.99057, 40.01593, 40.04109, 40.06606, 40.09083, 
    40.11541, 40.13978, 40.16396, 40.18795, 40.21173, 40.23532, 40.25871, 
    40.28189, 40.30489, 40.32767, 40.35027, 40.37266, 40.39485, 40.41684, 
    40.43863, 40.46022, 40.48161, 40.5028, 40.52378, 40.54456, 40.56514, 
    40.58552, 40.60569, 40.62567, 40.64544, 40.665, 40.68436, 40.70352, 
    40.72247, 40.74122, 40.75976, 40.7781, 40.79623, 40.81416, 40.83188, 
    40.8494, 40.8667, 40.88381, 40.9007, 40.91739, 40.93387, 40.95015, 
    40.96622, 40.98207, 40.99773, 41.01317, 41.0284, 41.04343, 41.05825, 
    41.07286, 41.08726, 41.10145, 41.11543, 41.1292, 41.14276, 41.15611, 
    41.16925, 41.18219, 41.1949, 41.20741, 41.21971, 41.2318, 41.24368, 
    41.25534, 41.26679, 41.27803, 41.28906, 41.29988, 41.31049, 41.32088, 
    41.33106, 41.34103, 41.35078, 41.36032, 41.36966, 41.37877, 41.38768, 
    41.39637, 41.40484, 41.41311, 41.42115, 41.42899, 41.43661, 41.44402, 
    41.45121, 41.45819, 41.46495, 41.47151, 41.47784, 41.48396, 41.48987, 
    41.49556, 41.50104, 41.5063, 41.51135, 41.51618, 41.5208, 41.5252, 
    41.52939, 41.53336, 41.53712, 41.54066, 41.54399, 41.5471, 41.54999, 
    41.55267, 41.55513, 41.55738, 41.55941, 41.56123, 41.56283, 41.56422, 
    41.56539, 41.56634, 41.56708, 41.5676, 41.56791, 41.568, 41.56787, 
    41.56754, 41.56698, 41.5662, 41.56522, 41.56401, 41.56259, 41.56096, 
    41.55911, 41.55704, 41.55476, 41.55226, 41.54955, 41.54662, 41.54347, 
    41.54012, 41.53654, 41.53275, 41.52874, 41.52452, 41.52008, 41.51543, 
    41.51057, 41.50549, 41.50019, 41.49468, 41.48895, 41.48301, 41.47685, 
    41.47049, 41.4639, 41.4571, 41.45009, 41.44286, 41.43542, 41.42776, 
    41.4199, 41.41181, 41.40351, 41.395, 41.38628, 41.37734, 41.36819, 
    41.35883, 41.34925, 41.33947, 41.32946, 41.31925, 41.30882, 41.29818, 
    41.28733, 41.27627, 41.265, 41.25351, 41.24181, 41.2299, 41.21778, 
    41.20545, 41.19291, 41.18015, 41.16719, 41.15401, 41.14063, 41.12704, 
    41.11323, 41.09922, 41.085, 41.07056, 41.05592, 41.04107, 41.02601, 
    41.01074, 40.99527, 40.97958, 40.96369, 40.94759, 40.93128, 40.91476, 
    40.89804, 40.88111, 40.86398, 40.84664, 40.82909, 40.81134, 40.79338, 
    40.77521, 40.75684, 40.73827, 40.71949, 40.7005, 40.68131, 40.66192, 
    40.64232, 40.62252, 40.60252, 40.58231, 40.5619, 40.54129, 40.52047, 
    40.49946, 40.47824, 40.45682, 40.4352, 40.41338, 40.39135, 40.36913, 
    40.34671, 40.32409, 40.30126, 40.27824, 40.25502, 40.2316, 40.20798, 
    40.18417, 40.16015, 40.13594, 40.11153, 40.08693, 40.06212, 40.03712, 
    40.01193, 39.98654, 39.96095, 39.93517, 39.90919, 39.88302, 39.85666, 
    39.8301, 39.80335, 39.77641, 39.74926, 39.72194, 39.69441, 39.66669, 
    39.63879, 39.61069, 39.5824, 39.55392, 39.52525, 39.49639, 39.46734, 
    39.43811, 39.40868, 39.37906, 39.34925, 39.31926, 39.28908, 39.25872, 
    39.22816, 39.19742, 39.16649, 39.13538, 39.10408, 39.0726, 39.04093, 
    39.00908, 38.97704, 38.94482, 38.91241, 38.87983, 38.84706, 38.81411, 
    38.78097, 38.74766, 38.71416, 38.68048, 38.64663, 38.61259, 38.57837, 
    38.54397, 38.5094,
  34.67091, 34.72047, 34.76989, 34.81917, 34.86831, 34.9173, 34.96614, 
    35.01485, 35.0634, 35.11182, 35.16009, 35.20821, 35.25618, 35.30401, 
    35.3517, 35.39923, 35.44662, 35.49385, 35.54094, 35.58788, 35.63467, 
    35.68131, 35.7278, 35.77414, 35.82033, 35.86637, 35.91225, 35.95798, 
    36.00356, 36.04898, 36.09426, 36.13938, 36.18434, 36.22915, 36.2738, 
    36.3183, 36.36264, 36.40683, 36.45086, 36.49472, 36.53844, 36.58199, 
    36.62539, 36.66863, 36.71171, 36.75463, 36.79739, 36.83998, 36.88242, 
    36.9247, 36.96681, 37.00876, 37.05055, 37.09218, 37.13364, 37.17494, 
    37.21608, 37.25705, 37.29786, 37.3385, 37.37897, 37.41928, 37.45942, 
    37.4994, 37.53921, 37.57885, 37.61832, 37.65763, 37.69676, 37.73573, 
    37.77452, 37.81315, 37.8516, 37.88989, 37.92801, 37.96595, 38.00372, 
    38.04132, 38.07874, 38.11599, 38.15307, 38.18998, 38.22671, 38.26326, 
    38.29964, 38.33585, 38.37188, 38.40773, 38.44341, 38.4789, 38.51423, 
    38.54937, 38.58434, 38.61913, 38.65373, 38.68816, 38.72241, 38.75648, 
    38.79037, 38.82408, 38.8576, 38.89095, 38.92412, 38.9571, 38.9899, 
    39.02251, 39.05495, 39.0872, 39.11926, 39.15114, 39.18284, 39.21435, 
    39.24567, 39.27682, 39.30777, 39.33854, 39.36912, 39.39951, 39.42971, 
    39.45973, 39.48956, 39.5192, 39.54866, 39.57792, 39.60699, 39.63587, 
    39.66457, 39.69307, 39.72138, 39.7495, 39.77743, 39.80516, 39.83271, 
    39.86006, 39.88721, 39.91418, 39.94095, 39.96753, 39.99391, 40.0201, 
    40.0461, 40.07189, 40.0975, 40.12291, 40.14812, 40.17313, 40.19795, 
    40.22257, 40.24699, 40.27122, 40.29525, 40.31908, 40.34271, 40.36614, 
    40.38937, 40.41241, 40.43524, 40.45788, 40.48031, 40.50254, 40.52458, 
    40.54641, 40.56804, 40.58947, 40.6107, 40.63172, 40.65255, 40.67316, 
    40.69358, 40.71379, 40.73381, 40.75361, 40.77322, 40.79261, 40.81181, 
    40.8308, 40.84958, 40.86816, 40.88653, 40.9047, 40.92266, 40.94042, 
    40.95797, 40.97531, 40.99245, 41.00938, 41.0261, 41.04261, 41.05892, 
    41.07502, 41.09091, 41.10659, 41.12207, 41.13733, 41.15239, 41.16723, 
    41.18187, 41.1963, 41.21052, 41.22453, 41.23832, 41.25191, 41.26529, 
    41.27846, 41.29141, 41.30416, 41.31669, 41.32901, 41.34113, 41.35303, 
    41.36472, 41.37619, 41.38745, 41.39851, 41.40934, 41.41997, 41.43039, 
    41.44059, 41.45057, 41.46035, 41.46991, 41.47926, 41.48839, 41.49731, 
    41.50602, 41.51451, 41.52279, 41.53086, 41.53871, 41.54634, 41.55377, 
    41.56098, 41.56797, 41.57475, 41.58131, 41.58766, 41.5938, 41.59971, 
    41.60542, 41.6109, 41.61618, 41.62123, 41.62608, 41.63071, 41.63512, 
    41.63931, 41.64329, 41.64706, 41.6506, 41.65394, 41.65705, 41.65995, 
    41.66264, 41.66511, 41.66736, 41.6694, 41.67122, 41.67282, 41.67421, 
    41.67538, 41.67634, 41.67708, 41.6776, 41.67791, 41.678, 41.67788, 
    41.67753, 41.67698, 41.6762, 41.67521, 41.674, 41.67258, 41.67094, 
    41.66909, 41.66702, 41.66473, 41.66223, 41.65951, 41.65657, 41.65342, 
    41.65006, 41.64648, 41.64268, 41.63866, 41.63443, 41.62999, 41.62533, 
    41.62045, 41.61536, 41.61005, 41.60453, 41.59879, 41.59284, 41.58667, 
    41.58029, 41.57369, 41.56688, 41.55985, 41.55261, 41.54515, 41.53748, 
    41.5296, 41.5215, 41.51318, 41.50466, 41.49591, 41.48696, 41.47779, 
    41.46841, 41.45882, 41.44901, 41.43898, 41.42875, 41.4183, 41.40764, 
    41.39677, 41.38568, 41.37439, 41.36288, 41.35116, 41.33923, 41.32708, 
    41.31472, 41.30215, 41.28938, 41.27639, 41.26319, 41.24978, 41.23616, 
    41.22232, 41.20828, 41.19403, 41.17957, 41.1649, 41.15002, 41.13493, 
    41.11963, 41.10413, 41.08841, 41.07249, 41.05635, 41.04002, 41.02347, 
    41.00671, 40.98975, 40.97258, 40.95521, 40.93763, 40.91983, 40.90184, 
    40.88364, 40.86523, 40.84662, 40.8278, 40.80878, 40.78956, 40.77013, 
    40.75049, 40.73066, 40.71061, 40.69036, 40.66992, 40.64927, 40.62841, 
    40.60735, 40.58609, 40.56463, 40.54297, 40.52111, 40.49904, 40.47678, 
    40.45431, 40.43164, 40.40878, 40.38571, 40.36245, 40.33898, 40.31532, 
    40.29146, 40.2674, 40.24314, 40.21869, 40.19403, 40.16919, 40.14414, 
    40.1189, 40.09346, 40.06783, 40.042, 40.01597, 39.98975, 39.96334, 
    39.93673, 39.90993, 39.88293, 39.85574, 39.82836, 39.80079, 39.77302, 
    39.74506, 39.71692, 39.68857, 39.66004, 39.63132, 39.60241, 39.5733, 
    39.54401, 39.51453, 39.48486, 39.455, 39.42495, 39.39471, 39.36429, 
    39.33368, 39.30289, 39.2719, 39.24073, 39.20938, 39.17784, 39.14611, 
    39.1142, 39.08211, 39.04983, 39.01737, 38.98472, 38.95189, 38.91888, 
    38.88569, 38.85231, 38.81876, 38.78502, 38.7511, 38.71701, 38.68273, 
    38.64827, 38.61363,
  34.76873, 34.81837, 34.86787, 34.91722, 34.96643, 35.0155, 35.06441, 
    35.11319, 35.16182, 35.21031, 35.25865, 35.30685, 35.3549, 35.4028, 
    35.45055, 35.49816, 35.54562, 35.59293, 35.64009, 35.6871, 35.73397, 
    35.78068, 35.82724, 35.87365, 35.91991, 35.96602, 36.01198, 36.05778, 
    36.10343, 36.14893, 36.19427, 36.23946, 36.2845, 36.32938, 36.3741, 
    36.41867, 36.46308, 36.50734, 36.55144, 36.59538, 36.63916, 36.68279, 
    36.72625, 36.76956, 36.81271, 36.8557, 36.89853, 36.94119, 36.9837, 
    37.02605, 37.06823, 37.11025, 37.15211, 37.19381, 37.23534, 37.2767, 
    37.31791, 37.35895, 37.39982, 37.44053, 37.48107, 37.52145, 37.56166, 
    37.6017, 37.64158, 37.68129, 37.72083, 37.76019, 37.7994, 37.83843, 
    37.87729, 37.91598, 37.95451, 37.99286, 38.03103, 38.06904, 38.10688, 
    38.14454, 38.18203, 38.21935, 38.25648, 38.29345, 38.33025, 38.36687, 
    38.40331, 38.43958, 38.47567, 38.51159, 38.54733, 38.58289, 38.61827, 
    38.65348, 38.6885, 38.72335, 38.75802, 38.79251, 38.82682, 38.86095, 
    38.8949, 38.92867, 38.96226, 38.99566, 39.02888, 39.06193, 39.09478, 
    39.12746, 39.15995, 39.19226, 39.22438, 39.25632, 39.28807, 39.31964, 
    39.35102, 39.38222, 39.41323, 39.44405, 39.47469, 39.50514, 39.5354, 
    39.56547, 39.59536, 39.62505, 39.65456, 39.68387, 39.713, 39.74194, 
    39.77068, 39.79923, 39.8276, 39.85577, 39.88375, 39.91154, 39.93913, 
    39.96653, 39.99374, 40.02076, 40.04758, 40.07421, 40.10064, 40.12688, 
    40.15292, 40.17876, 40.20442, 40.22987, 40.25513, 40.28019, 40.30506, 
    40.32972, 40.35419, 40.37847, 40.40254, 40.42641, 40.45009, 40.47357, 
    40.49685, 40.51992, 40.5428, 40.56548, 40.58796, 40.61023, 40.63231, 
    40.65418, 40.67585, 40.69733, 40.71859, 40.73966, 40.76052, 40.78118, 
    40.80164, 40.82189, 40.84194, 40.86179, 40.88142, 40.90086, 40.92009, 
    40.93912, 40.95794, 40.97655, 40.99496, 41.01317, 41.03116, 41.04895, 
    41.06654, 41.08392, 41.10109, 41.11805, 41.1348, 41.15135, 41.16769, 
    41.18382, 41.19974, 41.21545, 41.23096, 41.24625, 41.26134, 41.27621, 
    41.29088, 41.30534, 41.31958, 41.33362, 41.34745, 41.36106, 41.37447, 
    41.38766, 41.40064, 41.41341, 41.42597, 41.43832, 41.45045, 41.46238, 
    41.47409, 41.48558, 41.49687, 41.50794, 41.51881, 41.52945, 41.53989, 
    41.55011, 41.56012, 41.56991, 41.57949, 41.58886, 41.59801, 41.60695, 
    41.61567, 41.62418, 41.63248, 41.64056, 41.64843, 41.65608, 41.66352, 
    41.67074, 41.67775, 41.68454, 41.69112, 41.69748, 41.70362, 41.70956, 
    41.71527, 41.72077, 41.72606, 41.73112, 41.73597, 41.74061, 41.74503, 
    41.74923, 41.75322, 41.75699, 41.76055, 41.76389, 41.76701, 41.76992, 
    41.77261, 41.77508, 41.77734, 41.77938, 41.7812, 41.78281, 41.7842, 
    41.78538, 41.78633, 41.78708, 41.7876, 41.78791, 41.788, 41.78787, 
    41.78753, 41.78697, 41.7862, 41.78521, 41.784, 41.78257, 41.78093, 
    41.77907, 41.777, 41.7747, 41.7722, 41.76947, 41.76653, 41.76337, 41.76, 
    41.75641, 41.75261, 41.74858, 41.74435, 41.73989, 41.73522, 41.73034, 
    41.72523, 41.71991, 41.71438, 41.70863, 41.70267, 41.69649, 41.69009, 
    41.68348, 41.67665, 41.66961, 41.66236, 41.65488, 41.6472, 41.6393, 
    41.63118, 41.62285, 41.61431, 41.60555, 41.59658, 41.58739, 41.57799, 
    41.56837, 41.55855, 41.5485, 41.53825, 41.52778, 41.5171, 41.50621, 
    41.4951, 41.48378, 41.47225, 41.4605, 41.44855, 41.43638, 41.424, 
    41.4114, 41.3986, 41.38559, 41.37236, 41.35892, 41.34527, 41.33141, 
    41.31734, 41.30306, 41.28857, 41.27388, 41.25896, 41.24385, 41.22852, 
    41.21298, 41.19724, 41.18128, 41.16512, 41.14875, 41.13216, 41.11538, 
    41.09838, 41.08118, 41.06377, 41.04615, 41.02833, 41.0103, 40.99207, 
    40.97363, 40.95498, 40.93612, 40.91706, 40.8978, 40.87833, 40.85866, 
    40.83878, 40.8187, 40.79842, 40.77793, 40.75724, 40.73634, 40.71524, 
    40.69394, 40.67244, 40.65074, 40.62883, 40.60672, 40.58442, 40.56191, 
    40.5392, 40.51629, 40.49318, 40.46987, 40.44636, 40.42265, 40.39875, 
    40.37464, 40.35034, 40.32584, 40.30114, 40.27624, 40.25115, 40.22586, 
    40.20037, 40.17469, 40.14881, 40.12274, 40.09647, 40.07001, 40.04335, 
    40.0165, 39.98945, 39.96221, 39.93478, 39.90715, 39.87934, 39.85133, 
    39.82312, 39.79473, 39.76614, 39.73737, 39.7084, 39.67924, 39.6499, 
    39.62037, 39.59064, 39.56073, 39.53062, 39.50033, 39.46986, 39.43919, 
    39.40834, 39.3773, 39.34607, 39.31466, 39.28306, 39.25128, 39.21931, 
    39.18716, 39.15482, 39.1223, 39.0896, 39.05671, 39.02364, 38.99039, 
    38.95695, 38.92334, 38.88954, 38.85556, 38.82141, 38.78707, 38.75255, 
    38.71785,
  34.86653, 34.91624, 34.96581, 35.01524, 35.06452, 35.11366, 35.16266, 
    35.21151, 35.26021, 35.30877, 35.35719, 35.40546, 35.45358, 35.50155, 
    35.54938, 35.59706, 35.6446, 35.69198, 35.73921, 35.7863, 35.83323, 
    35.88002, 35.92665, 35.97314, 36.01947, 36.06565, 36.11168, 36.15755, 
    36.20327, 36.24884, 36.29426, 36.33952, 36.38462, 36.42958, 36.47437, 
    36.51901, 36.5635, 36.60782, 36.65199, 36.696, 36.73986, 36.78355, 
    36.82709, 36.87047, 36.91368, 36.95675, 36.99964, 37.04238, 37.08496, 
    37.12737, 37.16962, 37.21171, 37.25364, 37.29541, 37.33701, 37.37844, 
    37.41972, 37.46082, 37.50176, 37.54254, 37.58315, 37.6236, 37.66387, 
    37.70398, 37.74392, 37.7837, 37.8233, 37.86274, 37.90201, 37.94111, 
    37.98004, 38.0188, 38.05738, 38.0958, 38.13404, 38.17212, 38.21001, 
    38.24774, 38.2853, 38.32268, 38.35988, 38.39692, 38.43377, 38.47046, 
    38.50696, 38.54329, 38.57945, 38.61543, 38.65123, 38.68685, 38.7223, 
    38.75756, 38.79265, 38.82756, 38.86229, 38.89684, 38.93122, 38.9654, 
    38.99942, 39.03325, 39.06689, 39.10036, 39.13364, 39.16674, 39.19966, 
    39.23239, 39.26494, 39.29731, 39.32949, 39.36148, 39.39329, 39.42492, 
    39.45636, 39.48761, 39.51868, 39.54956, 39.58025, 39.61075, 39.64107, 
    39.6712, 39.70113, 39.73088, 39.76044, 39.78981, 39.81899, 39.84798, 
    39.87678, 39.90539, 39.9338, 39.96203, 39.99006, 40.0179, 40.04554, 
    40.073, 40.10026, 40.12732, 40.15419, 40.18087, 40.20735, 40.23364, 
    40.25973, 40.28563, 40.31133, 40.33683, 40.36214, 40.38725, 40.41216, 
    40.43687, 40.46139, 40.48571, 40.50983, 40.53374, 40.55747, 40.58099, 
    40.60431, 40.62743, 40.65036, 40.67308, 40.69559, 40.71791, 40.74003, 
    40.76195, 40.78366, 40.80518, 40.82648, 40.84759, 40.86849, 40.88919, 
    40.90969, 40.92998, 40.95007, 40.96995, 40.98963, 41.0091, 41.02837, 
    41.04744, 41.06629, 41.08494, 41.10339, 41.12163, 41.13966, 41.15749, 
    41.1751, 41.19251, 41.20972, 41.22671, 41.2435, 41.26008, 41.27645, 
    41.29261, 41.30857, 41.32431, 41.33984, 41.35517, 41.37029, 41.38519, 
    41.39989, 41.41437, 41.42865, 41.44271, 41.45656, 41.47021, 41.48363, 
    41.49686, 41.50986, 41.52266, 41.53524, 41.54762, 41.55977, 41.57172, 
    41.58345, 41.59498, 41.60629, 41.61738, 41.62827, 41.63893, 41.64939, 
    41.65963, 41.66966, 41.67947, 41.68907, 41.69846, 41.70763, 41.71658, 
    41.72533, 41.73386, 41.74217, 41.75027, 41.75815, 41.76582, 41.77327, 
    41.78051, 41.78753, 41.79433, 41.80092, 41.8073, 41.81345, 41.8194, 
    41.82512, 41.83064, 41.83593, 41.84101, 41.84587, 41.85051, 41.85494, 
    41.85916, 41.86315, 41.86693, 41.87049, 41.87384, 41.87697, 41.87988, 
    41.88258, 41.88506, 41.88732, 41.88936, 41.89119, 41.8928, 41.8942, 
    41.89537, 41.89633, 41.89708, 41.8976, 41.89791, 41.898, 41.89787, 
    41.89753, 41.89697, 41.89619, 41.8952, 41.89399, 41.89256, 41.89091, 
    41.88905, 41.88697, 41.88468, 41.88216, 41.87944, 41.87649, 41.87333, 
    41.86995, 41.86635, 41.86253, 41.85851, 41.85426, 41.84979, 41.84512, 
    41.84022, 41.83511, 41.82978, 41.82423, 41.81847, 41.8125, 41.8063, 
    41.79989, 41.79327, 41.78643, 41.77937, 41.7721, 41.76462, 41.75692, 
    41.749, 41.74087, 41.73252, 41.72396, 41.71518, 41.70619, 41.69699, 
    41.68757, 41.67793, 41.66809, 41.65802, 41.64775, 41.63726, 41.62656, 
    41.61564, 41.60451, 41.59317, 41.58161, 41.56985, 41.55787, 41.54567, 
    41.53327, 41.52065, 41.50782, 41.49478, 41.48153, 41.46806, 41.45439, 
    41.4405, 41.4264, 41.41209, 41.39758, 41.38285, 41.36791, 41.35276, 
    41.3374, 41.32183, 41.30606, 41.29007, 41.27388, 41.25747, 41.24086, 
    41.22404, 41.20701, 41.18977, 41.17233, 41.15468, 41.13682, 41.11876, 
    41.10048, 41.08201, 41.06332, 41.04443, 41.02534, 41.00603, 40.98653, 
    40.96682, 40.9469, 40.92678, 40.90646, 40.88593, 40.8652, 40.84426, 
    40.82312, 40.80178, 40.78024, 40.7585, 40.73655, 40.7144, 40.69205, 
    40.66949, 40.64674, 40.62379, 40.60064, 40.57728, 40.55373, 40.52998, 
    40.50602, 40.48187, 40.45752, 40.43298, 40.40823, 40.38329, 40.35815, 
    40.33281, 40.30727, 40.28154, 40.25562, 40.2295, 40.20318, 40.17666, 
    40.14996, 40.12305, 40.09596, 40.06867, 40.04118, 40.01351, 39.98564, 
    39.95758, 39.92932, 39.90088, 39.87224, 39.84341, 39.81439, 39.78518, 
    39.75578, 39.72619, 39.69641, 39.66644, 39.63628, 39.60594, 39.57541, 
    39.54468, 39.51377, 39.48268, 39.4514, 39.41993, 39.38827, 39.35643, 
    39.32441, 39.2922, 39.2598, 39.22722, 39.19446, 39.16151, 39.12839, 
    39.09507, 39.06158, 39.0279, 38.99405, 38.96001, 38.92579, 38.89139, 
    38.85681, 38.82205,
  34.9643, 35.01409, 35.06373, 35.11323, 35.16259, 35.2118, 35.26087, 
    35.30979, 35.35857, 35.40721, 35.4557, 35.50404, 35.55223, 35.60028, 
    35.64818, 35.69593, 35.74354, 35.791, 35.8383, 35.88546, 35.93247, 
    35.97933, 36.02604, 36.07259, 36.119, 36.16525, 36.21135, 36.25729, 
    36.30309, 36.34873, 36.39422, 36.43955, 36.48473, 36.52975, 36.57462, 
    36.61933, 36.66388, 36.70828, 36.75252, 36.7966, 36.84053, 36.8843, 
    36.9279, 36.97135, 37.01464, 37.05777, 37.10073, 37.14354, 37.18619, 
    37.22867, 37.27099, 37.31315, 37.35515, 37.39698, 37.43865, 37.48016, 
    37.5215, 37.56268, 37.60368, 37.64453, 37.68521, 37.72572, 37.76606, 
    37.80624, 37.84625, 37.88609, 37.92577, 37.96527, 38.0046, 38.04377, 
    38.08276, 38.12159, 38.16024, 38.19872, 38.23703, 38.27517, 38.31313, 
    38.35093, 38.38854, 38.42599, 38.46326, 38.50035, 38.53728, 38.57402, 
    38.61059, 38.64699, 38.6832, 38.71925, 38.75511, 38.79079, 38.82631, 
    38.86163, 38.89679, 38.93176, 38.96655, 39.00116, 39.03559, 39.06984, 
    39.10391, 39.1378, 39.17151, 39.20504, 39.23838, 39.27153, 39.30451, 
    39.3373, 39.36991, 39.40234, 39.43457, 39.46663, 39.4985, 39.53018, 
    39.56168, 39.59299, 39.62411, 39.65504, 39.68579, 39.71635, 39.74672, 
    39.77691, 39.8069, 39.8367, 39.86632, 39.89574, 39.92498, 39.95402, 
    39.98287, 40.01153, 40.04, 40.06828, 40.09636, 40.12425, 40.15195, 
    40.17945, 40.20676, 40.23388, 40.2608, 40.28753, 40.31406, 40.34039, 
    40.36654, 40.39248, 40.41823, 40.44378, 40.46913, 40.49429, 40.51925, 
    40.54401, 40.56857, 40.59293, 40.6171, 40.64107, 40.66483, 40.6884, 
    40.71177, 40.73493, 40.7579, 40.78066, 40.80323, 40.82559, 40.84775, 
    40.86971, 40.89146, 40.91301, 40.93436, 40.95551, 40.97646, 40.9972, 
    41.01773, 41.03806, 41.05819, 41.07811, 41.09783, 41.11734, 41.13665, 
    41.15575, 41.17464, 41.19333, 41.21181, 41.23008, 41.24815, 41.26601, 
    41.28366, 41.30111, 41.31834, 41.33537, 41.3522, 41.3688, 41.38521, 
    41.40141, 41.41739, 41.43316, 41.44873, 41.46408, 41.47923, 41.49416, 
    41.50889, 41.5234, 41.5377, 41.5518, 41.56568, 41.57935, 41.5928, 
    41.60605, 41.61908, 41.6319, 41.64452, 41.65691, 41.66909, 41.68106, 
    41.69282, 41.70437, 41.7157, 41.72682, 41.73772, 41.74841, 41.75889, 
    41.76915, 41.7792, 41.78903, 41.79865, 41.80806, 41.81725, 41.82622, 
    41.83498, 41.84352, 41.85185, 41.85997, 41.86787, 41.87555, 41.88301, 
    41.89027, 41.8973, 41.90412, 41.91072, 41.91711, 41.92328, 41.92924, 
    41.93498, 41.9405, 41.9458, 41.95089, 41.95576, 41.96042, 41.96486, 
    41.96908, 41.97308, 41.97687, 41.98044, 41.98379, 41.98693, 41.98985, 
    41.99255, 41.99503, 41.9973, 41.99934, 42.00117, 42.00279, 42.00419, 
    42.00537, 42.00633, 42.00707, 42.0076, 42.00791, 42.008, 42.00787, 
    42.00753, 42.00697, 42.00619, 42.0052, 42.00398, 42.00255, 42.0009, 
    41.99903, 41.99695, 41.99465, 41.99213, 41.9894, 41.98645, 41.98328, 
    41.97989, 41.97628, 41.97246, 41.96843, 41.96417, 41.9597, 41.95501, 
    41.9501, 41.94498, 41.93964, 41.93408, 41.92831, 41.92232, 41.91612, 
    41.90969, 41.90306, 41.89621, 41.88913, 41.88185, 41.87435, 41.86663, 
    41.8587, 41.85055, 41.84219, 41.83361, 41.82481, 41.8158, 41.80658, 
    41.79714, 41.78749, 41.77762, 41.76754, 41.75724, 41.74673, 41.73601, 
    41.72507, 41.71392, 41.70256, 41.69098, 41.67919, 41.66718, 41.65496, 
    41.64253, 41.62989, 41.61703, 41.60397, 41.59069, 41.5772, 41.5635, 
    41.54958, 41.53546, 41.52112, 41.50657, 41.49182, 41.47685, 41.46167, 
    41.44628, 41.43068, 41.41488, 41.39886, 41.38263, 41.36619, 41.34955, 
    41.3327, 41.31563, 41.29836, 41.28088, 41.2632, 41.24531, 41.22721, 
    41.2089, 41.19038, 41.17167, 41.15274, 41.13361, 41.11427, 41.09472, 
    41.07497, 41.05502, 41.03486, 41.0145, 40.99393, 40.97316, 40.95218, 
    40.931, 40.90962, 40.88803, 40.86625, 40.84426, 40.82206, 40.79967, 
    40.77708, 40.75428, 40.73128, 40.70808, 40.68468, 40.66109, 40.63729, 
    40.61329, 40.5891, 40.5647, 40.5401, 40.51531, 40.49032, 40.46513, 
    40.43975, 40.41417, 40.38839, 40.36241, 40.33624, 40.30988, 40.28331, 
    40.25655, 40.2296, 40.20245, 40.17511, 40.14758, 40.11985, 40.09193, 
    40.06382, 40.03551, 40.00701, 39.97832, 39.94944, 39.92036, 39.8911, 
    39.86164, 39.832, 39.80217, 39.77214, 39.74193, 39.71153, 39.68094, 
    39.65016, 39.6192, 39.58805, 39.55671, 39.52518, 39.49347, 39.46157, 
    39.42949, 39.39722, 39.36477, 39.33213, 39.29931, 39.2663, 39.23312, 
    39.19975, 39.16619, 39.13245, 39.09854, 39.06444, 39.03016, 38.9957, 
    38.96106, 38.92624,
  35.06204, 35.1119, 35.16161, 35.21119, 35.26062, 35.30991, 35.35905, 
    35.40805, 35.4569, 35.50561, 35.55417, 35.60259, 35.65086, 35.69898, 
    35.74695, 35.79478, 35.84246, 35.88999, 35.93737, 35.9846, 36.03168, 
    36.07861, 36.12539, 36.17202, 36.21849, 36.26482, 36.31099, 36.35701, 
    36.40288, 36.44859, 36.49415, 36.53955, 36.5848, 36.6299, 36.67484, 
    36.71962, 36.76424, 36.80871, 36.85302, 36.89718, 36.94117, 36.98501, 
    37.02869, 37.07221, 37.11557, 37.15876, 37.2018, 37.24468, 37.2874, 
    37.32995, 37.37234, 37.41457, 37.45663, 37.49854, 37.54028, 37.58185, 
    37.62326, 37.6645, 37.70558, 37.74649, 37.78724, 37.82782, 37.86823, 
    37.90848, 37.94855, 37.98846, 38.0282, 38.06777, 38.10717, 38.1464, 
    38.18547, 38.22436, 38.26307, 38.30162, 38.34, 38.3782, 38.41623, 
    38.45409, 38.49177, 38.52928, 38.56662, 38.60378, 38.64076, 38.67757, 
    38.71421, 38.75066, 38.78695, 38.82305, 38.85897, 38.89473, 38.93029, 
    38.96569, 39.0009, 39.03593, 39.07079, 39.10546, 39.13995, 39.17426, 
    39.2084, 39.24234, 39.27611, 39.3097, 39.3431, 39.37632, 39.40935, 
    39.4422, 39.47487, 39.50735, 39.53965, 39.57176, 39.60369, 39.63543, 
    39.66698, 39.69835, 39.72953, 39.76052, 39.79132, 39.82194, 39.85236, 
    39.8826, 39.91265, 39.94251, 39.97218, 40.00166, 40.03094, 40.06004, 
    40.08895, 40.11766, 40.14618, 40.17451, 40.20264, 40.23059, 40.25834, 
    40.28589, 40.31326, 40.34042, 40.36739, 40.39417, 40.42075, 40.44714, 
    40.47333, 40.49932, 40.52512, 40.55072, 40.57612, 40.60132, 40.62633, 
    40.65114, 40.67575, 40.70016, 40.72437, 40.74838, 40.77219, 40.7958, 
    40.81921, 40.84243, 40.86543, 40.88824, 40.91085, 40.93325, 40.95546, 
    40.97746, 40.99926, 41.02085, 41.04224, 41.06343, 41.08441, 41.10519, 
    41.12577, 41.14614, 41.1663, 41.18626, 41.20602, 41.22557, 41.24491, 
    41.26405, 41.28298, 41.3017, 41.32022, 41.33853, 41.35664, 41.37453, 
    41.39222, 41.4097, 41.42697, 41.44403, 41.46088, 41.47753, 41.49397, 
    41.51019, 41.52621, 41.54201, 41.55761, 41.57299, 41.58817, 41.60313, 
    41.61789, 41.63243, 41.64676, 41.66088, 41.67479, 41.68849, 41.70197, 
    41.71524, 41.7283, 41.74115, 41.75378, 41.7662, 41.77841, 41.79041, 
    41.80219, 41.81376, 41.82511, 41.83625, 41.84718, 41.85789, 41.86839, 
    41.87867, 41.88874, 41.89859, 41.90823, 41.91765, 41.92686, 41.93585, 
    41.94463, 41.95319, 41.96154, 41.96967, 41.97758, 41.98528, 41.99276, 
    42.00003, 42.00708, 42.01391, 42.02053, 42.02693, 42.03311, 42.03908, 
    42.04483, 42.05036, 42.05568, 42.06078, 42.06566, 42.07032, 42.07477, 
    42.079, 42.08301, 42.0868, 42.09038, 42.09374, 42.09689, 42.09981, 
    42.10252, 42.105, 42.10727, 42.10933, 42.11116, 42.11278, 42.11418, 
    42.11536, 42.11633, 42.11707, 42.1176, 42.11791, 42.118, 42.11787, 
    42.11753, 42.11697, 42.11619, 42.11519, 42.11397, 42.11254, 42.11089, 
    42.10902, 42.10693, 42.10463, 42.1021, 42.09936, 42.0964, 42.09322, 
    42.08983, 42.08622, 42.08239, 42.07834, 42.07408, 42.0696, 42.0649, 
    42.05998, 42.05485, 42.0495, 42.04393, 42.03815, 42.03215, 42.02593, 
    42.0195, 42.01284, 42.00598, 41.99889, 41.99159, 41.98408, 41.97635, 
    41.9684, 41.96023, 41.95185, 41.94326, 41.93444, 41.92542, 41.91618, 
    41.90672, 41.89705, 41.88716, 41.87706, 41.86674, 41.85621, 41.84546, 
    41.8345, 41.82333, 41.81194, 41.80034, 41.78852, 41.7765, 41.76426, 
    41.7518, 41.73913, 41.72625, 41.71316, 41.69985, 41.68633, 41.6726, 
    41.65866, 41.64451, 41.63015, 41.61557, 41.60078, 41.58578, 41.57058, 
    41.55516, 41.53953, 41.52369, 41.50764, 41.49138, 41.47491, 41.45823, 
    41.44135, 41.42425, 41.40695, 41.38943, 41.37172, 41.35379, 41.33565, 
    41.31731, 41.29876, 41.28, 41.26104, 41.24187, 41.22249, 41.20291, 
    41.18312, 41.16313, 41.14293, 41.12252, 41.10192, 41.0811, 41.06009, 
    41.03887, 41.01745, 40.99582, 40.97399, 40.95196, 40.92972, 40.90729, 
    40.88465, 40.86181, 40.83877, 40.81553, 40.79208, 40.76844, 40.74459, 
    40.72055, 40.69631, 40.67187, 40.64722, 40.62239, 40.59735, 40.57211, 
    40.54668, 40.52105, 40.49522, 40.4692, 40.44298, 40.41656, 40.38995, 
    40.36314, 40.33614, 40.30894, 40.28155, 40.25396, 40.22618, 40.19821, 
    40.17004, 40.14168, 40.11313, 40.08438, 40.05545, 40.02633, 39.99701, 
    39.9675, 39.9378, 39.90791, 39.87783, 39.84756, 39.81711, 39.78646, 
    39.75563, 39.72461, 39.6934, 39.662, 39.63042, 39.59865, 39.56669, 
    39.53455, 39.50223, 39.46972, 39.43702, 39.40414, 39.37107, 39.33783, 
    39.3044, 39.27078, 39.23699, 39.20301, 39.16885, 39.13451, 39.09999, 
    39.06528, 39.0304,
  35.15974, 35.20968, 35.25947, 35.30912, 35.35862, 35.40798, 35.4572, 
    35.50627, 35.5552, 35.60398, 35.65262, 35.70111, 35.74945, 35.79765, 
    35.84569, 35.89359, 35.94135, 35.98895, 36.0364, 36.08371, 36.13086, 
    36.17786, 36.22472, 36.27142, 36.31797, 36.36436, 36.41061, 36.4567, 
    36.50264, 36.54842, 36.59406, 36.63953, 36.68485, 36.73002, 36.77503, 
    36.81988, 36.86458, 36.90912, 36.9535, 36.99773, 37.04179, 37.0857, 
    37.12945, 37.17304, 37.21647, 37.25974, 37.30285, 37.34579, 37.38858, 
    37.4312, 37.47366, 37.51596, 37.55809, 37.60007, 37.64187, 37.68352, 
    37.72499, 37.76631, 37.80745, 37.84843, 37.88925, 37.9299, 37.97038, 
    38.01069, 38.05083, 38.09081, 38.13062, 38.17025, 38.20972, 38.24902, 
    38.28815, 38.32711, 38.36589, 38.4045, 38.44294, 38.48121, 38.51931, 
    38.55723, 38.59498, 38.63255, 38.66995, 38.70718, 38.74423, 38.7811, 
    38.8178, 38.85432, 38.89067, 38.92683, 38.96282, 38.99863, 39.03427, 
    39.06972, 39.105, 39.14009, 39.17501, 39.20974, 39.2443, 39.27867, 
    39.31286, 39.34687, 39.3807, 39.41434, 39.4478, 39.48108, 39.51418, 
    39.54708, 39.57981, 39.61235, 39.64471, 39.67688, 39.70886, 39.74066, 
    39.77227, 39.80369, 39.83493, 39.86598, 39.89684, 39.92751, 39.95799, 
    39.98829, 40.01839, 40.0483, 40.07803, 40.10756, 40.1369, 40.16605, 
    40.19501, 40.22378, 40.25235, 40.28073, 40.30892, 40.33691, 40.36472, 
    40.39232, 40.41973, 40.44695, 40.47398, 40.5008, 40.52744, 40.55387, 
    40.58011, 40.60615, 40.632, 40.65764, 40.68309, 40.70835, 40.7334, 
    40.75826, 40.78291, 40.80737, 40.83163, 40.85568, 40.87954, 40.9032, 
    40.92665, 40.94991, 40.97296, 40.99582, 41.01846, 41.04091, 41.06316, 
    41.0852, 41.10704, 41.12868, 41.15011, 41.17134, 41.19236, 41.21318, 
    41.2338, 41.25421, 41.27441, 41.29441, 41.31421, 41.33379, 41.35318, 
    41.37235, 41.39132, 41.41008, 41.42863, 41.44698, 41.46511, 41.48305, 
    41.50077, 41.51828, 41.53559, 41.55268, 41.56957, 41.58625, 41.60271, 
    41.61897, 41.63502, 41.65086, 41.66648, 41.6819, 41.69711, 41.7121, 
    41.72688, 41.74146, 41.75582, 41.76996, 41.7839, 41.79762, 41.81113, 
    41.82443, 41.83752, 41.85039, 41.86305, 41.8755, 41.88773, 41.89975, 
    41.91155, 41.92314, 41.93452, 41.94568, 41.95663, 41.96736, 41.97788, 
    41.98819, 41.99827, 42.00814, 42.0178, 42.02724, 42.03647, 42.04548, 
    42.05428, 42.06286, 42.07122, 42.07937, 42.0873, 42.09501, 42.10251, 
    42.10979, 42.11686, 42.1237, 42.13033, 42.13675, 42.14294, 42.14892, 
    42.15468, 42.16022, 42.16555, 42.17066, 42.17555, 42.18023, 42.18468, 
    42.18892, 42.19294, 42.19674, 42.20033, 42.20369, 42.20684, 42.20977, 
    42.21248, 42.21498, 42.21725, 42.21931, 42.22115, 42.22277, 42.22417, 
    42.22536, 42.22632, 42.22707, 42.2276, 42.22791, 42.228, 42.22787, 
    42.22753, 42.22696, 42.22618, 42.22518, 42.22396, 42.22253, 42.22087, 
    42.219, 42.21691, 42.2146, 42.21207, 42.20932, 42.20636, 42.20317, 
    42.19978, 42.19616, 42.19232, 42.18826, 42.18399, 42.1795, 42.17479, 
    42.16986, 42.16472, 42.15936, 42.15378, 42.14799, 42.14198, 42.13575, 
    42.1293, 42.12263, 42.11575, 42.10865, 42.10134, 42.09381, 42.08606, 
    42.07809, 42.06991, 42.06152, 42.0529, 42.04407, 42.03503, 42.02577, 
    42.01629, 42.0066, 41.99669, 41.98657, 41.97623, 41.96568, 41.95491, 
    41.94393, 41.93274, 41.92132, 41.9097, 41.89786, 41.88581, 41.87354, 
    41.86106, 41.84837, 41.83546, 41.82234, 41.80901, 41.79547, 41.78171, 
    41.76774, 41.75356, 41.73917, 41.72456, 41.70974, 41.69472, 41.67948, 
    41.66403, 41.64837, 41.6325, 41.61642, 41.60012, 41.58362, 41.56691, 
    41.54999, 41.53286, 41.51553, 41.49798, 41.48022, 41.46226, 41.44409, 
    41.42571, 41.40712, 41.38833, 41.36933, 41.35012, 41.33071, 41.31109, 
    41.29126, 41.27123, 41.25099, 41.23055, 41.2099, 41.18905, 41.16799, 
    41.14673, 41.12527, 41.1036, 41.08173, 41.05965, 41.03738, 41.0149, 
    40.99221, 40.96933, 40.94624, 40.92296, 40.89947, 40.87578, 40.85189, 
    40.8278, 40.80351, 40.77903, 40.75434, 40.72945, 40.70436, 40.67908, 
    40.6536, 40.62792, 40.60204, 40.57597, 40.5497, 40.52324, 40.49657, 
    40.46972, 40.44266, 40.41541, 40.38797, 40.36033, 40.3325, 40.30447, 
    40.27626, 40.24784, 40.21924, 40.19044, 40.16145, 40.13227, 40.1029, 
    40.07334, 40.04358, 40.01364, 39.98351, 39.95318, 39.92267, 39.89197, 
    39.86108, 39.83, 39.79874, 39.76728, 39.73564, 39.70382, 39.6718, 
    39.6396, 39.60722, 39.57465, 39.54189, 39.50895, 39.47583, 39.44252, 
    39.40903, 39.37536, 39.3415, 39.30746, 39.27324, 39.23884, 39.20426, 
    39.16949, 39.13455,
  35.25742, 35.30743, 35.35729, 35.40702, 35.45659, 35.50603, 35.55532, 
    35.60447, 35.65347, 35.70232, 35.75103, 35.7996, 35.84801, 35.89628, 
    35.9444, 35.99238, 36.0402, 36.08788, 36.13541, 36.18278, 36.23001, 
    36.27709, 36.32401, 36.37078, 36.41741, 36.46388, 36.5102, 36.55636, 
    36.60237, 36.64823, 36.69393, 36.73948, 36.78487, 36.83011, 36.87519, 
    36.92012, 36.96489, 37.0095, 37.05396, 37.09825, 37.14239, 37.18637, 
    37.23019, 37.27385, 37.31734, 37.36068, 37.40386, 37.44688, 37.48973, 
    37.53243, 37.57496, 37.61733, 37.65953, 37.70157, 37.74345, 37.78516, 
    37.82671, 37.86809, 37.90931, 37.95036, 37.99124, 38.03195, 38.0725, 
    38.11288, 38.1531, 38.19314, 38.23301, 38.27272, 38.31225, 38.35162, 
    38.39081, 38.42983, 38.46869, 38.50736, 38.54587, 38.58421, 38.62236, 
    38.66035, 38.69817, 38.73581, 38.77327, 38.81056, 38.84768, 38.88461, 
    38.92138, 38.95796, 38.99437, 39.0306, 39.06665, 39.10252, 39.13822, 
    39.17374, 39.20907, 39.24423, 39.27921, 39.31401, 39.34862, 39.38306, 
    39.41731, 39.45138, 39.48526, 39.51897, 39.55249, 39.58583, 39.61898, 
    39.65195, 39.68474, 39.71734, 39.74975, 39.78198, 39.81402, 39.84587, 
    39.87754, 39.90903, 39.94032, 39.97142, 40.00234, 40.03307, 40.06361, 
    40.09396, 40.12411, 40.15408, 40.18386, 40.21345, 40.24284, 40.27205, 
    40.30106, 40.32988, 40.35851, 40.38694, 40.41518, 40.44323, 40.47108, 
    40.49874, 40.52621, 40.55347, 40.58055, 40.60743, 40.63411, 40.66059, 
    40.68688, 40.71297, 40.73886, 40.76456, 40.79006, 40.81536, 40.84046, 
    40.86536, 40.89007, 40.91457, 40.93887, 40.96298, 40.98688, 41.01058, 
    41.03408, 41.05738, 41.08048, 41.10338, 41.12607, 41.14856, 41.17085, 
    41.19294, 41.21482, 41.2365, 41.25797, 41.27924, 41.3003, 41.32116, 
    41.34182, 41.36227, 41.38251, 41.40255, 41.42239, 41.44201, 41.46143, 
    41.48064, 41.49965, 41.51844, 41.53704, 41.55542, 41.57359, 41.59156, 
    41.60931, 41.62686, 41.6442, 41.66133, 41.67825, 41.69496, 41.71146, 
    41.72775, 41.74383, 41.7597, 41.77536, 41.79081, 41.80604, 41.82106, 
    41.83588, 41.85048, 41.86486, 41.87904, 41.89301, 41.90676, 41.9203, 
    41.93362, 41.94673, 41.95963, 41.97231, 41.98478, 41.99704, 42.00908, 
    42.02091, 42.03253, 42.04393, 42.05511, 42.06608, 42.07684, 42.08738, 
    42.0977, 42.10781, 42.1177, 42.12738, 42.13684, 42.14608, 42.15511, 
    42.16393, 42.17252, 42.1809, 42.18907, 42.19701, 42.20474, 42.21225, 
    42.21955, 42.22663, 42.23349, 42.24013, 42.24656, 42.25277, 42.25876, 
    42.26453, 42.27009, 42.27542, 42.28054, 42.28545, 42.29013, 42.29459, 
    42.29884, 42.30287, 42.30668, 42.31027, 42.31364, 42.3168, 42.31973, 
    42.32245, 42.32495, 42.32723, 42.32929, 42.33113, 42.33276, 42.33416, 
    42.33535, 42.33632, 42.33707, 42.3376, 42.33791, 42.338, 42.33787, 
    42.33753, 42.33696, 42.33618, 42.33518, 42.33396, 42.33252, 42.33086, 
    42.32898, 42.32689, 42.32457, 42.32204, 42.31928, 42.31631, 42.31313, 
    42.30972, 42.30609, 42.30225, 42.29818, 42.2939, 42.2894, 42.28468, 
    42.27975, 42.27459, 42.26922, 42.26363, 42.25782, 42.2518, 42.24556, 
    42.2391, 42.23242, 42.22552, 42.21841, 42.21108, 42.20353, 42.19577, 
    42.18779, 42.17959, 42.17118, 42.16255, 42.1537, 42.14464, 42.13536, 
    42.12586, 42.11615, 42.10622, 42.09608, 42.08572, 42.07515, 42.06436, 
    42.05336, 42.04214, 42.0307, 42.01905, 42.00719, 41.99512, 41.98283, 
    41.97032, 41.9576, 41.94467, 41.93153, 41.91817, 41.90459, 41.89081, 
    41.87681, 41.8626, 41.84818, 41.83355, 41.8187, 41.80365, 41.78838, 
    41.7729, 41.7572, 41.7413, 41.72519, 41.70887, 41.69233, 41.67559, 
    41.65863, 41.64147, 41.6241, 41.60652, 41.58873, 41.57073, 41.55252, 
    41.53411, 41.51549, 41.49665, 41.47762, 41.45837, 41.43892, 41.41926, 
    41.3994, 41.37933, 41.35905, 41.33857, 41.31788, 41.29699, 41.27589, 
    41.25459, 41.23308, 41.21137, 41.18946, 41.16734, 41.14502, 41.12249, 
    41.09977, 41.07684, 41.05371, 41.03038, 41.00685, 40.98311, 40.95918, 
    40.93504, 40.91071, 40.88617, 40.86144, 40.83651, 40.81137, 40.78604, 
    40.76051, 40.73478, 40.70886, 40.68274, 40.65642, 40.6299, 40.60319, 
    40.57628, 40.54918, 40.52187, 40.49438, 40.46669, 40.43881, 40.41073, 
    40.38246, 40.35399, 40.32534, 40.29649, 40.26744, 40.23821, 40.20878, 
    40.17916, 40.14936, 40.11936, 40.08917, 40.05879, 40.02822, 39.99746, 
    39.96651, 39.93538, 39.90406, 39.87255, 39.84085, 39.80896, 39.77689, 
    39.74464, 39.71219, 39.67957, 39.64675, 39.61375, 39.58057, 39.5472, 
    39.51365, 39.47992, 39.446, 39.4119, 39.37762, 39.34316, 39.30851, 
    39.27369, 39.23868,
  35.35506, 35.40514, 35.45508, 35.50488, 35.55453, 35.60405, 35.65341, 
    35.70263, 35.75171, 35.80064, 35.84942, 35.89806, 35.94655, 35.99489, 
    36.04309, 36.09113, 36.13903, 36.18678, 36.23438, 36.28183, 36.32913, 
    36.37628, 36.42328, 36.47013, 36.51682, 36.56337, 36.60976, 36.65599, 
    36.70208, 36.74801, 36.79378, 36.8394, 36.88487, 36.93018, 36.97533, 
    37.02033, 37.06517, 37.10985, 37.15438, 37.19875, 37.24295, 37.287, 
    37.33089, 37.37463, 37.4182, 37.46161, 37.50486, 37.54794, 37.59087, 
    37.63363, 37.67623, 37.71867, 37.76094, 37.80305, 37.845, 37.88678, 
    37.9284, 37.96985, 38.01113, 38.05225, 38.0932, 38.13398, 38.1746, 
    38.21505, 38.25533, 38.29544, 38.33538, 38.37516, 38.41476, 38.45419, 
    38.49345, 38.53254, 38.57146, 38.6102, 38.64877, 38.68718, 38.7254, 
    38.76345, 38.80133, 38.83904, 38.87657, 38.91392, 38.9511, 38.9881, 
    39.02493, 39.06158, 39.09805, 39.13434, 39.17046, 39.2064, 39.24216, 
    39.27774, 39.31313, 39.34835, 39.38339, 39.41825, 39.45293, 39.48742, 
    39.52174, 39.55587, 39.58982, 39.62358, 39.65717, 39.69056, 39.72377, 
    39.75681, 39.78965, 39.82231, 39.85478, 39.88707, 39.91917, 39.95108, 
    39.9828, 40.01434, 40.04569, 40.07685, 40.10783, 40.13861, 40.16921, 
    40.19961, 40.22983, 40.25985, 40.28968, 40.31932, 40.34877, 40.37803, 
    40.4071, 40.43597, 40.46465, 40.49314, 40.52143, 40.54953, 40.57744, 
    40.60515, 40.63266, 40.65998, 40.68711, 40.71404, 40.74077, 40.7673, 
    40.79364, 40.81978, 40.84573, 40.87147, 40.89702, 40.92237, 40.94751, 
    40.97247, 40.99722, 41.02176, 41.04612, 41.07026, 41.09421, 41.11796, 
    41.14151, 41.16485, 41.18799, 41.21093, 41.23367, 41.25621, 41.27854, 
    41.30066, 41.32259, 41.34431, 41.36582, 41.38713, 41.40824, 41.42914, 
    41.44984, 41.47033, 41.49061, 41.51069, 41.53056, 41.55022, 41.56968, 
    41.58893, 41.60797, 41.62681, 41.64544, 41.66385, 41.68206, 41.70006, 
    41.71785, 41.73544, 41.75281, 41.76997, 41.78693, 41.80367, 41.8202, 
    41.83652, 41.85264, 41.86854, 41.88423, 41.8997, 41.91497, 41.93002, 
    41.94487, 41.9595, 41.97391, 41.98812, 42.00211, 42.01589, 42.02945, 
    42.0428, 42.05594, 42.06887, 42.08157, 42.09407, 42.10635, 42.11842, 
    42.13027, 42.14191, 42.15333, 42.16454, 42.17553, 42.18631, 42.19687, 
    42.20721, 42.21734, 42.22725, 42.23695, 42.24643, 42.2557, 42.26474, 
    42.27357, 42.28219, 42.29058, 42.29876, 42.30673, 42.31447, 42.322, 
    42.32931, 42.3364, 42.34328, 42.34993, 42.35637, 42.36259, 42.3686, 
    42.37438, 42.37995, 42.3853, 42.39043, 42.39534, 42.40003, 42.40451, 
    42.40876, 42.4128, 42.41661, 42.42021, 42.4236, 42.42675, 42.4297, 
    42.43242, 42.43493, 42.43721, 42.43927, 42.44112, 42.44275, 42.44416, 
    42.44534, 42.44632, 42.44706, 42.44759, 42.44791, 42.448, 42.44787, 
    42.44753, 42.44696, 42.44617, 42.44517, 42.44395, 42.4425, 42.44084, 
    42.43896, 42.43686, 42.43454, 42.432, 42.42924, 42.42627, 42.42307, 
    42.41966, 42.41603, 42.41217, 42.4081, 42.40381, 42.3993, 42.39458, 
    42.38963, 42.38446, 42.37908, 42.37348, 42.36766, 42.36163, 42.35537, 
    42.3489, 42.34221, 42.3353, 42.32817, 42.32082, 42.31326, 42.30548, 
    42.29749, 42.28927, 42.28084, 42.27219, 42.26332, 42.25425, 42.24495, 
    42.23543, 42.2257, 42.21576, 42.20559, 42.19521, 42.18462, 42.17381, 
    42.16278, 42.15154, 42.14008, 42.12841, 42.11652, 42.10442, 42.09211, 
    42.07958, 42.06683, 42.05388, 42.04071, 42.02732, 42.01372, 41.99991, 
    41.98589, 41.97165, 41.9572, 41.94253, 41.92766, 41.91257, 41.89727, 
    41.88176, 41.86604, 41.8501, 41.83396, 41.8176, 41.80104, 41.78426, 
    41.76727, 41.75008, 41.73267, 41.71505, 41.69723, 41.6792, 41.66095, 
    41.6425, 41.62384, 41.60497, 41.5859, 41.56662, 41.54713, 41.52743, 
    41.50753, 41.48742, 41.4671, 41.44658, 41.42585, 41.40491, 41.38378, 
    41.36243, 41.34089, 41.31913, 41.29718, 41.27502, 41.25266, 41.23009, 
    41.20732, 41.18435, 41.16117, 41.13779, 41.11422, 41.09044, 41.06646, 
    41.04227, 41.01789, 40.99331, 40.96853, 40.94355, 40.91837, 40.89299, 
    40.86741, 40.84164, 40.81566, 40.78949, 40.76312, 40.73655, 40.70979, 
    40.68283, 40.65568, 40.62833, 40.60078, 40.57304, 40.5451, 40.51697, 
    40.48865, 40.46013, 40.43142, 40.40252, 40.37342, 40.34413, 40.31465, 
    40.28498, 40.25512, 40.22506, 40.19481, 40.16438, 40.13375, 40.10294, 
    40.07194, 40.04074, 40.00937, 39.9778, 39.94604, 39.9141, 39.88197, 
    39.84966, 39.81715, 39.78447, 39.75159, 39.71853, 39.68529, 39.65186, 
    39.61825, 39.58446, 39.55048, 39.51632, 39.48198, 39.44746, 39.41275, 
    39.37786, 39.3428,
  35.45267, 35.50283, 35.55285, 35.60271, 35.65244, 35.70203, 35.75147, 
    35.80076, 35.84991, 35.89892, 35.94777, 35.99649, 36.04505, 36.09347, 
    36.14174, 36.18986, 36.23783, 36.28565, 36.33333, 36.38085, 36.42823, 
    36.47545, 36.52252, 36.56944, 36.61621, 36.66282, 36.70929, 36.7556, 
    36.80175, 36.84776, 36.8936, 36.9393, 36.98484, 37.03022, 37.07544, 
    37.12051, 37.16542, 37.21018, 37.25478, 37.29921, 37.34349, 37.38762, 
    37.43158, 37.47538, 37.51902, 37.5625, 37.60582, 37.64898, 37.69197, 
    37.73481, 37.77748, 37.81999, 37.86233, 37.90451, 37.94653, 37.98838, 
    38.03006, 38.07158, 38.11293, 38.15412, 38.19514, 38.23599, 38.27668, 
    38.3172, 38.35754, 38.39772, 38.43773, 38.47757, 38.51724, 38.55674, 
    38.59607, 38.63522, 38.67421, 38.71302, 38.75166, 38.79012, 38.82842, 
    38.86654, 38.90448, 38.94225, 38.97984, 39.01727, 39.05451, 39.09158, 
    39.12846, 39.16518, 39.20171, 39.23807, 39.27425, 39.31025, 39.34607, 
    39.38171, 39.41718, 39.45246, 39.48756, 39.52248, 39.55722, 39.59177, 
    39.62615, 39.66034, 39.69435, 39.72818, 39.76182, 39.79528, 39.82855, 
    39.86164, 39.89454, 39.92726, 39.95979, 39.99214, 40.0243, 40.05627, 
    40.08805, 40.11964, 40.15105, 40.18227, 40.2133, 40.24414, 40.27479, 
    40.30525, 40.33553, 40.3656, 40.39549, 40.42519, 40.45469, 40.484, 
    40.51313, 40.54205, 40.57079, 40.59933, 40.62767, 40.65583, 40.68378, 
    40.71154, 40.73911, 40.76648, 40.79366, 40.82064, 40.84742, 40.874, 
    40.90039, 40.92658, 40.95258, 40.97837, 41.00396, 41.02936, 41.05456, 
    41.07956, 41.10435, 41.12895, 41.15335, 41.17754, 41.20153, 41.22533, 
    41.24892, 41.27231, 41.2955, 41.31848, 41.34126, 41.36384, 41.38622, 
    41.40839, 41.43035, 41.45211, 41.47367, 41.49502, 41.51617, 41.53711, 
    41.55785, 41.57838, 41.5987, 41.61882, 41.63873, 41.65843, 41.67793, 
    41.69721, 41.71629, 41.73516, 41.75383, 41.77228, 41.79053, 41.80856, 
    41.82639, 41.84401, 41.86142, 41.87861, 41.8956, 41.91238, 41.92894, 
    41.9453, 41.96144, 41.97737, 41.99309, 42.0086, 42.0239, 42.03898, 
    42.05385, 42.06851, 42.08295, 42.09719, 42.11121, 42.12502, 42.13861, 
    42.15199, 42.16515, 42.1781, 42.19083, 42.20335, 42.21566, 42.22775, 
    42.23963, 42.25129, 42.26273, 42.27396, 42.28498, 42.29578, 42.30636, 
    42.31672, 42.32687, 42.33681, 42.34652, 42.35602, 42.36531, 42.37437, 
    42.38322, 42.39185, 42.40026, 42.40846, 42.41644, 42.4242, 42.43174, 
    42.43907, 42.44617, 42.45306, 42.45974, 42.46619, 42.47242, 42.47844, 
    42.48423, 42.48981, 42.49517, 42.50031, 42.50523, 42.50993, 42.51442, 
    42.51868, 42.52272, 42.52655, 42.53016, 42.53354, 42.53671, 42.53966, 
    42.54239, 42.5449, 42.54719, 42.54926, 42.55111, 42.55274, 42.55415, 
    42.55534, 42.55631, 42.55706, 42.55759, 42.55791, 42.558, 42.55787, 
    42.55753, 42.55696, 42.55617, 42.55516, 42.55394, 42.55249, 42.55083, 
    42.54894, 42.54684, 42.54451, 42.54197, 42.53921, 42.53622, 42.53302, 
    42.5296, 42.52596, 42.5221, 42.51802, 42.51372, 42.5092, 42.50447, 
    42.49951, 42.49434, 42.48894, 42.48333, 42.4775, 42.47145, 42.46518, 
    42.45869, 42.45199, 42.44506, 42.43792, 42.43056, 42.42299, 42.41519, 
    42.40718, 42.39895, 42.3905, 42.38184, 42.37295, 42.36385, 42.35453, 
    42.345, 42.33525, 42.32528, 42.3151, 42.3047, 42.29408, 42.28325, 
    42.2722, 42.26094, 42.24946, 42.23776, 42.22585, 42.21373, 42.20139, 
    42.18884, 42.17606, 42.16308, 42.14988, 42.13647, 42.12284, 42.109, 
    42.09495, 42.08068, 42.0662, 42.05151, 42.03661, 42.02149, 42.00616, 
    41.99062, 41.97486, 41.9589, 41.94272, 41.92633, 41.90974, 41.89293, 
    41.87591, 41.85868, 41.84124, 41.82359, 41.80573, 41.78765, 41.76937, 
    41.75089, 41.73219, 41.71329, 41.69418, 41.67485, 41.65533, 41.63559, 
    41.61565, 41.5955, 41.57514, 41.55458, 41.53381, 41.51284, 41.49166, 
    41.47028, 41.44868, 41.42689, 41.40489, 41.38269, 41.36028, 41.33767, 
    41.31486, 41.29184, 41.26862, 41.2452, 41.22158, 41.19775, 41.17373, 
    41.1495, 41.12507, 41.10044, 41.07561, 41.05058, 41.02536, 40.99993, 
    40.9743, 40.94847, 40.92245, 40.89623, 40.86981, 40.8432, 40.81638, 
    40.78937, 40.76217, 40.73476, 40.70717, 40.67937, 40.65139, 40.6232, 
    40.59483, 40.56625, 40.53749, 40.50853, 40.47938, 40.45004, 40.42051, 
    40.39078, 40.36086, 40.33075, 40.30045, 40.26996, 40.23928, 40.2084, 
    40.17735, 40.1461, 40.11466, 40.08303, 40.05122, 40.01922, 39.98703, 
    39.95466, 39.9221, 39.88935, 39.85642, 39.8233, 39.79, 39.75651, 
    39.72284, 39.68898, 39.65495, 39.62072, 39.58632, 39.55173, 39.51697, 
    39.48202, 39.44689,
  35.55025, 35.60048, 35.65057, 35.70052, 35.75032, 35.79998, 35.84949, 
    35.89886, 35.94809, 35.99717, 36.0461, 36.09488, 36.14352, 36.19201, 
    36.24036, 36.28855, 36.3366, 36.38449, 36.43224, 36.47984, 36.52729, 
    36.57458, 36.62173, 36.66872, 36.71556, 36.76225, 36.80879, 36.85518, 
    36.9014, 36.94748, 36.9934, 37.03917, 37.08477, 37.13023, 37.17553, 
    37.22067, 37.26565, 37.31048, 37.35515, 37.39966, 37.44401, 37.4882, 
    37.53223, 37.57611, 37.61982, 37.66337, 37.70676, 37.74999, 37.79306, 
    37.83596, 37.8787, 37.92128, 37.9637, 38.00594, 38.04803, 38.08995, 
    38.1317, 38.17329, 38.21471, 38.25597, 38.29706, 38.33798, 38.37873, 
    38.41932, 38.45973, 38.49998, 38.54006, 38.57996, 38.6197, 38.65927, 
    38.69866, 38.73788, 38.77694, 38.81581, 38.85452, 38.89305, 38.93141, 
    38.9696, 39.00761, 39.04544, 39.0831, 39.12059, 39.15789, 39.19503, 
    39.23198, 39.26876, 39.30536, 39.34178, 39.37802, 39.41409, 39.44997, 
    39.48568, 39.5212, 39.55655, 39.59171, 39.62669, 39.66149, 39.69611, 
    39.73055, 39.7648, 39.79887, 39.83276, 39.86646, 39.89997, 39.93331, 
    39.96646, 39.99942, 40.0322, 40.06479, 40.09719, 40.12941, 40.16144, 
    40.19328, 40.22493, 40.2564, 40.28767, 40.31876, 40.34966, 40.38036, 
    40.41088, 40.44121, 40.47134, 40.50129, 40.53104, 40.5606, 40.58997, 
    40.61914, 40.64812, 40.67691, 40.7055, 40.7339, 40.7621, 40.79012, 
    40.81793, 40.84555, 40.87297, 40.9002, 40.92723, 40.95406, 40.98069, 
    41.00713, 41.03337, 41.05941, 41.08526, 41.1109, 41.13634, 41.16159, 
    41.18663, 41.21148, 41.23612, 41.26057, 41.28481, 41.30885, 41.33269, 
    41.35632, 41.37976, 41.40299, 41.42602, 41.44884, 41.47147, 41.49389, 
    41.5161, 41.53811, 41.55991, 41.58151, 41.60291, 41.62409, 41.64507, 
    41.66585, 41.68642, 41.70678, 41.72694, 41.74689, 41.76663, 41.78616, 
    41.80549, 41.8246, 41.84351, 41.86221, 41.88071, 41.89899, 41.91706, 
    41.93492, 41.95257, 41.97002, 41.98725, 42.00427, 42.02108, 42.03767, 
    42.05406, 42.07024, 42.0862, 42.10195, 42.11749, 42.13282, 42.14793, 
    42.16283, 42.17752, 42.192, 42.20626, 42.22031, 42.23414, 42.24776, 
    42.26116, 42.27435, 42.28733, 42.30009, 42.31264, 42.32497, 42.33708, 
    42.34898, 42.36067, 42.37214, 42.38339, 42.39442, 42.40524, 42.41585, 
    42.42624, 42.43641, 42.44636, 42.45609, 42.46561, 42.47491, 42.484, 
    42.49286, 42.50151, 42.50994, 42.51816, 42.52615, 42.53393, 42.54148, 
    42.54882, 42.55595, 42.56285, 42.56953, 42.576, 42.58224, 42.58827, 
    42.59408, 42.59967, 42.60504, 42.61019, 42.61512, 42.61983, 42.62433, 
    42.6286, 42.63265, 42.63649, 42.6401, 42.64349, 42.64667, 42.64962, 
    42.65236, 42.65487, 42.65717, 42.65924, 42.66109, 42.66273, 42.66414, 
    42.66533, 42.66631, 42.66706, 42.66759, 42.66791, 42.668, 42.66787, 
    42.66752, 42.66696, 42.66617, 42.66516, 42.66393, 42.66248, 42.66081, 
    42.65892, 42.65681, 42.65449, 42.65194, 42.64917, 42.64618, 42.64297, 
    42.63954, 42.63589, 42.63203, 42.62794, 42.62363, 42.6191, 42.61436, 
    42.60939, 42.60421, 42.5988, 42.59318, 42.58733, 42.58127, 42.57499, 
    42.56849, 42.56177, 42.55484, 42.54768, 42.54031, 42.53271, 42.5249, 
    42.51687, 42.50863, 42.50016, 42.49147, 42.48257, 42.47346, 42.46412, 
    42.45457, 42.4448, 42.43481, 42.42461, 42.41418, 42.40355, 42.39269, 
    42.38162, 42.37033, 42.35883, 42.34711, 42.33518, 42.32303, 42.31067, 
    42.29808, 42.28529, 42.27228, 42.25906, 42.24562, 42.23196, 42.2181, 
    42.20402, 42.18972, 42.17521, 42.16049, 42.14556, 42.13041, 42.11505, 
    42.09948, 42.08369, 42.06769, 42.05148, 42.03506, 42.01843, 42.00159, 
    41.98454, 41.96727, 41.94979, 41.93211, 41.91422, 41.89611, 41.87779, 
    41.85927, 41.84054, 41.82159, 41.80244, 41.78309, 41.76352, 41.74375, 
    41.72377, 41.70358, 41.68318, 41.66258, 41.64177, 41.62075, 41.59953, 
    41.57811, 41.55648, 41.53464, 41.5126, 41.49035, 41.4679, 41.44525, 
    41.42239, 41.39933, 41.37606, 41.3526, 41.32893, 41.30506, 41.28099, 
    41.25671, 41.23224, 41.20756, 41.18269, 41.15761, 41.13233, 41.10686, 
    41.08118, 41.05531, 41.02924, 41.00296, 40.97649, 40.94983, 40.92297, 
    40.8959, 40.86864, 40.84119, 40.81354, 40.7857, 40.75766, 40.72942, 
    40.70099, 40.67237, 40.64355, 40.61454, 40.58533, 40.55593, 40.52634, 
    40.49656, 40.46659, 40.43642, 40.40607, 40.37552, 40.34478, 40.31386, 
    40.28274, 40.25143, 40.21994, 40.18826, 40.15638, 40.12432, 40.09208, 
    40.05965, 40.02703, 39.99422, 39.96123, 39.92805, 39.89469, 39.86114, 
    39.82741, 39.79349, 39.75939, 39.72511, 39.69065, 39.656, 39.62117, 
    39.58616, 39.55096,
  35.6478, 35.6981, 35.74827, 35.79829, 35.84817, 35.8979, 35.94749, 
    35.99693, 36.04623, 36.09539, 36.14439, 36.19325, 36.24197, 36.29053, 
    36.33895, 36.38722, 36.43534, 36.48331, 36.53113, 36.5788, 36.62632, 
    36.67369, 36.72091, 36.76798, 36.81489, 36.86166, 36.90826, 36.95472, 
    37.00102, 37.04717, 37.09316, 37.139, 37.18468, 37.23021, 37.27558, 
    37.3208, 37.36585, 37.41075, 37.45549, 37.50007, 37.5445, 37.58876, 
    37.63287, 37.67681, 37.72059, 37.76422, 37.80768, 37.85098, 37.89412, 
    37.93709, 37.9799, 38.02255, 38.06503, 38.10735, 38.14951, 38.1915, 
    38.23332, 38.27498, 38.31647, 38.3578, 38.39895, 38.43994, 38.48076, 
    38.52142, 38.5619, 38.60221, 38.64236, 38.68233, 38.72214, 38.76178, 
    38.80124, 38.84053, 38.87964, 38.91859, 38.95736, 38.99596, 39.03439, 
    39.07264, 39.11071, 39.14861, 39.18634, 39.22389, 39.26126, 39.29846, 
    39.33548, 39.37232, 39.40898, 39.44547, 39.48177, 39.5179, 39.55385, 
    39.58962, 39.62521, 39.66061, 39.69584, 39.73088, 39.76575, 39.80043, 
    39.83492, 39.86924, 39.90337, 39.93732, 39.97108, 40.00466, 40.03805, 
    40.07126, 40.10428, 40.13712, 40.16977, 40.20223, 40.23451, 40.26659, 
    40.2985, 40.33021, 40.36173, 40.39306, 40.42421, 40.45516, 40.48592, 
    40.51649, 40.54688, 40.57707, 40.60707, 40.63688, 40.66649, 40.69591, 
    40.72514, 40.75417, 40.78302, 40.81166, 40.84011, 40.86837, 40.89643, 
    40.9243, 40.95197, 40.97945, 41.00673, 41.03381, 41.06069, 41.08738, 
    41.11386, 41.14015, 41.16624, 41.19213, 41.21783, 41.24332, 41.26861, 
    41.2937, 41.3186, 41.34329, 41.36778, 41.39207, 41.41615, 41.44004, 
    41.46372, 41.4872, 41.51048, 41.53355, 41.55642, 41.57909, 41.60155, 
    41.6238, 41.64585, 41.6677, 41.68934, 41.71078, 41.73201, 41.75303, 
    41.77385, 41.79446, 41.81486, 41.83506, 41.85505, 41.87482, 41.89439, 
    41.91376, 41.93291, 41.95186, 41.9706, 41.98912, 42.00744, 42.02555, 
    42.04345, 42.06113, 42.07861, 42.09587, 42.11293, 42.12977, 42.1464, 
    42.16282, 42.17903, 42.19503, 42.21081, 42.22638, 42.24174, 42.25688, 
    42.27181, 42.28653, 42.30103, 42.31532, 42.3294, 42.34326, 42.35691, 
    42.37034, 42.38356, 42.39656, 42.40934, 42.42192, 42.43427, 42.44641, 
    42.45834, 42.47004, 42.48153, 42.49281, 42.50387, 42.51471, 42.52533, 
    42.53574, 42.54593, 42.5559, 42.56566, 42.5752, 42.58452, 42.59362, 
    42.60251, 42.61117, 42.61962, 42.62785, 42.63586, 42.64365, 42.65123, 
    42.65858, 42.66572, 42.67263, 42.67933, 42.68581, 42.69207, 42.69811, 
    42.70393, 42.70953, 42.71491, 42.72007, 42.72501, 42.72974, 42.73424, 
    42.73852, 42.74258, 42.74642, 42.75004, 42.75344, 42.75663, 42.75959, 
    42.76233, 42.76484, 42.76714, 42.76922, 42.77108, 42.77272, 42.77413, 
    42.77533, 42.7763, 42.77706, 42.77759, 42.77791, 42.778, 42.77787, 
    42.77752, 42.77695, 42.77617, 42.77515, 42.77392, 42.77247, 42.7708, 
    42.76891, 42.76679, 42.76446, 42.76191, 42.75913, 42.75613, 42.75292, 
    42.74949, 42.74583, 42.74195, 42.73786, 42.73354, 42.729, 42.72425, 
    42.71927, 42.71408, 42.70866, 42.70303, 42.69717, 42.6911, 42.6848, 
    42.67829, 42.67155, 42.6646, 42.65743, 42.65004, 42.64244, 42.63461, 
    42.62656, 42.6183, 42.60982, 42.60112, 42.5922, 42.58306, 42.5737, 
    42.56413, 42.55434, 42.54433, 42.53411, 42.52367, 42.51301, 42.50213, 
    42.49104, 42.47973, 42.4682, 42.45646, 42.4445, 42.43233, 42.41994, 
    42.40734, 42.39452, 42.38148, 42.36823, 42.35476, 42.34108, 42.32719, 
    42.31308, 42.29875, 42.28421, 42.26947, 42.2545, 42.23932, 42.22393, 
    42.20833, 42.19251, 42.17648, 42.16024, 42.14379, 42.12712, 42.11024, 
    42.09316, 42.07586, 42.05835, 42.04063, 42.0227, 42.00456, 41.98621, 
    41.96765, 41.94888, 41.9299, 41.91071, 41.89131, 41.87171, 41.85189, 
    41.83187, 41.81165, 41.79121, 41.77057, 41.74972, 41.72866, 41.7074, 
    41.68593, 41.66426, 41.64238, 41.6203, 41.59801, 41.57551, 41.55281, 
    41.52991, 41.50681, 41.4835, 41.45999, 41.43628, 41.41236, 41.38824, 
    41.36392, 41.3394, 41.31467, 41.28975, 41.26463, 41.2393, 41.21378, 
    41.18805, 41.16213, 41.13601, 41.10968, 41.08316, 41.05645, 41.02953, 
    41.00242, 40.97511, 40.94761, 40.91991, 40.89201, 40.86391, 40.83563, 
    40.80714, 40.77847, 40.7496, 40.72053, 40.69127, 40.66182, 40.63217, 
    40.60234, 40.57231, 40.54208, 40.51167, 40.48107, 40.45028, 40.41929, 
    40.38812, 40.35675, 40.3252, 40.29346, 40.26153, 40.22942, 40.19711, 
    40.16462, 40.13194, 40.09907, 40.06602, 40.03278, 39.99936, 39.96575, 
    39.93196, 39.89798, 39.86382, 39.82948, 39.79495, 39.76024, 39.72535, 
    39.69028, 39.65503,
  35.74531, 35.79569, 35.84593, 35.89603, 35.94598, 35.99579, 36.04546, 
    36.09497, 36.14435, 36.19357, 36.24266, 36.29159, 36.34038, 36.38902, 
    36.43751, 36.48585, 36.53405, 36.58209, 36.62999, 36.67773, 36.72533, 
    36.77277, 36.82006, 36.8672, 36.91419, 36.96103, 37.00771, 37.05424, 
    37.10061, 37.14684, 37.1929, 37.23881, 37.28457, 37.33017, 37.37561, 
    37.42089, 37.46603, 37.51099, 37.55581, 37.60046, 37.64496, 37.68929, 
    37.73347, 37.77748, 37.82134, 37.86504, 37.90857, 37.95194, 37.99514, 
    38.03819, 38.08107, 38.12379, 38.16634, 38.20873, 38.25096, 38.29302, 
    38.33491, 38.37664, 38.4182, 38.45959, 38.50082, 38.54188, 38.58277, 
    38.62349, 38.66405, 38.70443, 38.74464, 38.78469, 38.82456, 38.86426, 
    38.90379, 38.94315, 38.98233, 39.02134, 39.06018, 39.09885, 39.13734, 
    39.17566, 39.21379, 39.25176, 39.28955, 39.32717, 39.36461, 39.40187, 
    39.43895, 39.47586, 39.51259, 39.54914, 39.58551, 39.6217, 39.65771, 
    39.69354, 39.72919, 39.76466, 39.79995, 39.83506, 39.86998, 39.90472, 
    39.93929, 39.97366, 40.00785, 40.04186, 40.07569, 40.10933, 40.14278, 
    40.17605, 40.20913, 40.24202, 40.27473, 40.30725, 40.33959, 40.37173, 
    40.40369, 40.43546, 40.46704, 40.49844, 40.52964, 40.56065, 40.59147, 
    40.6221, 40.65253, 40.68278, 40.71284, 40.7427, 40.77237, 40.80185, 
    40.83113, 40.86022, 40.88911, 40.91781, 40.94632, 40.97463, 41.00274, 
    41.03066, 41.05838, 41.08591, 41.11324, 41.14037, 41.1673, 41.19404, 
    41.22058, 41.24692, 41.27306, 41.299, 41.32474, 41.35028, 41.37563, 
    41.40077, 41.4257, 41.45045, 41.47498, 41.49932, 41.52345, 41.54738, 
    41.57111, 41.59464, 41.61795, 41.64107, 41.66399, 41.6867, 41.7092, 
    41.7315, 41.75359, 41.77548, 41.79717, 41.81865, 41.83992, 41.86098, 
    41.88184, 41.90249, 41.92293, 41.94316, 41.96319, 41.98301, 42.00262, 
    42.02202, 42.04121, 42.0602, 42.07897, 42.09754, 42.11589, 42.13403, 
    42.15197, 42.16969, 42.1872, 42.2045, 42.22159, 42.23846, 42.25513, 
    42.27158, 42.28782, 42.30385, 42.31966, 42.33526, 42.35065, 42.36583, 
    42.38079, 42.39553, 42.41007, 42.42439, 42.43849, 42.45238, 42.46605, 
    42.47951, 42.49276, 42.50578, 42.5186, 42.53119, 42.54357, 42.55574, 
    42.56768, 42.57942, 42.59093, 42.60223, 42.61331, 42.62417, 42.63482, 
    42.64525, 42.65546, 42.66545, 42.67523, 42.68479, 42.69413, 42.70325, 
    42.71215, 42.72083, 42.7293, 42.73755, 42.74557, 42.75338, 42.76097, 
    42.76834, 42.77549, 42.78242, 42.78913, 42.79562, 42.8019, 42.80795, 
    42.81378, 42.81939, 42.82478, 42.82996, 42.83491, 42.83964, 42.84415, 
    42.84844, 42.85251, 42.85636, 42.85999, 42.86339, 42.86658, 42.86954, 
    42.87229, 42.87482, 42.87712, 42.8792, 42.88107, 42.88271, 42.88412, 
    42.88532, 42.8863, 42.88706, 42.88759, 42.88791, 42.888, 42.88787, 
    42.88752, 42.88695, 42.88616, 42.88515, 42.88391, 42.88246, 42.88078, 
    42.87889, 42.87677, 42.87443, 42.87187, 42.86909, 42.86609, 42.86287, 
    42.85943, 42.85576, 42.85188, 42.84777, 42.84345, 42.83891, 42.83414, 
    42.82915, 42.82394, 42.81852, 42.81287, 42.807, 42.80092, 42.79461, 
    42.78809, 42.78134, 42.77437, 42.76719, 42.75978, 42.75216, 42.74432, 
    42.73626, 42.72797, 42.71947, 42.71075, 42.70182, 42.69266, 42.68329, 
    42.6737, 42.66389, 42.65386, 42.64361, 42.63315, 42.62247, 42.61157, 
    42.60046, 42.58912, 42.57758, 42.56581, 42.55383, 42.54163, 42.52921, 
    42.51658, 42.50373, 42.49067, 42.4774, 42.4639, 42.4502, 42.43627, 
    42.42213, 42.40778, 42.39322, 42.37843, 42.36344, 42.34823, 42.33281, 
    42.31718, 42.30133, 42.28527, 42.26899, 42.25251, 42.23581, 42.2189, 
    42.20178, 42.18444, 42.1669, 42.14914, 42.13118, 42.113, 42.09461, 
    42.07602, 42.05721, 42.03819, 42.01897, 41.99953, 41.97989, 41.96004, 
    41.93998, 41.91971, 41.89923, 41.87855, 41.85766, 41.83656, 41.81526, 
    41.79375, 41.77203, 41.75011, 41.72799, 41.70565, 41.68312, 41.66037, 
    41.63743, 41.61428, 41.59093, 41.56737, 41.54361, 41.51965, 41.49548, 
    41.47112, 41.44654, 41.42178, 41.3968, 41.37163, 41.34626, 41.32068, 
    41.29491, 41.26894, 41.24277, 41.2164, 41.18983, 41.16306, 41.13609, 
    41.10893, 41.08157, 41.05401, 41.02626, 40.99831, 40.97016, 40.94182, 
    40.91328, 40.88455, 40.85563, 40.82651, 40.7972, 40.76769, 40.73799, 
    40.7081, 40.67801, 40.64773, 40.61726, 40.58661, 40.55576, 40.52471, 
    40.49348, 40.46206, 40.43045, 40.39865, 40.36666, 40.33449, 40.30212, 
    40.26957, 40.23684, 40.20391, 40.1708, 40.1375, 40.10402, 40.07035, 
    40.0365, 40.00246, 39.96824, 39.93383, 39.89924, 39.86447, 39.82952, 
    39.79438, 39.75906,
  35.84279, 35.89325, 35.94357, 35.99374, 36.04376, 36.09365, 36.14339, 
    36.19298, 36.24243, 36.29173, 36.34089, 36.3899, 36.43876, 36.48747, 
    36.53604, 36.58445, 36.63272, 36.68084, 36.72881, 36.77663, 36.8243, 
    36.87182, 36.91919, 36.9664, 37.01346, 37.06037, 37.10712, 37.15373, 
    37.20018, 37.24647, 37.29261, 37.3386, 37.38442, 37.4301, 37.47561, 
    37.52097, 37.56617, 37.61121, 37.6561, 37.70082, 37.74539, 37.7898, 
    37.83405, 37.87814, 37.92206, 37.96582, 38.00943, 38.05287, 38.09615, 
    38.13927, 38.18222, 38.22501, 38.26763, 38.31009, 38.35239, 38.39452, 
    38.43648, 38.47828, 38.51991, 38.56137, 38.60267, 38.6438, 38.68475, 
    38.72554, 38.76617, 38.80662, 38.8469, 38.88701, 38.92695, 38.96672, 
    39.00632, 39.04574, 39.085, 39.12407, 39.16298, 39.20171, 39.24027, 
    39.27865, 39.31686, 39.35489, 39.39275, 39.43043, 39.46793, 39.50526, 
    39.54241, 39.57938, 39.61617, 39.65279, 39.68922, 39.72548, 39.76155, 
    39.79745, 39.83316, 39.86869, 39.90405, 39.93922, 39.9742, 40.00901, 
    40.04363, 40.07807, 40.11232, 40.14639, 40.18027, 40.21397, 40.24749, 
    40.28082, 40.31396, 40.34691, 40.37968, 40.41226, 40.44466, 40.47686, 
    40.50888, 40.54071, 40.57235, 40.60379, 40.63505, 40.66612, 40.69699, 
    40.72768, 40.75818, 40.78848, 40.81859, 40.84851, 40.87823, 40.90776, 
    40.9371, 40.96624, 40.99519, 41.02395, 41.05251, 41.08087, 41.10904, 
    41.13701, 41.16478, 41.19236, 41.21975, 41.24693, 41.27391, 41.3007, 
    41.32729, 41.35368, 41.37987, 41.40586, 41.43165, 41.45724, 41.48263, 
    41.50782, 41.53281, 41.55759, 41.58218, 41.60656, 41.63074, 41.65471, 
    41.67849, 41.70206, 41.72543, 41.74859, 41.77155, 41.7943, 41.81684, 
    41.83919, 41.86133, 41.88326, 41.90498, 41.9265, 41.94781, 41.96892, 
    41.98982, 42.01051, 42.03099, 42.05127, 42.07133, 42.09119, 42.11084, 
    42.13028, 42.14951, 42.16853, 42.18734, 42.20594, 42.22433, 42.24251, 
    42.26048, 42.27824, 42.29578, 42.31312, 42.33024, 42.34715, 42.36385, 
    42.38033, 42.39661, 42.41267, 42.42851, 42.44415, 42.45956, 42.47477, 
    42.48976, 42.50454, 42.5191, 42.53344, 42.54758, 42.56149, 42.5752, 
    42.58868, 42.60195, 42.61501, 42.62784, 42.64046, 42.65287, 42.66506, 
    42.67703, 42.68879, 42.70033, 42.71165, 42.72275, 42.73363, 42.7443, 
    42.75475, 42.76498, 42.775, 42.78479, 42.79437, 42.80373, 42.81287, 
    42.82179, 42.83049, 42.83897, 42.84724, 42.85528, 42.86311, 42.87071, 
    42.87809, 42.88526, 42.8922, 42.89893, 42.90543, 42.91172, 42.91778, 
    42.92363, 42.92925, 42.93465, 42.93983, 42.9448, 42.94954, 42.95406, 
    42.95836, 42.96244, 42.96629, 42.96993, 42.97334, 42.97654, 42.97951, 
    42.98226, 42.98479, 42.9871, 42.98919, 42.99105, 42.99269, 42.99412, 
    42.99532, 42.9963, 42.99706, 42.99759, 42.99791, 42.998, 42.99787, 
    42.99752, 42.99695, 42.99616, 42.99514, 42.99391, 42.99245, 42.99077, 
    42.98887, 42.98675, 42.98441, 42.98184, 42.97905, 42.97605, 42.97282, 
    42.96937, 42.9657, 42.9618, 42.95769, 42.95336, 42.9488, 42.94403, 
    42.93903, 42.93382, 42.92838, 42.92272, 42.91684, 42.91074, 42.90442, 
    42.89788, 42.89112, 42.88414, 42.87694, 42.86952, 42.86188, 42.85402, 
    42.84594, 42.83765, 42.82913, 42.82039, 42.81144, 42.80227, 42.79287, 
    42.78326, 42.77343, 42.76338, 42.75312, 42.74263, 42.73193, 42.72101, 
    42.70987, 42.69852, 42.68694, 42.67515, 42.66315, 42.65092, 42.63848, 
    42.62583, 42.61295, 42.59986, 42.58656, 42.57304, 42.55931, 42.54536, 
    42.53119, 42.51681, 42.50221, 42.4874, 42.47238, 42.45714, 42.44168, 
    42.42602, 42.41014, 42.39405, 42.37774, 42.36122, 42.34449, 42.32755, 
    42.31039, 42.29302, 42.27544, 42.25765, 42.23965, 42.22144, 42.20301, 
    42.18438, 42.16554, 42.14648, 42.12722, 42.10775, 42.08807, 42.06818, 
    42.04808, 42.02777, 42.00725, 41.98653, 41.9656, 41.94446, 41.92311, 
    41.90156, 41.8798, 41.85784, 41.83567, 41.81329, 41.79071, 41.76793, 
    41.74494, 41.72174, 41.69834, 41.67474, 41.65094, 41.62693, 41.60271, 
    41.5783, 41.55368, 41.52887, 41.50385, 41.47863, 41.45321, 41.42758, 
    41.40176, 41.37574, 41.34952, 41.32309, 41.29647, 41.26966, 41.24264, 
    41.21543, 41.18801, 41.1604, 41.1326, 41.1046, 41.0764, 41.048, 41.01941, 
    40.99063, 40.96165, 40.93247, 40.90311, 40.87354, 40.84379, 40.81384, 
    40.7837, 40.75336, 40.72284, 40.69212, 40.66122, 40.63012, 40.59883, 
    40.56735, 40.53568, 40.50383, 40.47178, 40.43954, 40.40712, 40.37451, 
    40.34171, 40.30873, 40.27556, 40.2422, 40.20866, 40.17493, 40.14101, 
    40.10691, 40.07263, 40.03816, 40.00351, 39.96868, 39.93366, 39.89846, 
    39.86309,
  35.94024, 35.99077, 36.04116, 36.09141, 36.14151, 36.19147, 36.24129, 
    36.29095, 36.34048, 36.38985, 36.43909, 36.48817, 36.53711, 36.5859, 
    36.63454, 36.68303, 36.73137, 36.77956, 36.82761, 36.8755, 36.92324, 
    36.97084, 37.01828, 37.06556, 37.1127, 37.15968, 37.20651, 37.25319, 
    37.29971, 37.34608, 37.39229, 37.43835, 37.48425, 37.52999, 37.57558, 
    37.62101, 37.66629, 37.7114, 37.75636, 37.80116, 37.8458, 37.89028, 
    37.9346, 37.97876, 38.02275, 38.06659, 38.11027, 38.15378, 38.19713, 
    38.24031, 38.28334, 38.3262, 38.36889, 38.41143, 38.45379, 38.49599, 
    38.53802, 38.57989, 38.62159, 38.66312, 38.70449, 38.74569, 38.78672, 
    38.82758, 38.86826, 38.90878, 38.94913, 38.98932, 39.02932, 39.06916, 
    39.10883, 39.14832, 39.18764, 39.22678, 39.26575, 39.30455, 39.34318, 
    39.38163, 39.4199, 39.458, 39.49592, 39.53367, 39.57124, 39.60863, 
    39.64584, 39.68288, 39.71974, 39.75642, 39.79292, 39.82924, 39.86538, 
    39.90133, 39.93711, 39.97271, 40.00812, 40.04335, 40.0784, 40.11327, 
    40.14795, 40.18245, 40.21677, 40.2509, 40.28485, 40.31861, 40.35218, 
    40.38557, 40.41877, 40.45179, 40.48462, 40.51726, 40.54971, 40.58197, 
    40.61405, 40.64593, 40.67763, 40.70914, 40.74045, 40.77158, 40.80251, 
    40.83326, 40.8638, 40.89417, 40.92433, 40.9543, 40.98409, 41.01367, 
    41.04306, 41.07226, 41.10126, 41.13007, 41.15868, 41.1871, 41.21532, 
    41.24335, 41.27118, 41.29881, 41.32624, 41.35347, 41.38051, 41.40734, 
    41.43398, 41.46042, 41.48666, 41.5127, 41.53854, 41.56418, 41.58962, 
    41.61486, 41.6399, 41.66473, 41.68936, 41.71379, 41.73801, 41.76204, 
    41.78586, 41.80947, 41.83289, 41.85609, 41.87909, 41.90189, 41.92448, 
    41.94687, 41.96905, 41.99103, 42.01279, 42.03436, 42.05571, 42.07686, 
    42.0978, 42.11853, 42.13905, 42.15937, 42.17947, 42.19937, 42.21906, 
    42.23853, 42.2578, 42.27686, 42.29571, 42.31435, 42.33277, 42.35099, 
    42.36899, 42.38678, 42.40437, 42.42173, 42.43889, 42.45583, 42.47256, 
    42.48908, 42.50539, 42.52148, 42.53736, 42.55302, 42.56847, 42.58371, 
    42.59873, 42.61353, 42.62812, 42.6425, 42.65666, 42.6706, 42.68433, 
    42.69785, 42.71114, 42.72422, 42.73709, 42.74974, 42.76217, 42.77438, 
    42.78638, 42.79816, 42.80972, 42.82106, 42.83219, 42.84309, 42.85379, 
    42.86426, 42.87451, 42.88454, 42.89436, 42.90395, 42.91333, 42.92249, 
    42.93143, 42.94015, 42.94865, 42.95693, 42.96499, 42.97283, 42.98045, 
    42.98785, 42.99503, 43.00199, 43.00873, 43.01524, 43.02154, 43.02762, 
    43.03347, 43.03911, 43.04453, 43.04972, 43.05469, 43.05944, 43.06397, 
    43.06828, 43.07236, 43.07623, 43.07987, 43.08329, 43.08649, 43.08947, 
    43.09223, 43.09476, 43.09708, 43.09917, 43.10104, 43.10268, 43.10411, 
    43.10531, 43.10629, 43.10705, 43.10759, 43.10791, 43.108, 43.10787, 
    43.10752, 43.10695, 43.10615, 43.10514, 43.1039, 43.10244, 43.10075, 
    43.09885, 43.09673, 43.09438, 43.0918, 43.08902, 43.086, 43.08277, 
    43.07931, 43.07563, 43.07173, 43.06761, 43.06327, 43.0587, 43.05392, 
    43.04891, 43.04368, 43.03823, 43.03256, 43.02667, 43.02056, 43.01423, 
    43.00768, 43.0009, 42.99391, 42.98669, 42.97926, 42.9716, 42.96373, 
    42.95563, 42.94732, 42.93878, 42.93003, 42.92105, 42.91186, 42.90245, 
    42.89282, 42.88297, 42.8729, 42.86261, 42.85211, 42.84138, 42.83044, 
    42.81928, 42.8079, 42.79631, 42.7845, 42.77246, 42.76022, 42.74775, 
    42.73507, 42.72217, 42.70906, 42.69572, 42.68218, 42.66842, 42.65443, 
    42.64024, 42.62583, 42.61121, 42.59636, 42.58131, 42.56604, 42.55056, 
    42.53486, 42.51895, 42.50282, 42.48648, 42.46993, 42.45317, 42.43619, 
    42.419, 42.4016, 42.38398, 42.36616, 42.34812, 42.32987, 42.31141, 
    42.29274, 42.27386, 42.25477, 42.23547, 42.21595, 42.19624, 42.1763, 
    42.15617, 42.13582, 42.11526, 42.0945, 42.07352, 42.05235, 42.03096, 
    42.00937, 41.98756, 41.96556, 41.94334, 41.92093, 41.8983, 41.87547, 
    41.85244, 41.8292, 41.80575, 41.7821, 41.75825, 41.7342, 41.70994, 
    41.68548, 41.66081, 41.63595, 41.61088, 41.58561, 41.56014, 41.53447, 
    41.5086, 41.48253, 41.45626, 41.42978, 41.40311, 41.37624, 41.34917, 
    41.32191, 41.29445, 41.26678, 41.23893, 41.21087, 41.18262, 41.15417, 
    41.12553, 41.09669, 41.06765, 41.03843, 41.009, 40.97939, 40.94957, 
    40.91957, 40.88937, 40.85899, 40.8284, 40.79763, 40.76667, 40.73551, 
    40.70417, 40.67263, 40.6409, 40.60899, 40.57688, 40.54459, 40.5121, 
    40.47943, 40.44658, 40.41353, 40.3803, 40.34688, 40.31328, 40.27949, 
    40.24551, 40.21135, 40.17701, 40.14248, 40.10777, 40.07287, 40.03779, 
    40.00253, 39.96709,
  36.03765, 36.08826, 36.13873, 36.18905, 36.23923, 36.28926, 36.33915, 
    36.3889, 36.4385, 36.48795, 36.53725, 36.58641, 36.63543, 36.68429, 
    36.733, 36.78157, 36.82999, 36.87825, 36.92637, 36.97434, 37.02216, 
    37.06982, 37.11734, 37.1647, 37.21191, 37.25897, 37.30587, 37.35262, 
    37.39922, 37.44566, 37.49194, 37.53807, 37.58405, 37.62986, 37.67553, 
    37.72103, 37.76638, 37.81157, 37.85659, 37.90147, 37.94618, 37.99073, 
    38.03512, 38.07935, 38.12342, 38.16733, 38.21107, 38.25466, 38.29808, 
    38.34134, 38.38443, 38.42736, 38.47013, 38.51273, 38.55517, 38.59744, 
    38.63954, 38.68148, 38.72325, 38.76485, 38.80629, 38.84755, 38.88865, 
    38.92958, 38.97034, 39.01093, 39.05135, 39.09159, 39.13167, 39.17157, 
    39.21131, 39.25087, 39.29026, 39.32947, 39.36851, 39.40738, 39.44607, 
    39.48458, 39.52292, 39.56109, 39.59908, 39.63689, 39.67452, 39.71198, 
    39.74926, 39.78636, 39.82328, 39.86003, 39.89659, 39.93298, 39.96918, 
    40.0052, 40.04104, 40.0767, 40.11218, 40.14747, 40.18259, 40.21751, 
    40.25226, 40.28682, 40.3212, 40.35539, 40.3894, 40.42322, 40.45686, 
    40.49031, 40.52357, 40.55664, 40.58953, 40.62223, 40.65474, 40.68707, 
    40.7192, 40.75114, 40.7829, 40.81446, 40.84584, 40.87702, 40.90801, 
    40.93881, 40.96942, 40.99984, 41.03006, 41.06009, 41.08992, 41.11956, 
    41.14901, 41.17826, 41.20732, 41.23618, 41.26485, 41.29332, 41.32159, 
    41.34967, 41.37755, 41.40523, 41.43272, 41.46, 41.48709, 41.51398, 
    41.54067, 41.56716, 41.59345, 41.61954, 41.64543, 41.67112, 41.69661, 
    41.72189, 41.74697, 41.77185, 41.79654, 41.82101, 41.84528, 41.86935, 
    41.89322, 41.91688, 41.94034, 41.96359, 41.98664, 42.00948, 42.03212, 
    42.05455, 42.07677, 42.09879, 42.1206, 42.1422, 42.1636, 42.18478, 
    42.20576, 42.22654, 42.2471, 42.26746, 42.2876, 42.30754, 42.32726, 
    42.34678, 42.36609, 42.38518, 42.40407, 42.42274, 42.4412, 42.45946, 
    42.4775, 42.49532, 42.51294, 42.53034, 42.54753, 42.56451, 42.58128, 
    42.59783, 42.61417, 42.63029, 42.6462, 42.66189, 42.67737, 42.69264, 
    42.70769, 42.72253, 42.73715, 42.75155, 42.76574, 42.77971, 42.79347, 
    42.80701, 42.82034, 42.83344, 42.84633, 42.859, 42.87146, 42.8837, 
    42.89572, 42.90752, 42.91911, 42.93048, 42.94162, 42.95255, 42.96326, 
    42.97376, 42.98403, 42.99409, 43.00392, 43.01354, 43.02293, 43.03211, 
    43.04107, 43.0498, 43.05832, 43.06662, 43.0747, 43.08255, 43.09019, 
    43.0976, 43.1048, 43.11177, 43.11852, 43.12505, 43.13136, 43.13745, 
    43.14332, 43.14897, 43.15439, 43.1596, 43.16458, 43.16934, 43.17388, 
    43.1782, 43.18229, 43.18616, 43.18981, 43.19324, 43.19645, 43.19943, 
    43.20219, 43.20473, 43.20705, 43.20915, 43.21102, 43.21267, 43.2141, 
    43.21531, 43.21629, 43.21705, 43.21759, 43.21791, 43.218, 43.21787, 
    43.21752, 43.21695, 43.21615, 43.21513, 43.21389, 43.21243, 43.21074, 
    43.20883, 43.2067, 43.20435, 43.20177, 43.19897, 43.19596, 43.19271, 
    43.18925, 43.18557, 43.18166, 43.17752, 43.17318, 43.1686, 43.16381, 
    43.15879, 43.15355, 43.14809, 43.14241, 43.13651, 43.13038, 43.12403, 
    43.11747, 43.11068, 43.10367, 43.09644, 43.08899, 43.08132, 43.07343, 
    43.06532, 43.05699, 43.04844, 43.03967, 43.03067, 43.02146, 43.01203, 
    43.00238, 42.99251, 42.98242, 42.97211, 42.96159, 42.95084, 42.93988, 
    42.92869, 42.91729, 42.90567, 42.89383, 42.88178, 42.86951, 42.85701, 
    42.84431, 42.83138, 42.81824, 42.80488, 42.79131, 42.77752, 42.76351, 
    42.74929, 42.73485, 42.7202, 42.70533, 42.69024, 42.67494, 42.65942, 
    42.6437, 42.62775, 42.6116, 42.59522, 42.57864, 42.56184, 42.54483, 
    42.52761, 42.51017, 42.49252, 42.47466, 42.45658, 42.4383, 42.4198, 
    42.4011, 42.38218, 42.36305, 42.34371, 42.32416, 42.3044, 42.28443, 
    42.26425, 42.24386, 42.22327, 42.20246, 42.18145, 42.16022, 42.1388, 
    42.11716, 42.09532, 42.07327, 42.05101, 42.02855, 42.00588, 41.98301, 
    41.95993, 41.93664, 41.91315, 41.88946, 41.86556, 41.84146, 41.81715, 
    41.79264, 41.76793, 41.74302, 41.7179, 41.69258, 41.66707, 41.64135, 
    41.61543, 41.58931, 41.56298, 41.53646, 41.50974, 41.48282, 41.4557, 
    41.42838, 41.40087, 41.37315, 41.34524, 41.31713, 41.28883, 41.26033, 
    41.23163, 41.20274, 41.17365, 41.14436, 41.11489, 41.08522, 41.05535, 
    41.02529, 40.99504, 40.96459, 40.93395, 40.90312, 40.8721, 40.84089, 
    40.80948, 40.77789, 40.74611, 40.71413, 40.68196, 40.64961, 40.61707, 
    40.58434, 40.55143, 40.51832, 40.48503, 40.45155, 40.41788, 40.38403, 
    40.34999, 40.31577, 40.28137, 40.24678, 40.212, 40.17704, 40.1419, 
    40.10658, 40.07107,
  36.13504, 36.18572, 36.23626, 36.28666, 36.33691, 36.38702, 36.43699, 
    36.48681, 36.53648, 36.58601, 36.63539, 36.68462, 36.73371, 36.78265, 
    36.83144, 36.88008, 36.92857, 36.97691, 37.02511, 37.07315, 37.12104, 
    37.16878, 37.21637, 37.26381, 37.31109, 37.35822, 37.4052, 37.45202, 
    37.49869, 37.5452, 37.59156, 37.63777, 37.68382, 37.72971, 37.77544, 
    37.82102, 37.86644, 37.9117, 37.9568, 38.00174, 38.04653, 38.09115, 
    38.13562, 38.17992, 38.22406, 38.26804, 38.31186, 38.35551, 38.39901, 
    38.44234, 38.4855, 38.5285, 38.57134, 38.61401, 38.65652, 38.69886, 
    38.74104, 38.78304, 38.82488, 38.86655, 38.90806, 38.94939, 38.99056, 
    39.03156, 39.07239, 39.11305, 39.15353, 39.19385, 39.234, 39.27397, 
    39.31377, 39.3534, 39.39285, 39.43213, 39.47124, 39.51017, 39.54893, 
    39.58752, 39.62592, 39.66415, 39.70221, 39.74009, 39.77779, 39.81531, 
    39.85266, 39.88982, 39.92681, 39.96362, 40.00024, 40.03669, 40.07296, 
    40.10905, 40.14495, 40.18068, 40.21622, 40.25158, 40.28675, 40.32174, 
    40.35655, 40.39117, 40.42561, 40.45987, 40.49393, 40.52782, 40.56152, 
    40.59502, 40.62835, 40.66148, 40.69443, 40.72719, 40.75976, 40.79214, 
    40.82434, 40.85634, 40.88815, 40.91978, 40.95121, 40.98245, 41.0135, 
    41.04435, 41.07502, 41.10549, 41.13577, 41.16586, 41.19574, 41.22544, 
    41.25494, 41.28425, 41.31337, 41.34228, 41.371, 41.39952, 41.42785, 
    41.45598, 41.48391, 41.51165, 41.53918, 41.56652, 41.59366, 41.62061, 
    41.64734, 41.67389, 41.70023, 41.72636, 41.7523, 41.77804, 41.80358, 
    41.82891, 41.85404, 41.87897, 41.9037, 41.92822, 41.95254, 41.97666, 
    42.00057, 42.02428, 42.04778, 42.07108, 42.09417, 42.11706, 42.13974, 
    42.16221, 42.18448, 42.20654, 42.22839, 42.25004, 42.27148, 42.29271, 
    42.31373, 42.33454, 42.35514, 42.37554, 42.39573, 42.4157, 42.43547, 
    42.45502, 42.47437, 42.4935, 42.51242, 42.53113, 42.54963, 42.56792, 
    42.58599, 42.60386, 42.62151, 42.63895, 42.65617, 42.67318, 42.68998, 
    42.70657, 42.72294, 42.73909, 42.75504, 42.77076, 42.78627, 42.80157, 
    42.81665, 42.83152, 42.84617, 42.8606, 42.87482, 42.88882, 42.9026, 
    42.91617, 42.92952, 42.94266, 42.95557, 42.96827, 42.98075, 42.99302, 
    43.00506, 43.01689, 43.0285, 43.03989, 43.05106, 43.06201, 43.07274, 
    43.08326, 43.09355, 43.10363, 43.11348, 43.12312, 43.13253, 43.14173, 
    43.1507, 43.15946, 43.16799, 43.17631, 43.1844, 43.19227, 43.19992, 
    43.20736, 43.21456, 43.22155, 43.22832, 43.23486, 43.24118, 43.24729, 
    43.25317, 43.25883, 43.26426, 43.26948, 43.27447, 43.27924, 43.28379, 
    43.28811, 43.29222, 43.2961, 43.29976, 43.30319, 43.3064, 43.30939, 
    43.31216, 43.31471, 43.31703, 43.31913, 43.32101, 43.32266, 43.32409, 
    43.3253, 43.32629, 43.32705, 43.32759, 43.3279, 43.328, 43.32787, 
    43.32752, 43.32694, 43.32615, 43.32512, 43.32388, 43.32241, 43.32072, 
    43.31881, 43.31668, 43.31432, 43.31174, 43.30894, 43.30591, 43.30266, 
    43.29919, 43.2955, 43.29158, 43.28744, 43.28308, 43.2785, 43.27369, 
    43.26867, 43.26342, 43.25795, 43.25225, 43.24634, 43.2402, 43.23384, 
    43.22726, 43.22046, 43.21344, 43.20619, 43.19873, 43.19104, 43.18314, 
    43.17501, 43.16666, 43.15809, 43.1493, 43.14029, 43.13106, 43.12161, 
    43.11194, 43.10205, 43.09194, 43.08161, 43.07106, 43.06029, 43.0493, 
    43.0381, 43.02668, 43.01503, 43.00317, 42.99109, 42.97879, 42.96628, 
    42.95354, 42.94059, 42.92743, 42.91404, 42.90044, 42.88662, 42.87259, 
    42.85833, 42.84386, 42.82918, 42.81428, 42.79916, 42.78383, 42.76829, 
    42.75253, 42.73655, 42.72036, 42.70396, 42.68734, 42.67051, 42.65346, 
    42.6362, 42.61873, 42.60105, 42.58315, 42.56504, 42.54672, 42.52819, 
    42.50944, 42.49049, 42.47132, 42.45194, 42.43235, 42.41256, 42.39254, 
    42.37233, 42.3519, 42.33126, 42.31042, 42.28936, 42.2681, 42.24663, 
    42.22495, 42.20306, 42.18097, 42.15867, 42.13616, 42.11345, 42.09053, 
    42.06741, 42.04408, 42.02054, 41.9968, 41.97286, 41.94871, 41.92436, 
    41.8998, 41.87504, 41.85008, 41.82492, 41.79955, 41.77398, 41.74821, 
    41.72224, 41.69607, 41.6697, 41.64313, 41.61636, 41.58938, 41.56221, 
    41.53484, 41.50727, 41.47951, 41.45155, 41.42339, 41.39503, 41.36647, 
    41.33772, 41.30877, 41.27963, 41.25029, 41.22076, 41.19103, 41.16111, 
    41.13099, 41.10068, 41.07018, 41.03949, 41.0086, 40.97752, 40.94625, 
    40.91479, 40.88313, 40.85129, 40.81926, 40.78704, 40.75462, 40.72202, 
    40.68923, 40.65625, 40.62309, 40.58974, 40.5562, 40.52247, 40.48856, 
    40.45446, 40.42018, 40.38571, 40.35106, 40.31622, 40.2812, 40.24599, 
    40.21061, 40.17504,
  36.23239, 36.28315, 36.33376, 36.38424, 36.43457, 36.48475, 36.53479, 
    36.58469, 36.63443, 36.68404, 36.73349, 36.7828, 36.83196, 36.88098, 
    36.92984, 36.97856, 37.02713, 37.07554, 37.12381, 37.17193, 37.21989, 
    37.26771, 37.31537, 37.36288, 37.41024, 37.45744, 37.5045, 37.55139, 
    37.59814, 37.64473, 37.69116, 37.73743, 37.78355, 37.82952, 37.87533, 
    37.92098, 37.96647, 38.0118, 38.05698, 38.102, 38.14685, 38.19155, 
    38.23608, 38.28046, 38.32467, 38.36872, 38.41262, 38.45634, 38.49991, 
    38.54331, 38.58655, 38.62962, 38.67253, 38.71527, 38.75785, 38.80026, 
    38.8425, 38.88458, 38.92649, 38.96824, 39.00981, 39.05121, 39.09245, 
    39.13352, 39.17442, 39.21514, 39.2557, 39.29609, 39.3363, 39.37634, 
    39.41621, 39.45591, 39.49543, 39.53477, 39.57395, 39.61295, 39.65178, 
    39.69043, 39.7289, 39.7672, 39.80532, 39.84327, 39.88103, 39.91862, 
    39.95603, 39.99326, 40.03032, 40.06719, 40.10388, 40.14039, 40.17672, 
    40.21288, 40.24884, 40.28463, 40.32024, 40.35566, 40.3909, 40.42595, 
    40.46082, 40.49551, 40.53001, 40.56432, 40.59845, 40.6324, 40.66616, 
    40.69973, 40.73311, 40.76631, 40.79932, 40.83213, 40.86477, 40.89721, 
    40.92946, 40.96152, 40.99339, 41.02507, 41.05656, 41.08786, 41.11897, 
    41.14988, 41.1806, 41.21113, 41.24147, 41.27161, 41.30156, 41.33131, 
    41.36087, 41.39023, 41.4194, 41.44836, 41.47714, 41.50572, 41.5341, 
    41.56228, 41.59027, 41.61805, 41.64565, 41.67303, 41.70023, 41.72721, 
    41.75401, 41.7806, 41.80699, 41.83318, 41.85917, 41.88496, 41.91054, 
    41.93592, 41.96111, 41.98608, 42.01086, 42.03543, 42.05979, 42.08395, 
    42.10791, 42.13167, 42.15522, 42.17856, 42.20169, 42.22462, 42.24735, 
    42.26987, 42.29218, 42.31428, 42.33618, 42.35787, 42.37935, 42.40062, 
    42.42168, 42.44254, 42.46318, 42.48362, 42.50384, 42.52386, 42.54366, 
    42.56326, 42.58264, 42.60181, 42.62077, 42.63952, 42.65805, 42.67638, 
    42.69449, 42.71239, 42.73008, 42.74755, 42.76481, 42.78185, 42.79869, 
    42.8153, 42.83171, 42.84789, 42.86387, 42.87963, 42.89517, 42.9105, 
    42.92561, 42.9405, 42.95518, 42.96965, 42.98389, 42.99792, 43.01173, 
    43.02533, 43.03871, 43.05187, 43.06481, 43.07753, 43.09004, 43.10233, 
    43.1144, 43.12625, 43.13788, 43.1493, 43.16049, 43.17146, 43.18222, 
    43.19275, 43.20307, 43.21317, 43.22304, 43.2327, 43.24213, 43.25135, 
    43.26034, 43.26911, 43.27766, 43.286, 43.29411, 43.30199, 43.30966, 
    43.3171, 43.32433, 43.33133, 43.33811, 43.34467, 43.35101, 43.35712, 
    43.36301, 43.36868, 43.37413, 43.37936, 43.38436, 43.38914, 43.3937, 
    43.39803, 43.40214, 43.40603, 43.40969, 43.41314, 43.41636, 43.41936, 
    43.42213, 43.42468, 43.42701, 43.42911, 43.43099, 43.43265, 43.43409, 
    43.4353, 43.43628, 43.43705, 43.43759, 43.4379, 43.438, 43.43787, 
    43.43752, 43.43694, 43.43614, 43.43512, 43.43387, 43.4324, 43.43071, 
    43.42879, 43.42665, 43.42429, 43.42171, 43.4189, 43.41586, 43.41261, 
    43.40913, 43.40543, 43.4015, 43.39736, 43.39299, 43.3884, 43.38358, 
    43.37854, 43.37328, 43.3678, 43.36209, 43.35617, 43.35002, 43.34365, 
    43.33706, 43.33024, 43.3232, 43.31594, 43.30846, 43.30076, 43.29284, 
    43.28469, 43.27633, 43.26774, 43.25893, 43.2499, 43.24065, 43.23118, 
    43.22149, 43.21158, 43.20145, 43.1911, 43.18053, 43.16974, 43.15873, 
    43.14751, 43.13606, 43.12439, 43.1125, 43.1004, 43.08808, 43.07554, 
    43.06278, 43.0498, 43.03661, 43.02319, 43.00956, 42.99572, 42.98166, 
    42.96737, 42.95288, 42.93816, 42.92323, 42.90808, 42.89272, 42.87715, 
    42.86135, 42.84535, 42.82912, 42.81269, 42.79604, 42.77917, 42.76209, 
    42.7448, 42.72729, 42.70957, 42.69164, 42.6735, 42.65514, 42.63657, 
    42.61779, 42.59879, 42.57959, 42.56017, 42.54054, 42.5207, 42.50066, 
    42.4804, 42.45993, 42.43925, 42.41837, 42.39727, 42.37597, 42.35445, 
    42.33273, 42.3108, 42.28867, 42.26632, 42.24377, 42.22101, 42.19805, 
    42.17488, 42.1515, 42.12792, 42.10414, 42.08015, 42.05595, 42.03155, 
    42.00695, 41.98214, 41.95713, 41.93192, 41.90651, 41.88089, 41.85507, 
    41.82905, 41.80283, 41.77641, 41.74978, 41.72296, 41.69594, 41.66871, 
    41.64129, 41.61367, 41.58585, 41.55784, 41.52962, 41.50121, 41.4726, 
    41.44379, 41.41479, 41.3856, 41.3562, 41.32661, 41.29683, 41.26685, 
    41.23668, 41.20631, 41.17576, 41.145, 41.11406, 41.08292, 41.05159, 
    41.02008, 40.98837, 40.95646, 40.92437, 40.89209, 40.85962, 40.82696, 
    40.79411, 40.76107, 40.72784, 40.69443, 40.66083, 40.62704, 40.59307, 
    40.55891, 40.52456, 40.49003, 40.45532, 40.42042, 40.38533, 40.35007, 
    40.31462, 40.27898,
  36.3297, 36.38054, 36.43123, 36.48178, 36.53218, 36.58245, 36.63256, 
    36.68253, 36.73236, 36.78204, 36.83157, 36.88095, 36.93019, 36.97927, 
    37.02821, 37.07701, 37.12565, 37.17414, 37.22248, 37.27068, 37.31871, 
    37.3666, 37.41434, 37.46193, 37.50936, 37.55664, 37.60376, 37.65073, 
    37.69755, 37.74421, 37.79072, 37.83707, 37.88327, 37.92931, 37.97519, 
    38.02091, 38.06647, 38.11188, 38.15713, 38.20222, 38.24715, 38.29192, 
    38.33652, 38.38097, 38.42526, 38.46938, 38.51335, 38.55714, 38.60078, 
    38.64425, 38.68756, 38.73071, 38.77369, 38.8165, 38.85915, 38.90163, 
    38.94395, 38.98609, 39.02807, 39.06989, 39.11153, 39.15301, 39.19431, 
    39.23545, 39.27642, 39.31721, 39.35784, 39.39829, 39.43858, 39.47869, 
    39.51862, 39.55839, 39.59798, 39.63739, 39.67664, 39.71571, 39.7546, 
    39.79332, 39.83186, 39.87022, 39.90841, 39.94642, 39.98425, 40.02191, 
    40.05938, 40.09668, 40.1338, 40.17074, 40.2075, 40.24407, 40.28047, 
    40.31668, 40.35272, 40.38857, 40.42424, 40.45972, 40.49502, 40.53014, 
    40.56507, 40.59982, 40.63438, 40.66876, 40.70296, 40.73696, 40.77078, 
    40.80441, 40.83786, 40.87111, 40.90418, 40.93706, 40.96975, 41.00225, 
    41.03456, 41.06668, 41.09862, 41.13036, 41.1619, 41.19326, 41.22442, 
    41.25539, 41.28617, 41.31676, 41.34715, 41.37735, 41.40735, 41.43716, 
    41.46677, 41.49619, 41.52541, 41.55444, 41.58327, 41.6119, 41.64033, 
    41.66857, 41.69661, 41.72445, 41.75209, 41.77953, 41.80677, 41.83382, 
    41.86066, 41.8873, 41.91374, 41.93998, 41.96602, 41.99186, 42.01749, 
    42.04292, 42.06815, 42.09318, 42.118, 42.14262, 42.16703, 42.19124, 
    42.21525, 42.23905, 42.26264, 42.28603, 42.30921, 42.33219, 42.35496, 
    42.37752, 42.39987, 42.42202, 42.44396, 42.46569, 42.48721, 42.50853, 
    42.52963, 42.55053, 42.57121, 42.59169, 42.61195, 42.63201, 42.65185, 
    42.67148, 42.6909, 42.71011, 42.72911, 42.7479, 42.76647, 42.78483, 
    42.80298, 42.82092, 42.83864, 42.85614, 42.87344, 42.89052, 42.90738, 
    42.92403, 42.94047, 42.95669, 42.9727, 42.98849, 43.00406, 43.01942, 
    43.03456, 43.04949, 43.0642, 43.07869, 43.09296, 43.10702, 43.12086, 
    43.13448, 43.14789, 43.16108, 43.17405, 43.1868, 43.19933, 43.21164, 
    43.22374, 43.23561, 43.24726, 43.2587, 43.26992, 43.28092, 43.29169, 
    43.30225, 43.31259, 43.3227, 43.3326, 43.34227, 43.35173, 43.36096, 
    43.36997, 43.37877, 43.38733, 43.39568, 43.40381, 43.41171, 43.4194, 
    43.42686, 43.43409, 43.44111, 43.44791, 43.45448, 43.46083, 43.46695, 
    43.47286, 43.47854, 43.484, 43.48923, 43.49425, 43.49904, 43.5036, 
    43.50795, 43.51207, 43.51596, 43.51964, 43.52309, 43.52631, 43.52932, 
    43.5321, 43.53465, 43.53698, 43.53909, 43.54098, 43.54264, 43.54408, 
    43.54529, 43.54628, 43.54705, 43.54759, 43.5479, 43.548, 43.54787, 
    43.54752, 43.54694, 43.54614, 43.54511, 43.54387, 43.54239, 43.5407, 
    43.53878, 43.53663, 43.53426, 43.53167, 43.52886, 43.52582, 43.52256, 
    43.51907, 43.51536, 43.51143, 43.50727, 43.5029, 43.49829, 43.49347, 
    43.48842, 43.48315, 43.47766, 43.47194, 43.466, 43.45984, 43.45345, 
    43.44685, 43.44002, 43.43296, 43.42569, 43.41819, 43.41048, 43.40254, 
    43.39437, 43.38599, 43.37739, 43.36856, 43.35952, 43.35025, 43.34076, 
    43.33105, 43.32112, 43.31097, 43.30059, 43.29, 43.27919, 43.26816, 
    43.25691, 43.24544, 43.23375, 43.22184, 43.20971, 43.19736, 43.1848, 
    43.17201, 43.159, 43.14578, 43.13234, 43.11869, 43.10481, 43.09072, 
    43.07641, 43.06188, 43.04714, 43.03218, 43.017, 43.00161, 42.986, 
    42.97018, 42.95414, 42.93789, 42.92141, 42.90473, 42.88783, 42.87072, 
    42.85339, 42.83585, 42.81809, 42.80013, 42.78194, 42.76355, 42.74494, 
    42.72612, 42.70709, 42.68785, 42.66839, 42.64872, 42.62885, 42.60876, 
    42.58846, 42.56795, 42.54723, 42.52631, 42.50517, 42.48382, 42.46227, 
    42.4405, 42.41853, 42.39635, 42.37396, 42.35137, 42.32857, 42.30556, 
    42.28234, 42.25892, 42.23529, 42.21146, 42.18743, 42.16319, 42.13874, 
    42.11409, 42.08923, 42.06417, 42.03891, 42.01345, 41.98779, 41.96192, 
    41.93584, 41.90957, 41.8831, 41.85643, 41.82955, 41.80248, 41.7752, 
    41.74773, 41.72006, 41.69218, 41.66412, 41.63585, 41.60738, 41.57872, 
    41.54986, 41.5208, 41.49155, 41.4621, 41.43246, 41.40262, 41.37259, 
    41.34236, 41.31194, 41.28132, 41.25051, 41.21951, 41.18831, 41.15693, 
    41.12535, 41.09358, 41.06162, 41.02947, 40.99712, 40.9646, 40.93187, 
    40.89896, 40.86587, 40.83258, 40.79911, 40.76545, 40.73159, 40.69756, 
    40.66334, 40.62893, 40.59434, 40.55956, 40.5246, 40.48945, 40.45412, 
    40.41861, 40.38291,
  36.42699, 36.4779, 36.52867, 36.57929, 36.62977, 36.68011, 36.7303, 
    36.78035, 36.83025, 36.88, 36.9296, 36.97906, 37.02838, 37.07754, 
    37.12656, 37.17542, 37.22414, 37.27271, 37.32113, 37.36939, 37.41751, 
    37.46547, 37.51328, 37.56094, 37.60845, 37.6558, 37.703, 37.75005, 
    37.79694, 37.84367, 37.89025, 37.93668, 37.98295, 38.02906, 38.07501, 
    38.12081, 38.16645, 38.21193, 38.25725, 38.30241, 38.34742, 38.39226, 
    38.43694, 38.48146, 38.52582, 38.57001, 38.61405, 38.65792, 38.70163, 
    38.74517, 38.78855, 38.83177, 38.87482, 38.91771, 38.96042, 39.00298, 
    39.04536, 39.08758, 39.12963, 39.17152, 39.21323, 39.25478, 39.29615, 
    39.33736, 39.3784, 39.41926, 39.45996, 39.50048, 39.54083, 39.58101, 
    39.62101, 39.66085, 39.70051, 39.73999, 39.7793, 39.81844, 39.8574, 
    39.89618, 39.93479, 39.97322, 40.01148, 40.04956, 40.08746, 40.12518, 
    40.16272, 40.20008, 40.23726, 40.27427, 40.31109, 40.34773, 40.38419, 
    40.42048, 40.45657, 40.49249, 40.52822, 40.56377, 40.59913, 40.63431, 
    40.66931, 40.70412, 40.73875, 40.77319, 40.80744, 40.84151, 40.87539, 
    40.90908, 40.94258, 40.9759, 41.00903, 41.04197, 41.07472, 41.10728, 
    41.13966, 41.17184, 41.20382, 41.23562, 41.26723, 41.29865, 41.32986, 
    41.36089, 41.39173, 41.42237, 41.45282, 41.48307, 41.51313, 41.543, 
    41.57267, 41.60214, 41.63142, 41.6605, 41.68938, 41.71806, 41.74655, 
    41.77485, 41.80294, 41.83083, 41.85852, 41.88602, 41.91331, 41.94041, 
    41.9673, 41.99399, 42.02048, 42.04678, 42.07286, 42.09875, 42.12444, 
    42.14991, 42.17519, 42.20027, 42.22514, 42.2498, 42.27427, 42.29852, 
    42.32257, 42.34642, 42.37006, 42.39349, 42.41672, 42.43974, 42.46255, 
    42.48516, 42.50756, 42.52975, 42.55173, 42.57351, 42.59507, 42.61642, 
    42.63757, 42.65851, 42.67923, 42.69975, 42.72005, 42.74015, 42.76003, 
    42.77971, 42.79916, 42.81841, 42.83745, 42.85627, 42.87488, 42.89328, 
    42.91146, 42.92944, 42.94719, 42.96473, 42.98206, 42.99918, 43.01608, 
    43.03276, 43.04923, 43.06548, 43.08152, 43.09734, 43.11295, 43.12834, 
    43.14351, 43.15847, 43.17321, 43.18773, 43.20203, 43.21612, 43.22998, 
    43.24364, 43.25707, 43.27028, 43.28328, 43.29605, 43.30861, 43.32095, 
    43.33307, 43.34497, 43.35665, 43.36811, 43.37935, 43.39037, 43.40117, 
    43.41174, 43.4221, 43.43224, 43.44215, 43.45185, 43.46132, 43.47058, 
    43.47961, 43.48841, 43.497, 43.50537, 43.51351, 43.52143, 43.52913, 
    43.53661, 43.54386, 43.55089, 43.5577, 43.56429, 43.57065, 43.57679, 
    43.5827, 43.5884, 43.59387, 43.59911, 43.60414, 43.60894, 43.61351, 
    43.61787, 43.62199, 43.6259, 43.62958, 43.63304, 43.63627, 43.63928, 
    43.64206, 43.64463, 43.64696, 43.64907, 43.65096, 43.65263, 43.65407, 
    43.65528, 43.65628, 43.65704, 43.65759, 43.65791, 43.658, 43.65787, 
    43.65752, 43.65694, 43.65614, 43.65511, 43.65385, 43.65238, 43.65068, 
    43.64875, 43.64661, 43.64423, 43.64164, 43.63882, 43.63577, 43.6325, 
    43.62901, 43.62529, 43.62136, 43.61719, 43.6128, 43.60819, 43.60336, 
    43.5983, 43.59302, 43.58751, 43.58178, 43.57583, 43.56966, 43.56326, 
    43.55664, 43.54979, 43.54273, 43.53544, 43.52793, 43.5202, 43.51224, 
    43.50406, 43.49566, 43.48704, 43.47819, 43.46913, 43.45984, 43.45033, 
    43.4406, 43.43065, 43.42048, 43.41008, 43.39947, 43.38864, 43.37758, 
    43.36631, 43.35482, 43.3431, 43.33117, 43.31901, 43.30664, 43.29405, 
    43.28124, 43.26821, 43.25496, 43.24149, 43.22781, 43.21391, 43.19978, 
    43.18544, 43.17089, 43.15612, 43.14112, 43.12592, 43.11049, 43.09486, 
    43.079, 43.06293, 43.04664, 43.03014, 43.01342, 42.99648, 42.97934, 
    42.96198, 42.9444, 42.92661, 42.9086, 42.89038, 42.87195, 42.85331, 
    42.83445, 42.81538, 42.7961, 42.77661, 42.7569, 42.73698, 42.71686, 
    42.69652, 42.67597, 42.65521, 42.63424, 42.61306, 42.59167, 42.57008, 
    42.54827, 42.52625, 42.50403, 42.4816, 42.45896, 42.43611, 42.41306, 
    42.3898, 42.36633, 42.34266, 42.31878, 42.2947, 42.27041, 42.24591, 
    42.22122, 42.19632, 42.17121, 42.1459, 42.12038, 42.09467, 42.06875, 
    42.04263, 42.01631, 41.98978, 41.96306, 41.93613, 41.90901, 41.88168, 
    41.85416, 41.82643, 41.7985, 41.77038, 41.74206, 41.71354, 41.68482, 
    41.65591, 41.6268, 41.59749, 41.56799, 41.53829, 41.50839, 41.4783, 
    41.44802, 41.41754, 41.38686, 41.356, 41.32494, 41.29369, 41.26224, 
    41.23061, 41.19878, 41.16676, 41.13455, 41.10215, 41.06956, 41.03677, 
    41.00381, 40.97065, 40.9373, 40.90376, 40.87004, 40.83613, 40.80203, 
    40.76775, 40.73328, 40.69862, 40.66378, 40.62876, 40.59355, 40.55816, 
    40.52258, 40.48682,
  36.52423, 36.57522, 36.62606, 36.67677, 36.72732, 36.77774, 36.828, 
    36.87812, 36.9281, 36.97793, 37.02761, 37.07714, 37.12653, 37.17577, 
    37.22486, 37.2738, 37.3226, 37.37124, 37.41973, 37.46807, 37.51627, 
    37.5643, 37.61219, 37.65992, 37.7075, 37.75493, 37.80221, 37.84933, 
    37.89629, 37.9431, 37.98976, 38.03626, 38.0826, 38.12878, 38.17481, 
    38.22068, 38.2664, 38.31195, 38.35735, 38.40258, 38.44765, 38.49257, 
    38.53732, 38.58192, 38.62635, 38.67062, 38.71472, 38.75867, 38.80245, 
    38.84607, 38.88951, 38.9328, 38.97593, 39.01888, 39.06167, 39.1043, 
    39.14676, 39.18904, 39.23117, 39.27312, 39.3149, 39.35652, 39.39797, 
    39.43924, 39.48035, 39.52129, 39.56205, 39.60264, 39.64306, 39.68331, 
    39.72338, 39.76329, 39.80301, 39.84257, 39.88195, 39.92115, 39.96018, 
    39.99903, 40.0377, 40.0762, 40.11452, 40.15267, 40.19064, 40.22842, 
    40.26603, 40.30346, 40.34071, 40.37778, 40.41467, 40.45137, 40.4879, 
    40.52424, 40.56041, 40.59638, 40.63218, 40.66779, 40.70322, 40.73846, 
    40.77353, 40.8084, 40.84309, 40.87759, 40.91191, 40.94603, 40.97998, 
    41.01373, 41.0473, 41.08068, 41.11386, 41.14687, 41.17968, 41.2123, 
    41.24473, 41.27697, 41.30902, 41.34087, 41.37254, 41.40401, 41.43529, 
    41.46638, 41.49727, 41.52797, 41.55848, 41.58879, 41.6189, 41.64882, 
    41.67855, 41.70808, 41.73741, 41.76654, 41.79548, 41.82422, 41.85276, 
    41.88111, 41.90925, 41.9372, 41.96494, 41.99249, 42.01984, 42.04698, 
    42.07393, 42.10067, 42.12722, 42.15356, 42.1797, 42.20563, 42.23137, 
    42.2569, 42.28222, 42.30735, 42.33226, 42.35698, 42.38148, 42.40579, 
    42.42989, 42.45378, 42.47747, 42.50095, 42.52422, 42.54728, 42.57014, 
    42.59279, 42.61523, 42.63747, 42.6595, 42.68131, 42.70292, 42.72432, 
    42.7455, 42.76648, 42.78725, 42.8078, 42.82815, 42.84829, 42.86821, 
    42.88792, 42.90742, 42.9267, 42.94578, 42.96464, 42.98329, 43.00172, 
    43.01994, 43.03795, 43.05574, 43.07332, 43.09068, 43.10783, 43.12476, 
    43.14148, 43.15799, 43.17427, 43.19034, 43.2062, 43.22183, 43.23725, 
    43.25246, 43.26744, 43.28221, 43.29676, 43.3111, 43.32521, 43.33911, 
    43.35279, 43.36625, 43.37949, 43.39251, 43.40531, 43.41789, 43.43026, 
    43.4424, 43.45432, 43.46603, 43.47751, 43.48877, 43.49981, 43.51064, 
    43.52124, 43.53162, 43.54177, 43.55171, 43.56142, 43.57092, 43.58019, 
    43.58924, 43.59806, 43.60667, 43.61505, 43.62321, 43.63115, 43.63886, 
    43.64635, 43.65363, 43.66067, 43.66749, 43.67409, 43.68047, 43.68662, 
    43.69255, 43.69825, 43.70374, 43.70899, 43.71402, 43.71883, 43.72342, 
    43.72778, 43.73192, 43.73583, 43.73952, 43.74298, 43.74622, 43.74924, 
    43.75203, 43.7546, 43.75694, 43.75906, 43.76095, 43.76262, 43.76406, 
    43.76528, 43.76627, 43.76704, 43.76759, 43.76791, 43.768, 43.76787, 
    43.76751, 43.76693, 43.76613, 43.7651, 43.76385, 43.76237, 43.76067, 
    43.75874, 43.75658, 43.75421, 43.75161, 43.74878, 43.74573, 43.74245, 
    43.73895, 43.73523, 43.73128, 43.72711, 43.72271, 43.71809, 43.71325, 
    43.70818, 43.70288, 43.69736, 43.69162, 43.68566, 43.67947, 43.67306, 
    43.66643, 43.65957, 43.65249, 43.64518, 43.63766, 43.62991, 43.62194, 
    43.61374, 43.60532, 43.59668, 43.58782, 43.57874, 43.56943, 43.5599, 
    43.55015, 43.54018, 43.52999, 43.51957, 43.50894, 43.49808, 43.48701, 
    43.47571, 43.46419, 43.45245, 43.44049, 43.42831, 43.41592, 43.4033, 
    43.39046, 43.37741, 43.36413, 43.35064, 43.33692, 43.32299, 43.30884, 
    43.29448, 43.27989, 43.26509, 43.25006, 43.23483, 43.21937, 43.2037, 
    43.18781, 43.17171, 43.15539, 43.13885, 43.1221, 43.10513, 43.08795, 
    43.07055, 43.05294, 43.03511, 43.01707, 42.99882, 42.98035, 42.96167, 
    42.94278, 42.92367, 42.90435, 42.88482, 42.86507, 42.84512, 42.82495, 
    42.80457, 42.78398, 42.76318, 42.74217, 42.72095, 42.69952, 42.67788, 
    42.65602, 42.63396, 42.6117, 42.58922, 42.56654, 42.54365, 42.52055, 
    42.49725, 42.47373, 42.45002, 42.42609, 42.40196, 42.37762, 42.35308, 
    42.32833, 42.30338, 42.27823, 42.25287, 42.22731, 42.20154, 42.17558, 
    42.1494, 42.12303, 42.09645, 42.06968, 42.0427, 42.01553, 41.98815, 
    41.96057, 41.93279, 41.90481, 41.87664, 41.84826, 41.81969, 41.79092, 
    41.76195, 41.73278, 41.70342, 41.67386, 41.6441, 41.61415, 41.584, 
    41.55367, 41.52313, 41.4924, 41.46147, 41.43036, 41.39904, 41.36754, 
    41.33585, 41.30396, 41.27188, 41.23961, 41.20715, 41.1745, 41.14166, 
    41.10863, 41.07541, 41.042, 41.0084, 40.97462, 40.94065, 40.90649, 
    40.87214, 40.83761, 40.80289, 40.76799, 40.7329, 40.69763, 40.66217, 
    40.62653, 40.59071,
  36.62144, 36.67251, 36.72343, 36.77421, 36.82484, 36.87533, 36.92567, 
    36.97587, 37.02592, 37.07582, 37.12558, 37.17519, 37.22466, 37.27398, 
    37.32314, 37.37216, 37.42102, 37.46974, 37.51831, 37.56673, 37.61499, 
    37.66311, 37.71107, 37.75888, 37.80653, 37.85403, 37.90139, 37.94858, 
    37.99562, 38.0425, 38.08923, 38.13581, 38.18222, 38.22848, 38.27458, 
    38.32053, 38.36631, 38.41194, 38.45741, 38.50272, 38.54787, 38.59285, 
    38.63768, 38.68235, 38.72685, 38.77119, 38.81537, 38.85939, 38.90324, 
    38.94693, 38.99045, 39.03381, 39.077, 39.12003, 39.1629, 39.20559, 
    39.24812, 39.29048, 39.33267, 39.3747, 39.41655, 39.45824, 39.49976, 
    39.5411, 39.58228, 39.62328, 39.66412, 39.70478, 39.74527, 39.78559, 
    39.82573, 39.8657, 39.90549, 39.94512, 39.98457, 40.02383, 40.06293, 
    40.10185, 40.14059, 40.17916, 40.21755, 40.25576, 40.29379, 40.33165, 
    40.36932, 40.40681, 40.44413, 40.48127, 40.51822, 40.55499, 40.59158, 
    40.62799, 40.66422, 40.70026, 40.73612, 40.7718, 40.80729, 40.8426, 
    40.87772, 40.91266, 40.94741, 40.98198, 41.01635, 41.05054, 41.08455, 
    41.11837, 41.15199, 41.18543, 41.21868, 41.25174, 41.28461, 41.3173, 
    41.34978, 41.38208, 41.41419, 41.44611, 41.47783, 41.50937, 41.5407, 
    41.57185, 41.6028, 41.63355, 41.66412, 41.69448, 41.72466, 41.75463, 
    41.78441, 41.814, 41.84338, 41.87257, 41.90157, 41.93036, 41.95896, 
    41.98735, 42.01555, 42.04355, 42.07135, 42.09895, 42.12635, 42.15355, 
    42.18055, 42.20734, 42.23394, 42.26033, 42.28652, 42.3125, 42.33829, 
    42.36386, 42.38924, 42.41441, 42.43938, 42.46414, 42.4887, 42.51305, 
    42.53719, 42.56113, 42.58487, 42.60839, 42.63171, 42.65482, 42.67772, 
    42.70042, 42.7229, 42.74518, 42.76725, 42.78911, 42.81076, 42.8322, 
    42.85343, 42.87445, 42.89526, 42.91586, 42.93624, 42.95642, 42.97638, 
    42.99613, 43.01567, 43.03499, 43.0541, 43.073, 43.09169, 43.11016, 
    43.12841, 43.14646, 43.16429, 43.1819, 43.1993, 43.21648, 43.23345, 
    43.2502, 43.26674, 43.28305, 43.29916, 43.31504, 43.33071, 43.34616, 
    43.3614, 43.37642, 43.39121, 43.40579, 43.42015, 43.4343, 43.44822, 
    43.46193, 43.47542, 43.48869, 43.50174, 43.51456, 43.52717, 43.53956, 
    43.55173, 43.56367, 43.57541, 43.58691, 43.5982, 43.60926, 43.62011, 
    43.63073, 43.64113, 43.65131, 43.66126, 43.671, 43.68051, 43.6898, 
    43.69887, 43.70771, 43.71634, 43.72474, 43.73291, 43.74086, 43.7486, 
    43.7561, 43.76339, 43.77045, 43.77728, 43.7839, 43.79029, 43.79645, 
    43.80239, 43.80811, 43.8136, 43.81887, 43.82391, 43.82873, 43.83333, 
    43.8377, 43.84184, 43.84576, 43.84946, 43.85293, 43.85618, 43.8592, 
    43.862, 43.86457, 43.86692, 43.86904, 43.87093, 43.8726, 43.87405, 
    43.87527, 43.87627, 43.87704, 43.87759, 43.8779, 43.878, 43.87787, 
    43.87751, 43.87693, 43.87613, 43.8751, 43.87384, 43.87236, 43.87065, 
    43.86872, 43.86656, 43.86418, 43.86157, 43.85874, 43.85568, 43.8524, 
    43.84889, 43.84516, 43.8412, 43.83702, 43.83261, 43.82798, 43.82313, 
    43.81805, 43.81275, 43.80722, 43.80147, 43.79549, 43.78929, 43.78286, 
    43.77622, 43.76934, 43.76225, 43.75493, 43.74739, 43.73962, 43.73163, 
    43.72342, 43.71498, 43.70633, 43.69745, 43.68835, 43.67902, 43.66947, 
    43.6597, 43.64971, 43.6395, 43.62906, 43.6184, 43.60752, 43.59642, 
    43.58511, 43.57356, 43.5618, 43.54982, 43.53762, 43.52519, 43.51255, 
    43.49968, 43.4866, 43.4733, 43.45978, 43.44604, 43.43208, 43.4179, 
    43.4035, 43.38889, 43.37405, 43.359, 43.34373, 43.32825, 43.31255, 
    43.29662, 43.28049, 43.26413, 43.24757, 43.23078, 43.21378, 43.19656, 
    43.17913, 43.16148, 43.14362, 43.12554, 43.10725, 43.08875, 43.07003, 
    43.05109, 43.03195, 43.01259, 42.99302, 42.97324, 42.95324, 42.93303, 
    42.91261, 42.89198, 42.87114, 42.85009, 42.82882, 42.80735, 42.78567, 
    42.76377, 42.74167, 42.71936, 42.69684, 42.67411, 42.65118, 42.62803, 
    42.60468, 42.58112, 42.55736, 42.53339, 42.50921, 42.48483, 42.46024, 
    42.43544, 42.41044, 42.38524, 42.35983, 42.33422, 42.30841, 42.28239, 
    42.25617, 42.22974, 42.20312, 42.17629, 42.14926, 42.12203, 42.0946, 
    42.06697, 42.03914, 42.0111, 41.98288, 41.95445, 41.92582, 41.89699, 
    41.86797, 41.83875, 41.80933, 41.77972, 41.7499, 41.71989, 41.68969, 
    41.65929, 41.6287, 41.59792, 41.56693, 41.53576, 41.50439, 41.47283, 
    41.44107, 41.40913, 41.37699, 41.34466, 41.31214, 41.27943, 41.24653, 
    41.21344, 41.18016, 41.14669, 41.11303, 41.07918, 41.04515, 41.01093, 
    40.97652, 40.94193, 40.90714, 40.87218, 40.83702, 40.80169, 40.76617, 
    40.73046, 40.69457,
  36.71862, 36.76977, 36.82076, 36.87162, 36.92233, 36.97289, 37.02331, 
    37.07358, 37.12371, 37.17369, 37.22353, 37.27321, 37.32275, 37.37214, 
    37.42138, 37.47047, 37.51942, 37.56821, 37.61686, 37.66535, 37.71369, 
    37.76188, 37.80991, 37.8578, 37.90553, 37.95311, 38.00053, 38.0478, 
    38.09491, 38.14187, 38.18867, 38.23532, 38.28181, 38.32815, 38.37432, 
    38.42034, 38.4662, 38.5119, 38.55745, 38.60283, 38.64805, 38.69311, 
    38.73801, 38.78275, 38.82732, 38.87174, 38.91599, 38.96008, 39.00401, 
    39.04776, 39.09136, 39.13479, 39.17806, 39.22116, 39.26409, 39.30686, 
    39.34946, 39.39189, 39.43415, 39.47625, 39.51818, 39.55993, 39.60152, 
    39.64294, 39.68418, 39.72526, 39.76616, 39.80689, 39.84745, 39.88784, 
    39.92805, 39.96809, 40.00795, 40.04765, 40.08716, 40.1265, 40.16566, 
    40.20465, 40.24346, 40.2821, 40.32055, 40.35883, 40.39693, 40.43485, 
    40.47259, 40.51015, 40.54753, 40.58473, 40.62175, 40.65859, 40.69525, 
    40.73172, 40.76801, 40.80412, 40.84005, 40.87579, 40.91134, 40.94671, 
    40.9819, 41.0169, 41.05172, 41.08634, 41.12078, 41.15504, 41.1891, 
    41.22298, 41.25667, 41.29017, 41.32348, 41.35661, 41.38953, 41.42228, 
    41.45483, 41.48719, 41.51935, 41.55133, 41.58311, 41.6147, 41.6461, 
    41.6773, 41.70831, 41.73912, 41.76974, 41.80017, 41.83039, 41.86043, 
    41.89027, 41.91991, 41.94935, 41.97859, 42.00764, 42.03649, 42.06514, 
    42.09359, 42.12185, 42.1499, 42.17775, 42.2054, 42.23285, 42.26011, 
    42.28715, 42.314, 42.34064, 42.36709, 42.39333, 42.41936, 42.44519, 
    42.47083, 42.49625, 42.52147, 42.54649, 42.5713, 42.5959, 42.6203, 
    42.64449, 42.66848, 42.69225, 42.71583, 42.73919, 42.76235, 42.78529, 
    42.80803, 42.83057, 42.85289, 42.875, 42.8969, 42.91859, 42.94008, 
    42.96135, 42.98241, 43.00326, 43.0239, 43.04432, 43.06454, 43.08454, 
    43.10433, 43.12391, 43.14327, 43.16242, 43.18136, 43.20008, 43.21859, 
    43.23688, 43.25496, 43.27283, 43.29047, 43.30791, 43.32513, 43.34213, 
    43.35891, 43.37548, 43.39183, 43.40797, 43.42389, 43.43959, 43.45507, 
    43.47034, 43.48538, 43.50021, 43.51482, 43.52921, 43.54338, 43.55734, 
    43.57108, 43.58459, 43.59788, 43.61096, 43.62381, 43.63645, 43.64886, 
    43.66106, 43.67303, 43.68478, 43.69631, 43.70762, 43.7187, 43.72957, 
    43.74022, 43.75064, 43.76084, 43.77081, 43.78057, 43.7901, 43.79941, 
    43.80849, 43.81736, 43.826, 43.83442, 43.84261, 43.85058, 43.85833, 
    43.86585, 43.87315, 43.88022, 43.88707, 43.8937, 43.9001, 43.90628, 
    43.91224, 43.91796, 43.92347, 43.92875, 43.9338, 43.93863, 43.94323, 
    43.94761, 43.95177, 43.9557, 43.9594, 43.96288, 43.96613, 43.96916, 
    43.97197, 43.97454, 43.97689, 43.97902, 43.98092, 43.98259, 43.98404, 
    43.98527, 43.98626, 43.98704, 43.98758, 43.9879, 43.988, 43.98787, 
    43.98751, 43.98693, 43.98612, 43.98509, 43.98383, 43.98235, 43.98063, 
    43.9787, 43.97654, 43.97415, 43.97153, 43.9687, 43.96563, 43.96235, 
    43.95883, 43.95509, 43.95113, 43.94694, 43.94252, 43.93788, 43.93302, 
    43.92793, 43.92261, 43.91707, 43.91131, 43.90532, 43.89911, 43.89267, 
    43.88601, 43.87912, 43.87201, 43.86467, 43.85712, 43.84933, 43.84133, 
    43.8331, 43.82465, 43.81597, 43.80708, 43.79795, 43.78861, 43.77904, 
    43.76925, 43.75924, 43.749, 43.73854, 43.72787, 43.71696, 43.70584, 
    43.6945, 43.68293, 43.67115, 43.65914, 43.64691, 43.63446, 43.6218, 
    43.60891, 43.59579, 43.58247, 43.56892, 43.55515, 43.54116, 43.52695, 
    43.51252, 43.49788, 43.48302, 43.46794, 43.45264, 43.43712, 43.42138, 
    43.40543, 43.38926, 43.37288, 43.35627, 43.33945, 43.32242, 43.30516, 
    43.2877, 43.27002, 43.25212, 43.234, 43.21568, 43.19713, 43.17838, 
    43.1594, 43.14022, 43.12083, 43.10122, 43.08139, 43.06136, 43.04111, 
    43.02065, 42.99998, 42.97909, 42.958, 42.9367, 42.91518, 42.89345, 
    42.87152, 42.84937, 42.82701, 42.80445, 42.78168, 42.7587, 42.73551, 
    42.71211, 42.68851, 42.6647, 42.64068, 42.61645, 42.59202, 42.56738, 
    42.54254, 42.51749, 42.49224, 42.46679, 42.44112, 42.41526, 42.38919, 
    42.36292, 42.33644, 42.30976, 42.28289, 42.25581, 42.22852, 42.20104, 
    42.17336, 42.14547, 42.11739, 42.0891, 42.06062, 42.03194, 42.00306, 
    41.97398, 41.9447, 41.91523, 41.88556, 41.85569, 41.82563, 41.79537, 
    41.76491, 41.73426, 41.70341, 41.67238, 41.64114, 41.60972, 41.57809, 
    41.54628, 41.51428, 41.48208, 41.44969, 41.41711, 41.38434, 41.35138, 
    41.31823, 41.28489, 41.25135, 41.21764, 41.18373, 41.14963, 41.11535, 
    41.08088, 41.04622, 41.01138, 40.97635, 40.94113, 40.90573, 40.87014, 
    40.83437, 40.79842,
  36.81577, 36.86699, 36.91806, 36.96899, 37.01978, 37.07042, 37.12091, 
    37.17126, 37.22147, 37.27152, 37.32143, 37.3712, 37.42081, 37.47028, 
    37.51959, 37.56876, 37.61778, 37.66665, 37.71537, 37.76394, 37.81235, 
    37.86061, 37.90873, 37.95669, 38.00449, 38.05215, 38.09964, 38.14699, 
    38.19418, 38.24121, 38.28809, 38.33481, 38.38137, 38.42778, 38.47403, 
    38.52013, 38.56606, 38.61184, 38.65745, 38.70291, 38.7482, 38.79333, 
    38.83831, 38.88312, 38.92777, 38.97226, 39.01658, 39.06075, 39.10474, 
    39.14857, 39.19224, 39.23575, 39.27908, 39.32226, 39.36526, 39.4081, 
    39.45077, 39.49327, 39.53561, 39.57777, 39.61977, 39.6616, 39.70326, 
    39.74475, 39.78606, 39.82721, 39.86818, 39.90898, 39.94961, 39.99007, 
    40.03035, 40.07046, 40.11039, 40.15015, 40.18974, 40.22914, 40.26838, 
    40.30743, 40.34631, 40.38501, 40.42353, 40.46188, 40.50005, 40.53803, 
    40.57584, 40.61347, 40.65091, 40.68818, 40.72527, 40.76217, 40.79889, 
    40.83543, 40.87179, 40.90796, 40.94395, 40.97975, 41.01537, 41.05081, 
    41.08606, 41.12112, 41.156, 41.19069, 41.22519, 41.25951, 41.29364, 
    41.32758, 41.36133, 41.39489, 41.42826, 41.46145, 41.49444, 41.52724, 
    41.55985, 41.59227, 41.6245, 41.65653, 41.68837, 41.72002, 41.75148, 
    41.78274, 41.8138, 41.84468, 41.87535, 41.90583, 41.93612, 41.96621, 
    41.9961, 42.0258, 42.0553, 42.0846, 42.1137, 42.1426, 42.17131, 42.19981, 
    42.22812, 42.25623, 42.28413, 42.31184, 42.33934, 42.36665, 42.39375, 
    42.42065, 42.44734, 42.47383, 42.50013, 42.52621, 42.55209, 42.57777, 
    42.60325, 42.62852, 42.65358, 42.67844, 42.70309, 42.72754, 42.75178, 
    42.77581, 42.79964, 42.82325, 42.84666, 42.86987, 42.89286, 42.91564, 
    42.93822, 42.96058, 42.98274, 43.00468, 43.02642, 43.04795, 43.06926, 
    43.09036, 43.11126, 43.13194, 43.1524, 43.17266, 43.1927, 43.21253, 
    43.23214, 43.25154, 43.27073, 43.28971, 43.30847, 43.32701, 43.34534, 
    43.36346, 43.38136, 43.39904, 43.41651, 43.43377, 43.4508, 43.46762, 
    43.48422, 43.50061, 43.51678, 43.53273, 43.54846, 43.56397, 43.57927, 
    43.59435, 43.60921, 43.62385, 43.63827, 43.65247, 43.66645, 43.68021, 
    43.69376, 43.70708, 43.72018, 43.73306, 43.74572, 43.75816, 43.77038, 
    43.78238, 43.79415, 43.80571, 43.81704, 43.82815, 43.83904, 43.8497, 
    43.86015, 43.87037, 43.88036, 43.89014, 43.89969, 43.90902, 43.91813, 
    43.92701, 43.93567, 43.9441, 43.95231, 43.9603, 43.96806, 43.9756, 
    43.98291, 43.99, 43.99686, 44.00351, 44.00992, 44.01611, 44.02208, 
    44.02782, 44.03333, 44.03862, 44.04369, 44.04853, 44.05314, 44.05753, 
    44.06169, 44.06563, 44.06934, 44.07283, 44.07609, 44.07912, 44.08193, 
    44.08451, 44.08687, 44.089, 44.0909, 44.09258, 44.09404, 44.09526, 
    44.09626, 44.09703, 44.09758, 44.0979, 44.098, 44.09787, 44.09751, 
    44.09693, 44.09612, 44.09508, 44.09382, 44.09233, 44.09062, 44.08868, 
    44.08651, 44.08412, 44.0815, 44.07866, 44.07559, 44.07229, 44.06877, 
    44.06502, 44.06105, 44.05685, 44.05243, 44.04778, 44.0429, 44.0378, 
    44.03247, 44.02692, 44.02115, 44.01515, 44.00892, 44.00247, 43.99579, 
    43.98889, 43.98177, 43.97442, 43.96685, 43.95905, 43.95103, 43.94278, 
    43.93431, 43.92562, 43.9167, 43.90756, 43.89819, 43.88861, 43.8788, 
    43.86876, 43.85851, 43.84803, 43.83733, 43.8264, 43.81526, 43.80389, 
    43.7923, 43.78049, 43.76846, 43.75621, 43.74373, 43.73104, 43.71812, 
    43.70499, 43.69163, 43.67805, 43.66425, 43.65024, 43.636, 43.62154, 
    43.60687, 43.59198, 43.57687, 43.56153, 43.54599, 43.53022, 43.51423, 
    43.49803, 43.48161, 43.46497, 43.44812, 43.43105, 43.41376, 43.39626, 
    43.37854, 43.36061, 43.34246, 43.3241, 43.30552, 43.28672, 43.26771, 
    43.24849, 43.22905, 43.2094, 43.18954, 43.16947, 43.14918, 43.12868, 
    43.10796, 43.08704, 43.0659, 43.04456, 43.023, 43.00123, 42.97925, 
    42.95706, 42.93466, 42.91205, 42.88924, 42.86621, 42.84298, 42.81953, 
    42.79588, 42.77202, 42.74796, 42.72369, 42.69921, 42.67452, 42.64963, 
    42.62453, 42.59923, 42.57373, 42.54802, 42.5221, 42.49598, 42.46966, 
    42.44313, 42.4164, 42.38947, 42.36234, 42.33501, 42.30747, 42.27973, 
    42.2518, 42.22366, 42.19532, 42.16678, 42.13805, 42.10911, 42.07998, 
    42.05064, 42.02111, 41.99139, 41.96146, 41.93134, 41.90103, 41.87051, 
    41.83981, 41.8089, 41.77781, 41.74651, 41.71503, 41.68335, 41.65148, 
    41.61941, 41.58715, 41.55471, 41.52206, 41.48923, 41.45621, 41.423, 
    41.3896, 41.356, 41.32222, 41.28825, 41.25409, 41.21975, 41.18521, 
    41.15049, 41.11559, 41.08049, 41.04522, 41.00975, 40.9741, 40.93827, 
    40.90225,
  36.91288, 36.96417, 37.01532, 37.06633, 37.11719, 37.16791, 37.21848, 
    37.26891, 37.31919, 37.36932, 37.41931, 37.46914, 37.51884, 37.56838, 
    37.61777, 37.66702, 37.71611, 37.76506, 37.81385, 37.86249, 37.91098, 
    37.95932, 38.00751, 38.05555, 38.10343, 38.15115, 38.19873, 38.24615, 
    38.29341, 38.34052, 38.38747, 38.43427, 38.48091, 38.52739, 38.57372, 
    38.61988, 38.66589, 38.71174, 38.75743, 38.80296, 38.84832, 38.89353, 
    38.93858, 38.98347, 39.02819, 39.07275, 39.11715, 39.16138, 39.20545, 
    39.24936, 39.2931, 39.33667, 39.38008, 39.42333, 39.4664, 39.50932, 
    39.55206, 39.59463, 39.63704, 39.67928, 39.72134, 39.76324, 39.80497, 
    39.84653, 39.88792, 39.92913, 39.97018, 40.01105, 40.05175, 40.09227, 
    40.13262, 40.1728, 40.2128, 40.25263, 40.29228, 40.33176, 40.37106, 
    40.41018, 40.44913, 40.4879, 40.52649, 40.5649, 40.60314, 40.64119, 
    40.67907, 40.71676, 40.75427, 40.79161, 40.82876, 40.86573, 40.90252, 
    40.93912, 40.97554, 41.01178, 41.04783, 41.0837, 41.11938, 41.15488, 
    41.1902, 41.22533, 41.26027, 41.29502, 41.32959, 41.36397, 41.39816, 
    41.43216, 41.46597, 41.4996, 41.53303, 41.56627, 41.59933, 41.63219, 
    41.66486, 41.69734, 41.72963, 41.76172, 41.79362, 41.82533, 41.85684, 
    41.88816, 41.91928, 41.95021, 41.98095, 42.01149, 42.04183, 42.07198, 
    42.10193, 42.13168, 42.16123, 42.19059, 42.21975, 42.24871, 42.27747, 
    42.30603, 42.33438, 42.36255, 42.39051, 42.41826, 42.44582, 42.47318, 
    42.50033, 42.52728, 42.55403, 42.58057, 42.60691, 42.63305, 42.65899, 
    42.68471, 42.71024, 42.73555, 42.76067, 42.78557, 42.81028, 42.83477, 
    42.85905, 42.88313, 42.90701, 42.93067, 42.95413, 42.97738, 43.00041, 
    43.02324, 43.04586, 43.06827, 43.09047, 43.11246, 43.13424, 43.15581, 
    43.17717, 43.19831, 43.21924, 43.23996, 43.26047, 43.28077, 43.30085, 
    43.32072, 43.34037, 43.35981, 43.37904, 43.39805, 43.41685, 43.43543, 
    43.4538, 43.47195, 43.48989, 43.50761, 43.52511, 43.5424, 43.55947, 
    43.57632, 43.59296, 43.60938, 43.62558, 43.64156, 43.65733, 43.67287, 
    43.6882, 43.70331, 43.7182, 43.73287, 43.74732, 43.76155, 43.77556, 
    43.78935, 43.80292, 43.81627, 43.8294, 43.8423, 43.85499, 43.86745, 
    43.8797, 43.89172, 43.90352, 43.9151, 43.92646, 43.93759, 43.9485, 
    43.95919, 43.96965, 43.97989, 43.98991, 43.99971, 44.00928, 44.01863, 
    44.02775, 44.03665, 44.04533, 44.05378, 44.062, 44.07001, 44.07779, 
    44.08534, 44.09267, 44.09977, 44.10666, 44.11331, 44.11974, 44.12594, 
    44.13192, 44.13767, 44.1432, 44.1485, 44.15358, 44.15842, 44.16305, 
    44.16745, 44.17162, 44.17556, 44.17928, 44.18278, 44.18604, 44.18908, 
    44.1919, 44.19448, 44.19685, 44.19898, 44.20089, 44.20257, 44.20403, 
    44.20526, 44.20626, 44.20703, 44.20758, 44.2079, 44.208, 44.20787, 
    44.20751, 44.20692, 44.20612, 44.20508, 44.20381, 44.20232, 44.2006, 
    44.19866, 44.19649, 44.19409, 44.19147, 44.18862, 44.18554, 44.18224, 
    44.17871, 44.17495, 44.17097, 44.16676, 44.16233, 44.15767, 44.15279, 
    44.14767, 44.14234, 44.13678, 44.13099, 44.12497, 44.11874, 44.11227, 
    44.10558, 44.09867, 44.09153, 44.08416, 44.07657, 44.06876, 44.06072, 
    44.05246, 44.04397, 44.03526, 44.02632, 44.01716, 44.00778, 43.99817, 
    43.98834, 43.97829, 43.96801, 43.95751, 43.94679, 43.93584, 43.92467, 
    43.91328, 43.90167, 43.88984, 43.87778, 43.8655, 43.853, 43.84028, 
    43.82734, 43.81417, 43.80079, 43.78718, 43.77336, 43.75931, 43.74505, 
    43.73056, 43.71586, 43.70093, 43.68579, 43.67043, 43.65485, 43.63905, 
    43.62303, 43.6068, 43.59034, 43.57367, 43.55679, 43.53968, 43.52236, 
    43.50482, 43.48707, 43.4691, 43.45091, 43.43251, 43.41389, 43.39506, 
    43.37601, 43.35675, 43.33728, 43.31759, 43.29769, 43.27757, 43.25724, 
    43.2367, 43.21595, 43.19498, 43.1738, 43.15241, 43.13081, 43.109, 
    43.08698, 43.06474, 43.0423, 43.01965, 42.99678, 42.97371, 42.95043, 
    42.92694, 42.90324, 42.87934, 42.85523, 42.83091, 42.80638, 42.78165, 
    42.75671, 42.73156, 42.70621, 42.68066, 42.6549, 42.62893, 42.60276, 
    42.57639, 42.54981, 42.52303, 42.49605, 42.46886, 42.44147, 42.41389, 
    42.3861, 42.3581, 42.32991, 42.30152, 42.27293, 42.24414, 42.21515, 
    42.18596, 42.15657, 42.12699, 42.0972, 42.06722, 42.03704, 42.00667, 
    41.9761, 41.94534, 41.91438, 41.88322, 41.85187, 41.82032, 41.78859, 
    41.75666, 41.72453, 41.69221, 41.65971, 41.627, 41.59411, 41.56103, 
    41.52776, 41.49429, 41.46064, 41.42679, 41.39276, 41.35854, 41.32413, 
    41.28954, 41.25475, 41.21978, 41.18462, 41.14928, 41.11375, 41.07804, 
    41.04214, 41.00606,
  37.00995, 37.06133, 37.11255, 37.16364, 37.21457, 37.26537, 37.31601, 
    37.36652, 37.41687, 37.46708, 37.51715, 37.56706, 37.61683, 37.66645, 
    37.71592, 37.76524, 37.81441, 37.86343, 37.9123, 37.96102, 38.00958, 
    38.058, 38.10626, 38.15437, 38.20233, 38.25013, 38.29778, 38.34528, 
    38.39261, 38.4398, 38.48682, 38.5337, 38.58041, 38.62696, 38.67337, 
    38.7196, 38.76569, 38.81161, 38.85738, 38.90298, 38.94842, 38.9937, 
    39.03882, 39.08378, 39.12858, 39.17321, 39.21768, 39.26199, 39.30613, 
    39.35011, 39.39392, 39.43757, 39.48106, 39.52437, 39.56752, 39.6105, 
    39.65332, 39.69596, 39.73844, 39.78075, 39.82289, 39.86486, 39.90666, 
    39.94829, 39.98975, 40.03103, 40.07215, 40.11309, 40.15385, 40.19445, 
    40.23487, 40.27512, 40.31519, 40.35509, 40.39481, 40.43436, 40.47372, 
    40.51292, 40.55193, 40.59077, 40.62943, 40.66791, 40.70621, 40.74433, 
    40.78227, 40.82003, 40.85761, 40.89501, 40.93223, 40.96926, 41.00612, 
    41.04279, 41.07927, 41.11558, 41.1517, 41.18763, 41.22338, 41.25894, 
    41.29432, 41.32951, 41.36452, 41.39933, 41.43396, 41.4684, 41.50266, 
    41.53672, 41.5706, 41.60428, 41.63778, 41.67108, 41.7042, 41.73712, 
    41.76985, 41.80239, 41.83474, 41.86689, 41.89885, 41.93062, 41.96219, 
    41.99357, 42.02475, 42.05574, 42.08653, 42.11713, 42.14753, 42.17773, 
    42.20774, 42.23755, 42.26715, 42.29657, 42.32578, 42.35479, 42.38361, 
    42.41222, 42.44064, 42.46885, 42.49686, 42.52468, 42.55229, 42.57969, 
    42.6069, 42.6339, 42.6607, 42.6873, 42.71369, 42.73988, 42.76586, 
    42.79164, 42.81721, 42.84258, 42.86774, 42.8927, 42.91745, 42.94199, 
    42.96632, 42.99045, 43.01437, 43.03808, 43.06158, 43.08488, 43.10796, 
    43.13083, 43.1535, 43.17595, 43.1982, 43.22023, 43.24205, 43.26366, 
    43.28506, 43.30625, 43.32722, 43.34798, 43.36853, 43.38887, 43.40899, 
    43.4289, 43.44859, 43.46807, 43.48734, 43.50639, 43.52523, 43.54385, 
    43.56225, 43.58044, 43.59841, 43.61617, 43.63371, 43.65103, 43.66814, 
    43.68502, 43.70169, 43.71814, 43.73438, 43.75039, 43.76619, 43.78177, 
    43.79713, 43.81227, 43.82719, 43.84188, 43.85637, 43.87062, 43.88466, 
    43.89848, 43.91208, 43.92546, 43.93861, 43.95155, 43.96426, 43.97675, 
    43.98902, 44.00106, 44.01289, 44.02449, 44.03587, 44.04703, 44.05796, 
    44.06867, 44.07915, 44.08942, 44.09946, 44.10927, 44.11887, 44.12823, 
    44.13737, 44.14629, 44.15499, 44.16346, 44.1717, 44.17972, 44.18752, 
    44.19509, 44.20243, 44.20955, 44.21644, 44.22311, 44.22955, 44.23577, 
    44.24176, 44.24752, 44.25306, 44.25837, 44.26346, 44.26832, 44.27295, 
    44.27736, 44.28154, 44.2855, 44.28922, 44.29272, 44.296, 44.29905, 
    44.30186, 44.30446, 44.30682, 44.30896, 44.31087, 44.31256, 44.31402, 
    44.31525, 44.31625, 44.31703, 44.31758, 44.31791, 44.318, 44.31787, 
    44.31751, 44.31693, 44.31611, 44.31507, 44.3138, 44.31231, 44.31059, 
    44.30864, 44.30647, 44.30406, 44.30143, 44.29858, 44.29549, 44.29218, 
    44.28865, 44.28489, 44.2809, 44.27668, 44.27224, 44.26757, 44.26267, 
    44.25755, 44.2522, 44.24663, 44.24083, 44.2348, 44.22855, 44.22207, 
    44.21537, 44.20844, 44.20128, 44.1939, 44.1863, 44.17847, 44.17041, 
    44.16213, 44.15363, 44.1449, 44.13594, 44.12677, 44.11736, 44.10773, 
    44.09789, 44.08781, 44.07751, 44.06699, 44.05624, 44.04528, 44.03408, 
    44.02267, 44.01103, 43.99918, 43.98709, 43.97479, 43.96227, 43.94952, 
    43.93655, 43.92336, 43.90994, 43.89631, 43.88246, 43.86839, 43.85409, 
    43.83957, 43.82484, 43.80989, 43.79471, 43.77932, 43.76371, 43.74788, 
    43.73183, 43.71556, 43.69907, 43.68237, 43.66544, 43.6483, 43.63095, 
    43.61337, 43.59558, 43.57758, 43.55936, 43.54092, 43.52226, 43.50339, 
    43.48431, 43.46501, 43.4455, 43.42577, 43.40582, 43.38567, 43.3653, 
    43.34472, 43.32392, 43.30291, 43.28169, 43.26026, 43.23861, 43.21676, 
    43.19469, 43.17242, 43.14993, 43.12723, 43.10432, 43.0812, 43.05788, 
    43.03434, 43.0106, 42.98665, 42.96249, 42.93812, 42.91355, 42.88876, 
    42.86378, 42.83858, 42.81318, 42.78757, 42.76176, 42.73575, 42.70953, 
    42.68311, 42.65648, 42.62965, 42.60261, 42.57537, 42.54793, 42.52029, 
    42.49245, 42.4644, 42.43616, 42.40771, 42.37907, 42.35022, 42.32117, 
    42.29193, 42.26249, 42.23284, 42.203, 42.17297, 42.14273, 42.1123, 
    42.08167, 42.05085, 42.01983, 41.98862, 41.95721, 41.92561, 41.89381, 
    41.86182, 41.82963, 41.79726, 41.76469, 41.73193, 41.69897, 41.66583, 
    41.63249, 41.59896, 41.56525, 41.53135, 41.49725, 41.46297, 41.4285, 
    41.39384, 41.35899, 41.32396, 41.28873, 41.25333, 41.21774, 41.18196, 
    41.146, 41.10985,
  37.10699, 37.15844, 37.20974, 37.26091, 37.31192, 37.36279, 37.41351, 
    37.4641, 37.51453, 37.56481, 37.61495, 37.66494, 37.71479, 37.76448, 
    37.81403, 37.86343, 37.91267, 37.96177, 38.01071, 38.05951, 38.10815, 
    38.15664, 38.20498, 38.25317, 38.3012, 38.34908, 38.3968, 38.44437, 
    38.49178, 38.53904, 38.58614, 38.63309, 38.67988, 38.72651, 38.77298, 
    38.8193, 38.86546, 38.91145, 38.95729, 39.00297, 39.04848, 39.09384, 
    39.13904, 39.18407, 39.22894, 39.27365, 39.31819, 39.36257, 39.40679, 
    39.45084, 39.49472, 39.53844, 39.582, 39.62539, 39.66861, 39.71167, 
    39.75455, 39.79727, 39.83982, 39.8822, 39.92441, 39.96645, 40.00832, 
    40.05002, 40.09155, 40.13291, 40.17409, 40.2151, 40.25594, 40.29661, 
    40.3371, 40.37741, 40.41756, 40.45752, 40.49731, 40.53693, 40.57636, 
    40.61562, 40.65471, 40.69361, 40.73234, 40.77089, 40.80926, 40.84745, 
    40.88546, 40.92328, 40.96093, 40.99839, 41.03568, 41.07278, 41.1097, 
    41.14643, 41.18299, 41.21936, 41.25554, 41.29154, 41.32735, 41.36298, 
    41.39842, 41.43368, 41.46875, 41.50362, 41.53832, 41.57282, 41.60714, 
    41.64127, 41.6752, 41.70895, 41.74251, 41.77588, 41.80905, 41.84203, 
    41.87482, 41.90742, 41.93983, 41.97205, 42.00407, 42.03589, 42.06752, 
    42.09896, 42.1302, 42.16125, 42.1921, 42.22275, 42.25321, 42.28347, 
    42.31353, 42.3434, 42.37306, 42.40253, 42.4318, 42.46087, 42.48974, 
    42.51841, 42.54688, 42.57515, 42.60321, 42.63108, 42.65874, 42.6862, 
    42.71346, 42.74051, 42.76736, 42.79401, 42.82046, 42.84669, 42.87273, 
    42.89856, 42.92418, 42.9496, 42.97481, 42.99981, 43.02461, 43.0492, 
    43.07358, 43.09776, 43.12172, 43.14548, 43.16903, 43.19237, 43.2155, 
    43.23841, 43.26113, 43.28363, 43.30591, 43.32799, 43.34985, 43.37151, 
    43.39295, 43.41418, 43.4352, 43.456, 43.47659, 43.49697, 43.51713, 
    43.53708, 43.55681, 43.57633, 43.59563, 43.61472, 43.6336, 43.65226, 
    43.6707, 43.68892, 43.70693, 43.72472, 43.7423, 43.75965, 43.77679, 
    43.79372, 43.81042, 43.8269, 43.84317, 43.85922, 43.87505, 43.89066, 
    43.90605, 43.92122, 43.93617, 43.9509, 43.96541, 43.9797, 43.99377, 
    44.00761, 44.02124, 44.03464, 44.04782, 44.06079, 44.07352, 44.08604, 
    44.09834, 44.1104, 44.12225, 44.13388, 44.14528, 44.15646, 44.16742, 
    44.17815, 44.18866, 44.19894, 44.209, 44.21884, 44.22845, 44.23783, 
    44.247, 44.25594, 44.26465, 44.27313, 44.28139, 44.28943, 44.29725, 
    44.30483, 44.31219, 44.31932, 44.32623, 44.33291, 44.33937, 44.3456, 
    44.3516, 44.35738, 44.36293, 44.36825, 44.37335, 44.37822, 44.38286, 
    44.38728, 44.39146, 44.39543, 44.39916, 44.40267, 44.40595, 44.409, 
    44.41183, 44.41443, 44.4168, 44.41895, 44.42086, 44.42255, 44.42401, 
    44.42524, 44.42625, 44.42703, 44.42758, 44.4279, 44.428, 44.42787, 
    44.42751, 44.42692, 44.42611, 44.42506, 44.42379, 44.4223, 44.42057, 
    44.41862, 44.41644, 44.41403, 44.4114, 44.40854, 44.40545, 44.40213, 
    44.39859, 44.39482, 44.39082, 44.38659, 44.38214, 44.37746, 44.37255, 
    44.36742, 44.36206, 44.35648, 44.35067, 44.34463, 44.33836, 44.33187, 
    44.32515, 44.31821, 44.31104, 44.30364, 44.29602, 44.28818, 44.28011, 
    44.2718, 44.26328, 44.25454, 44.24556, 44.23637, 44.22694, 44.2173, 
    44.20742, 44.19733, 44.18701, 44.17647, 44.1657, 44.15471, 44.14349, 
    44.13206, 44.1204, 44.10851, 44.09641, 44.08408, 44.07153, 44.05875, 
    44.04575, 44.03254, 44.0191, 44.00544, 43.99155, 43.97745, 43.96313, 
    43.94859, 43.93382, 43.91883, 43.90363, 43.8882, 43.87256, 43.8567, 
    43.84061, 43.82431, 43.80779, 43.79105, 43.7741, 43.75692, 43.73953, 
    43.72192, 43.7041, 43.68605, 43.66779, 43.64932, 43.63063, 43.61172, 
    43.59259, 43.57326, 43.5537, 43.53394, 43.51395, 43.49376, 43.47335, 
    43.45272, 43.43188, 43.41084, 43.38957, 43.3681, 43.34641, 43.32451, 
    43.3024, 43.28008, 43.25755, 43.23481, 43.21185, 43.18869, 43.16532, 
    43.14174, 43.11795, 43.09394, 43.06974, 43.04532, 43.0207, 42.99587, 
    42.97083, 42.94559, 42.92014, 42.89449, 42.86863, 42.84256, 42.81629, 
    42.78981, 42.76313, 42.73625, 42.70916, 42.68187, 42.65438, 42.62668, 
    42.59879, 42.57069, 42.54239, 42.51389, 42.48519, 42.45628, 42.42719, 
    42.39788, 42.36839, 42.33869, 42.30879, 42.2787, 42.24841, 42.21792, 
    42.18723, 42.15635, 42.12527, 42.094, 42.06253, 42.03087, 41.99901, 
    41.96696, 41.93472, 41.90228, 41.86965, 41.83683, 41.80381, 41.77061, 
    41.73721, 41.70362, 41.66985, 41.63588, 41.60172, 41.56738, 41.53284, 
    41.49812, 41.46321, 41.42811, 41.39283, 41.35736, 41.3217, 41.28586, 
    41.24983, 41.21362,
  37.204, 37.25552, 37.3069, 37.35814, 37.40923, 37.46018, 37.51098, 
    37.56164, 37.61214, 37.66251, 37.71272, 37.76279, 37.81271, 37.86248, 
    37.91211, 37.96158, 38.0109, 38.06007, 38.1091, 38.15797, 38.20668, 
    38.25525, 38.30367, 38.35193, 38.40004, 38.44799, 38.49579, 38.54343, 
    38.59092, 38.63826, 38.68544, 38.73246, 38.77932, 38.82603, 38.87257, 
    38.91896, 38.96519, 39.01127, 39.05718, 39.10293, 39.14852, 39.19395, 
    39.23922, 39.28433, 39.32927, 39.37405, 39.41867, 39.46312, 39.50741, 
    39.55154, 39.5955, 39.63929, 39.68292, 39.72638, 39.76967, 39.8128, 
    39.85576, 39.89855, 39.94117, 39.98362, 40.02591, 40.06802, 40.10996, 
    40.15173, 40.19333, 40.23476, 40.27601, 40.31709, 40.358, 40.39874, 
    40.4393, 40.47968, 40.51989, 40.55993, 40.59979, 40.63947, 40.67898, 
    40.71831, 40.75746, 40.79644, 40.83523, 40.87385, 40.91228, 40.95054, 
    40.98862, 41.02651, 41.06422, 41.10176, 41.13911, 41.17628, 41.21326, 
    41.25006, 41.28668, 41.32312, 41.35936, 41.39543, 41.4313, 41.467, 
    41.5025, 41.53782, 41.57296, 41.6079, 41.64265, 41.67722, 41.7116, 
    41.74579, 41.77979, 41.8136, 41.84722, 41.88065, 41.91389, 41.94693, 
    41.97978, 42.01244, 42.04491, 42.07718, 42.10926, 42.14115, 42.17284, 
    42.20433, 42.23564, 42.26674, 42.29765, 42.32836, 42.35888, 42.38919, 
    42.41931, 42.44923, 42.47896, 42.50848, 42.53781, 42.56693, 42.59586, 
    42.62458, 42.6531, 42.68143, 42.70955, 42.73746, 42.76518, 42.79269, 
    42.82, 42.84711, 42.87402, 42.90071, 42.92721, 42.9535, 42.97958, 
    43.00546, 43.03114, 43.0566, 43.08186, 43.10691, 43.13176, 43.1564, 
    43.18083, 43.20505, 43.22906, 43.25287, 43.27647, 43.29985, 43.32302, 
    43.34599, 43.36874, 43.39129, 43.41362, 43.43574, 43.45765, 43.47935, 
    43.50083, 43.5221, 43.54316, 43.56401, 43.58464, 43.60506, 43.62526, 
    43.64525, 43.66502, 43.68458, 43.70392, 43.72305, 43.74196, 43.76066, 
    43.77914, 43.7974, 43.81544, 43.83327, 43.85088, 43.86827, 43.88545, 
    43.9024, 43.91914, 43.93566, 43.95196, 43.96804, 43.98391, 43.99955, 
    44.01497, 44.03017, 44.04515, 44.05991, 44.07445, 44.08877, 44.10286, 
    44.11674, 44.13039, 44.14383, 44.15704, 44.17002, 44.18279, 44.19533, 
    44.20765, 44.21975, 44.23162, 44.24327, 44.25469, 44.2659, 44.27687, 
    44.28763, 44.29816, 44.30846, 44.31855, 44.3284, 44.33803, 44.34744, 
    44.35662, 44.36557, 44.37431, 44.38281, 44.39109, 44.39914, 44.40697, 
    44.41457, 44.42195, 44.4291, 44.43602, 44.44271, 44.44918, 44.45543, 
    44.46144, 44.46723, 44.47279, 44.47813, 44.48323, 44.48811, 44.49276, 
    44.49719, 44.50139, 44.50536, 44.5091, 44.51262, 44.5159, 44.51896, 
    44.5218, 44.5244, 44.52678, 44.52893, 44.53085, 44.53254, 44.534, 
    44.53524, 44.53625, 44.53703, 44.53758, 44.5379, 44.538, 44.53787, 
    44.53751, 44.53692, 44.5361, 44.53506, 44.53379, 44.53228, 44.53056, 
    44.5286, 44.52642, 44.524, 44.52136, 44.51849, 44.5154, 44.51208, 
    44.50853, 44.50475, 44.50074, 44.49651, 44.49204, 44.48735, 44.48244, 
    44.47729, 44.47192, 44.46633, 44.4605, 44.45445, 44.44817, 44.44167, 
    44.43494, 44.42798, 44.4208, 44.41338, 44.40575, 44.39788, 44.38979, 
    44.38148, 44.37294, 44.36417, 44.35518, 44.34597, 44.33652, 44.32686, 
    44.31696, 44.30685, 44.29651, 44.28594, 44.27515, 44.26414, 44.2529, 
    44.24144, 44.22976, 44.21785, 44.20572, 44.19336, 44.18078, 44.16798, 
    44.15496, 44.14172, 44.12825, 44.11456, 44.10065, 44.08652, 44.07216, 
    44.05759, 44.04279, 44.02778, 44.01254, 43.99709, 43.98141, 43.96552, 
    43.9494, 43.93306, 43.91651, 43.89974, 43.88275, 43.86554, 43.84811, 
    43.83047, 43.8126, 43.79453, 43.77623, 43.75771, 43.73899, 43.72004, 
    43.70088, 43.6815, 43.66191, 43.6421, 43.62208, 43.60184, 43.58139, 
    43.56072, 43.53984, 43.51875, 43.49745, 43.47593, 43.4542, 43.43225, 
    43.4101, 43.38774, 43.36516, 43.34237, 43.31937, 43.29617, 43.27275, 
    43.24912, 43.22528, 43.20123, 43.17698, 43.15252, 43.12785, 43.10297, 
    43.07788, 43.05259, 43.02709, 43.00138, 42.97547, 42.94936, 42.92303, 
    42.8965, 42.86977, 42.84284, 42.8157, 42.78836, 42.76081, 42.73306, 
    42.70511, 42.67696, 42.64861, 42.62005, 42.59129, 42.56234, 42.53318, 
    42.50383, 42.47427, 42.44452, 42.41456, 42.38441, 42.35406, 42.32352, 
    42.29277, 42.26183, 42.2307, 42.19937, 42.16784, 42.13612, 42.1042, 
    42.07209, 42.03979, 42.00729, 41.9746, 41.94172, 41.90864, 41.87537, 
    41.84192, 41.80827, 41.77443, 41.74039, 41.70618, 41.67177, 41.63717, 
    41.60238, 41.56741, 41.53225, 41.4969, 41.46136, 41.42564, 41.38974, 
    41.35364, 41.31736,
  37.30096, 37.35257, 37.40403, 37.45534, 37.50651, 37.55753, 37.60841, 
    37.65915, 37.70973, 37.76017, 37.81046, 37.86061, 37.9106, 37.96045, 
    38.01015, 38.0597, 38.1091, 38.15835, 38.20745, 38.25639, 38.30519, 
    38.35383, 38.40232, 38.45066, 38.49884, 38.54687, 38.59475, 38.64247, 
    38.69003, 38.73744, 38.78469, 38.83179, 38.87873, 38.92551, 38.97213, 
    39.0186, 39.0649, 39.11105, 39.15704, 39.20286, 39.24853, 39.29403, 
    39.33937, 39.38456, 39.42957, 39.47443, 39.51912, 39.56364, 39.60801, 
    39.65221, 39.69624, 39.7401, 39.78381, 39.82734, 39.8707, 39.91391, 
    39.95694, 39.9998, 40.04249, 40.08502, 40.12737, 40.16956, 40.21157, 
    40.25341, 40.29508, 40.33658, 40.37791, 40.41906, 40.46004, 40.50084, 
    40.54147, 40.58193, 40.62221, 40.66232, 40.70225, 40.742, 40.78157, 
    40.82097, 40.86019, 40.89923, 40.9381, 40.97678, 41.01529, 41.05361, 
    41.09175, 41.12972, 41.1675, 41.2051, 41.24252, 41.27975, 41.3168, 
    41.35367, 41.39035, 41.42685, 41.46317, 41.49929, 41.53524, 41.571, 
    41.60657, 41.64195, 41.67715, 41.71215, 41.74697, 41.7816, 41.81605, 
    41.8503, 41.88436, 41.91823, 41.95192, 41.9854, 42.0187, 42.05181, 
    42.08472, 42.11744, 42.14997, 42.1823, 42.21445, 42.24639, 42.27814, 
    42.3097, 42.34106, 42.37222, 42.40319, 42.43396, 42.46453, 42.4949, 
    42.52508, 42.55506, 42.58484, 42.61442, 42.6438, 42.67298, 42.70196, 
    42.73074, 42.75932, 42.78769, 42.81587, 42.84384, 42.87161, 42.89918, 
    42.92654, 42.9537, 42.98066, 43.0074, 43.03395, 43.06029, 43.08643, 
    43.11236, 43.13808, 43.1636, 43.18891, 43.21401, 43.2389, 43.26359, 
    43.28807, 43.31234, 43.3364, 43.36025, 43.38389, 43.40733, 43.43055, 
    43.45356, 43.47636, 43.49894, 43.52132, 43.54348, 43.56544, 43.58718, 
    43.6087, 43.63002, 43.65112, 43.67201, 43.69268, 43.71314, 43.73338, 
    43.75341, 43.77322, 43.79282, 43.81221, 43.83137, 43.85032, 43.86905, 
    43.88757, 43.90587, 43.92395, 43.94181, 43.95946, 43.97689, 43.9941, 
    44.01109, 44.02786, 44.04441, 44.06075, 44.07686, 44.09275, 44.10843, 
    44.12388, 44.13911, 44.15413, 44.16891, 44.18349, 44.19783, 44.21196, 
    44.22586, 44.23954, 44.25301, 44.26624, 44.27925, 44.29205, 44.30462, 
    44.31696, 44.32908, 44.34098, 44.35265, 44.3641, 44.37533, 44.38633, 
    44.39711, 44.40766, 44.41798, 44.42809, 44.43796, 44.44761, 44.45704, 
    44.46624, 44.47522, 44.48396, 44.49249, 44.50078, 44.50885, 44.5167, 
    44.52431, 44.5317, 44.53887, 44.5458, 44.55251, 44.55899, 44.56525, 
    44.57128, 44.57708, 44.58265, 44.588, 44.59312, 44.59801, 44.60267, 
    44.60711, 44.61131, 44.61529, 44.61904, 44.62256, 44.62586, 44.62893, 
    44.63176, 44.63437, 44.63675, 44.6389, 44.64083, 44.64252, 44.64399, 
    44.64523, 44.64624, 44.64703, 44.64758, 44.6479, 44.648, 44.64787, 
    44.64751, 44.64692, 44.6461, 44.64505, 44.64378, 44.64227, 44.64054, 
    44.63858, 44.63639, 44.63398, 44.63133, 44.62846, 44.62535, 44.62202, 
    44.61846, 44.61468, 44.61066, 44.60642, 44.60195, 44.59725, 44.59232, 
    44.58717, 44.58179, 44.57618, 44.57034, 44.56428, 44.55798, 44.55147, 
    44.54472, 44.53775, 44.53055, 44.52312, 44.51547, 44.50759, 44.49949, 
    44.49115, 44.48259, 44.47381, 44.4648, 44.45556, 44.4461, 44.43642, 
    44.4265, 44.41637, 44.406, 44.39542, 44.3846, 44.37357, 44.3623, 
    44.35082, 44.33911, 44.32718, 44.31502, 44.30264, 44.29004, 44.27721, 
    44.26416, 44.25089, 44.2374, 44.22368, 44.20974, 44.19558, 44.18119, 
    44.16659, 44.15176, 44.13672, 44.12145, 44.10596, 44.09026, 44.07433, 
    44.05818, 44.04181, 44.02522, 44.00842, 43.99139, 43.97415, 43.95668, 
    43.939, 43.9211, 43.90299, 43.88465, 43.8661, 43.84734, 43.82835, 
    43.80915, 43.78974, 43.7701, 43.75026, 43.73019, 43.70992, 43.68942, 
    43.66872, 43.6478, 43.62666, 43.60532, 43.58375, 43.56198, 43.53999, 
    43.5178, 43.49538, 43.47276, 43.44993, 43.42689, 43.40363, 43.38017, 
    43.35649, 43.33261, 43.30851, 43.28421, 43.2597, 43.23498, 43.21005, 
    43.18492, 43.15958, 43.13403, 43.10827, 43.08231, 43.05614, 43.02977, 
    43.00319, 42.97641, 42.94942, 42.92223, 42.89483, 42.86723, 42.83943, 
    42.81142, 42.78322, 42.75481, 42.7262, 42.69739, 42.66838, 42.63916, 
    42.60975, 42.58014, 42.55033, 42.52032, 42.49011, 42.45971, 42.4291, 
    42.3983, 42.3673, 42.33611, 42.30472, 42.27313, 42.24135, 42.20937, 
    42.1772, 42.14484, 42.11228, 42.07953, 42.04659, 42.01345, 41.98012, 
    41.9466, 41.91289, 41.87899, 41.84489, 41.81061, 41.77614, 41.74148, 
    41.70663, 41.67159, 41.63636, 41.60095, 41.56535, 41.52956, 41.49359, 
    41.45744, 41.42109,
  37.3979, 37.44958, 37.50111, 37.5525, 37.60375, 37.65485, 37.70581, 
    37.75661, 37.80728, 37.8578, 37.90816, 37.95839, 38.00846, 38.05838, 
    38.10816, 38.15779, 38.20726, 38.25659, 38.30576, 38.35479, 38.40366, 
    38.45237, 38.50094, 38.54935, 38.59761, 38.64572, 38.69367, 38.74147, 
    38.78911, 38.83659, 38.88392, 38.93109, 38.97811, 39.02496, 39.07166, 
    39.1182, 39.16458, 39.2108, 39.25686, 39.30276, 39.3485, 39.39408, 
    39.4395, 39.48475, 39.52985, 39.57478, 39.61954, 39.66414, 39.70858, 
    39.75285, 39.79696, 39.84089, 39.88467, 39.92827, 39.97171, 40.01498, 
    40.05809, 40.10102, 40.14379, 40.18639, 40.22881, 40.27107, 40.31315, 
    40.35506, 40.39681, 40.43838, 40.47977, 40.521, 40.56205, 40.60292, 
    40.64362, 40.68415, 40.7245, 40.76468, 40.80468, 40.8445, 40.88414, 
    40.92361, 40.9629, 41.00201, 41.04094, 41.0797, 41.11827, 41.15666, 
    41.19487, 41.2329, 41.27075, 41.30842, 41.3459, 41.3832, 41.42032, 
    41.45726, 41.494, 41.53057, 41.56695, 41.60315, 41.63915, 41.67497, 
    41.71061, 41.74606, 41.78132, 41.81639, 41.85127, 41.88597, 41.92048, 
    41.95479, 41.98891, 42.02285, 42.05659, 42.09015, 42.1235, 42.15667, 
    42.18965, 42.22243, 42.25502, 42.28741, 42.31961, 42.35162, 42.38343, 
    42.41504, 42.44646, 42.47768, 42.50871, 42.53954, 42.57016, 42.6006, 
    42.63083, 42.66087, 42.6907, 42.72034, 42.74977, 42.77901, 42.80805, 
    42.83688, 42.86552, 42.89395, 42.92218, 42.9502, 42.97803, 43.00565, 
    43.03306, 43.06028, 43.08728, 43.11409, 43.14068, 43.16708, 43.19326, 
    43.21924, 43.24501, 43.27058, 43.29594, 43.32109, 43.34604, 43.37077, 
    43.3953, 43.41962, 43.44373, 43.46762, 43.49131, 43.51479, 43.53806, 
    43.56111, 43.58396, 43.60659, 43.62901, 43.65122, 43.67322, 43.695, 
    43.71657, 43.73793, 43.75907, 43.78, 43.80071, 43.82121, 43.8415, 
    43.86157, 43.88142, 43.90106, 43.92048, 43.93969, 43.95868, 43.97744, 
    43.996, 44.01434, 44.03246, 44.05035, 44.06804, 44.0855, 44.10275, 
    44.11977, 44.13658, 44.15316, 44.16953, 44.18568, 44.2016, 44.21731, 
    44.23279, 44.24805, 44.2631, 44.27792, 44.29252, 44.3069, 44.32105, 
    44.33498, 44.34869, 44.36218, 44.37545, 44.38848, 44.4013, 44.4139, 
    44.42627, 44.43842, 44.45034, 44.46204, 44.47351, 44.48476, 44.49578, 
    44.50658, 44.51715, 44.5275, 44.53762, 44.54752, 44.55719, 44.56664, 
    44.57586, 44.58485, 44.59362, 44.60216, 44.61047, 44.61856, 44.62642, 
    44.63405, 44.64146, 44.64864, 44.65559, 44.66231, 44.66881, 44.67508, 
    44.68112, 44.68693, 44.69252, 44.69787, 44.703, 44.7079, 44.71257, 
    44.71702, 44.72123, 44.72522, 44.72898, 44.73251, 44.73581, 44.73888, 
    44.74173, 44.74434, 44.74673, 44.74889, 44.75082, 44.75251, 44.75399, 
    44.75523, 44.75624, 44.75702, 44.75758, 44.7579, 44.758, 44.75787, 
    44.7575, 44.75692, 44.7561, 44.75505, 44.75377, 44.75226, 44.75053, 
    44.74856, 44.74637, 44.74395, 44.74129, 44.73841, 44.73531, 44.73197, 
    44.7284, 44.72461, 44.72058, 44.71633, 44.71185, 44.70714, 44.70221, 
    44.69704, 44.69165, 44.68603, 44.68018, 44.6741, 44.6678, 44.66126, 
    44.6545, 44.64752, 44.6403, 44.63286, 44.62519, 44.61729, 44.60917, 
    44.60082, 44.59225, 44.58344, 44.57442, 44.56516, 44.55568, 44.54597, 
    44.53604, 44.52588, 44.5155, 44.50489, 44.49405, 44.48299, 44.47171, 
    44.4602, 44.44847, 44.43651, 44.42433, 44.41192, 44.39929, 44.38644, 
    44.37336, 44.36006, 44.34654, 44.33279, 44.31882, 44.30463, 44.29022, 
    44.27559, 44.26073, 44.24566, 44.23036, 44.21484, 44.1991, 44.18314, 
    44.16695, 44.15055, 44.13393, 44.11709, 44.10003, 44.08275, 44.06525, 
    44.04754, 44.0296, 44.01145, 43.99308, 43.97449, 43.95568, 43.93666, 
    43.91742, 43.89797, 43.8783, 43.85841, 43.8383, 43.81799, 43.79745, 
    43.7767, 43.75574, 43.73457, 43.71317, 43.69157, 43.66975, 43.64772, 
    43.62548, 43.60302, 43.58036, 43.55748, 43.53439, 43.51109, 43.48758, 
    43.46386, 43.43992, 43.41578, 43.39143, 43.36687, 43.34211, 43.31713, 
    43.29194, 43.26655, 43.24095, 43.21515, 43.18913, 43.16291, 43.13649, 
    43.10986, 43.08302, 43.05598, 43.02874, 43.00129, 42.97364, 42.94578, 
    42.91772, 42.88946, 42.861, 42.83234, 42.80347, 42.7744, 42.74513, 
    42.71566, 42.686, 42.65613, 42.62606, 42.5958, 42.56533, 42.53467, 
    42.50381, 42.47276, 42.4415, 42.41005, 42.37841, 42.34657, 42.31453, 
    42.2823, 42.24987, 42.21725, 42.18444, 42.15144, 42.11824, 42.08485, 
    42.05127, 42.01749, 41.98353, 41.94937, 41.91503, 41.88049, 41.84577, 
    41.81086, 41.77575, 41.74046, 41.70499, 41.66932, 41.63347, 41.59743, 
    41.56121, 41.5248,
  37.49479, 37.54655, 37.59816, 37.64963, 37.70095, 37.75213, 37.80317, 
    37.85405, 37.90479, 37.95539, 38.00583, 38.05613, 38.10628, 38.15628, 
    38.20613, 38.25584, 38.30539, 38.35479, 38.40405, 38.45314, 38.50209, 
    38.55089, 38.59953, 38.64802, 38.69635, 38.74454, 38.79256, 38.84044, 
    38.88815, 38.93571, 38.98312, 39.03036, 39.07745, 39.12439, 39.17116, 
    39.21777, 39.26423, 39.31052, 39.35666, 39.40264, 39.44845, 39.4941, 
    39.5396, 39.58492, 39.63009, 39.67509, 39.71993, 39.76461, 39.80912, 
    39.85346, 39.89764, 39.94165, 39.9855, 40.02918, 40.07269, 40.11604, 
    40.15921, 40.20222, 40.24506, 40.28773, 40.33023, 40.37255, 40.41471, 
    40.4567, 40.49851, 40.54015, 40.58162, 40.62291, 40.66403, 40.70498, 
    40.74575, 40.78635, 40.82677, 40.86702, 40.90708, 40.94698, 40.98669, 
    41.02623, 41.06559, 41.10476, 41.14376, 41.18259, 41.22123, 41.25969, 
    41.29797, 41.33606, 41.37398, 41.41171, 41.44926, 41.48663, 41.52382, 
    41.56082, 41.59763, 41.63427, 41.67071, 41.70697, 41.74305, 41.77893, 
    41.81463, 41.85014, 41.88547, 41.9206, 41.95555, 41.99031, 42.02488, 
    42.05926, 42.09345, 42.12745, 42.16125, 42.19487, 42.22829, 42.26152, 
    42.29455, 42.3274, 42.36005, 42.3925, 42.42476, 42.45683, 42.4887, 
    42.52037, 42.55185, 42.58313, 42.61421, 42.6451, 42.67579, 42.70628, 
    42.73657, 42.76666, 42.79655, 42.82625, 42.85574, 42.88503, 42.91412, 
    42.94301, 42.9717, 43.00019, 43.02847, 43.05655, 43.08443, 43.1121, 
    43.13957, 43.16684, 43.1939, 43.22075, 43.2474, 43.27385, 43.30008, 
    43.32611, 43.35194, 43.37756, 43.40297, 43.42817, 43.45316, 43.47794, 
    43.50252, 43.52688, 43.55104, 43.57499, 43.59872, 43.62225, 43.64556, 
    43.66866, 43.69155, 43.71423, 43.73669, 43.75895, 43.78099, 43.80281, 
    43.82443, 43.84583, 43.86702, 43.88799, 43.90874, 43.92928, 43.94961, 
    43.96972, 43.98961, 44.00929, 44.02875, 44.04799, 44.06702, 44.08583, 
    44.10442, 44.1228, 44.14095, 44.15889, 44.17661, 44.1941, 44.21138, 
    44.22844, 44.24529, 44.26191, 44.27831, 44.29449, 44.31044, 44.32618, 
    44.3417, 44.35699, 44.37207, 44.38692, 44.40155, 44.41595, 44.43014, 
    44.4441, 44.45784, 44.47136, 44.48465, 44.49771, 44.51056, 44.52318, 
    44.53558, 44.54774, 44.55969, 44.57141, 44.58291, 44.59418, 44.60523, 
    44.61605, 44.62665, 44.63702, 44.64716, 44.65708, 44.66677, 44.67624, 
    44.68548, 44.69449, 44.70327, 44.71183, 44.72016, 44.72827, 44.73615, 
    44.74379, 44.75121, 44.75841, 44.76537, 44.77211, 44.77862, 44.7849, 
    44.79095, 44.79678, 44.80238, 44.80775, 44.81289, 44.8178, 44.82248, 
    44.82693, 44.83116, 44.83515, 44.83892, 44.84246, 44.84576, 44.84884, 
    44.85169, 44.85431, 44.8567, 44.85887, 44.8608, 44.8625, 44.86398, 
    44.86522, 44.86623, 44.86702, 44.86758, 44.8679, 44.868, 44.86787, 
    44.8675, 44.86691, 44.86609, 44.86504, 44.86376, 44.86225, 44.86051, 
    44.85854, 44.85634, 44.85392, 44.85126, 44.84837, 44.84526, 44.84191, 
    44.83834, 44.83454, 44.83051, 44.82624, 44.82175, 44.81704, 44.81209, 
    44.80691, 44.80151, 44.79588, 44.79001, 44.78392, 44.77761, 44.77106, 
    44.76429, 44.75729, 44.75005, 44.7426, 44.73491, 44.727, 44.71886, 
    44.71049, 44.7019, 44.69308, 44.68403, 44.67476, 44.66525, 44.65553, 
    44.64557, 44.6354, 44.62499, 44.61436, 44.6035, 44.59241, 44.58111, 
    44.56958, 44.55782, 44.54583, 44.53363, 44.5212, 44.50854, 44.49566, 
    44.48256, 44.46923, 44.45568, 44.44191, 44.42791, 44.41369, 44.39925, 
    44.38458, 44.3697, 44.35459, 44.33926, 44.32371, 44.30793, 44.29194, 
    44.27573, 44.25929, 44.24264, 44.22576, 44.20866, 44.19135, 44.17382, 
    44.15606, 44.13809, 44.1199, 44.10149, 44.08287, 44.06403, 44.04496, 
    44.02568, 44.00619, 43.98648, 43.96655, 43.94641, 43.92605, 43.90547, 
    43.88468, 43.86368, 43.84246, 43.82103, 43.79938, 43.77752, 43.75544, 
    43.73315, 43.71066, 43.68794, 43.66502, 43.64188, 43.61854, 43.59498, 
    43.57121, 43.54723, 43.52304, 43.49864, 43.47404, 43.44922, 43.42419, 
    43.39896, 43.37352, 43.34787, 43.32201, 43.29595, 43.26968, 43.2432, 
    43.21652, 43.18963, 43.16254, 43.13524, 43.10774, 43.08003, 43.05212, 
    43.02401, 42.9957, 42.96718, 42.93846, 42.90953, 42.88041, 42.85109, 
    42.82156, 42.79184, 42.76191, 42.73179, 42.70147, 42.67094, 42.64022, 
    42.60931, 42.57819, 42.54688, 42.51537, 42.48367, 42.45177, 42.41967, 
    42.38738, 42.35489, 42.32221, 42.28934, 42.25627, 42.22301, 42.18956, 
    42.15591, 42.12208, 42.08805, 42.05383, 42.01942, 41.98483, 41.95004, 
    41.91506, 41.87989, 41.84454, 41.809, 41.77327, 41.73735, 41.70125, 
    41.66496, 41.62848,
  37.59166, 37.64349, 37.69518, 37.74672, 37.79813, 37.84938, 37.90049, 
    37.95145, 38.00227, 38.05294, 38.10347, 38.15384, 38.20407, 38.25415, 
    38.30408, 38.35386, 38.40348, 38.45296, 38.50229, 38.55147, 38.60049, 
    38.64936, 38.69809, 38.74665, 38.79506, 38.84332, 38.89142, 38.93937, 
    38.98716, 39.0348, 39.08228, 39.1296, 39.17677, 39.22377, 39.27062, 
    39.31731, 39.36385, 39.41022, 39.45643, 39.50248, 39.54837, 39.59409, 
    39.63966, 39.68506, 39.7303, 39.77538, 39.82029, 39.86504, 39.90963, 
    39.95404, 39.9983, 40.04239, 40.0863, 40.13006, 40.17365, 40.21706, 
    40.26031, 40.30339, 40.3463, 40.38904, 40.43161, 40.47401, 40.51624, 
    40.5583, 40.60018, 40.6419, 40.68343, 40.7248, 40.76599, 40.80701, 
    40.84785, 40.88852, 40.92901, 40.96933, 41.00946, 41.04943, 41.08921, 
    41.12882, 41.16824, 41.20749, 41.24656, 41.28545, 41.32416, 41.36269, 
    41.40104, 41.43921, 41.47719, 41.51499, 41.55261, 41.59004, 41.62729, 
    41.66436, 41.70124, 41.73794, 41.77445, 41.81078, 41.84692, 41.88287, 
    41.91864, 41.95421, 41.9896, 42.0248, 42.05981, 42.09464, 42.12927, 
    42.16371, 42.19796, 42.23202, 42.26589, 42.29957, 42.33305, 42.36634, 
    42.39944, 42.43235, 42.46506, 42.49757, 42.52989, 42.56202, 42.59395, 
    42.62568, 42.65722, 42.68856, 42.7197, 42.75065, 42.78139, 42.81194, 
    42.84229, 42.87244, 42.90239, 42.93214, 42.96169, 42.99104, 43.02019, 
    43.04913, 43.07787, 43.10641, 43.13475, 43.16289, 43.19082, 43.21855, 
    43.24607, 43.27339, 43.3005, 43.32741, 43.35411, 43.38061, 43.40689, 
    43.43298, 43.45885, 43.48452, 43.50998, 43.53523, 43.56027, 43.5851, 
    43.60973, 43.63414, 43.65834, 43.68233, 43.70612, 43.72969, 43.75305, 
    43.7762, 43.79913, 43.82186, 43.84437, 43.86667, 43.88875, 43.91062, 
    43.93228, 43.95372, 43.97495, 43.99596, 44.01676, 44.03734, 44.05771, 
    44.07786, 44.09779, 44.11751, 44.13701, 44.1563, 44.17536, 44.19421, 
    44.21284, 44.23125, 44.24944, 44.26741, 44.28517, 44.3027, 44.32002, 
    44.33711, 44.35399, 44.37064, 44.38708, 44.40329, 44.41928, 44.43505, 
    44.4506, 44.46593, 44.48103, 44.49591, 44.51057, 44.52501, 44.53922, 
    44.55322, 44.56698, 44.58052, 44.59384, 44.60694, 44.61981, 44.63245, 
    44.64488, 44.65707, 44.66904, 44.68079, 44.69231, 44.70361, 44.71468, 
    44.72552, 44.73614, 44.74653, 44.7567, 44.76664, 44.77635, 44.78584, 
    44.79509, 44.80412, 44.81293, 44.8215, 44.82985, 44.83797, 44.84587, 
    44.85353, 44.86097, 44.86818, 44.87516, 44.88191, 44.88843, 44.89473, 
    44.90079, 44.90663, 44.91224, 44.91762, 44.92277, 44.92769, 44.93238, 
    44.93684, 44.94108, 44.94508, 44.94886, 44.9524, 44.95572, 44.95881, 
    44.96166, 44.96429, 44.96668, 44.96885, 44.97078, 44.97249, 44.97397, 
    44.97522, 44.97623, 44.97702, 44.97758, 44.9779, 44.978, 44.97787, 
    44.9775, 44.97691, 44.97609, 44.97503, 44.97375, 44.97224, 44.97049, 
    44.96852, 44.96632, 44.96389, 44.96122, 44.95833, 44.95521, 44.95186, 
    44.94828, 44.94447, 44.94043, 44.93615, 44.93166, 44.92693, 44.92197, 
    44.91678, 44.91137, 44.90572, 44.89985, 44.89375, 44.88742, 44.88086, 
    44.87407, 44.86705, 44.85981, 44.85233, 44.84463, 44.8367, 44.82854, 
    44.82016, 44.81155, 44.80271, 44.79364, 44.78435, 44.77483, 44.76508, 
    44.7551, 44.7449, 44.73448, 44.72382, 44.71294, 44.70184, 44.69051, 
    44.67895, 44.66717, 44.65516, 44.64293, 44.63047, 44.61779, 44.60488, 
    44.59175, 44.5784, 44.56482, 44.55101, 44.53699, 44.52274, 44.50827, 
    44.49358, 44.47866, 44.46352, 44.44815, 44.43257, 44.41677, 44.40074, 
    44.38449, 44.36802, 44.35133, 44.33442, 44.3173, 44.29995, 44.28238, 
    44.26459, 44.24658, 44.22835, 44.2099, 44.19124, 44.17236, 44.15326, 
    44.13394, 44.11441, 44.09465, 44.07469, 44.0545, 44.0341, 44.01348, 
    43.99265, 43.97161, 43.95034, 43.92887, 43.90718, 43.88527, 43.86316, 
    43.84082, 43.81828, 43.79552, 43.77255, 43.74937, 43.72598, 43.70237, 
    43.67855, 43.65453, 43.63029, 43.60585, 43.58119, 43.55632, 43.53125, 
    43.50596, 43.48047, 43.45477, 43.42886, 43.40275, 43.37643, 43.3499, 
    43.32317, 43.29623, 43.26908, 43.24173, 43.21418, 43.18642, 43.15845, 
    43.13028, 43.10191, 43.07334, 43.04457, 43.01559, 42.98641, 42.95703, 
    42.92745, 42.89767, 42.86768, 42.83751, 42.80712, 42.77654, 42.74577, 
    42.71479, 42.68361, 42.65224, 42.62067, 42.58891, 42.55695, 42.52479, 
    42.49244, 42.4599, 42.42715, 42.39422, 42.36109, 42.32777, 42.29425, 
    42.26055, 42.22665, 42.19256, 42.15828, 42.1238, 42.08914, 42.05429, 
    42.01925, 41.98402, 41.9486, 41.91299, 41.8772, 41.84121, 41.80505, 
    41.76869, 41.73215,
  37.68848, 37.74039, 37.79216, 37.84378, 37.89526, 37.94659, 37.99778, 
    38.04882, 38.09972, 38.15046, 38.20107, 38.25152, 38.30182, 38.35198, 
    38.40199, 38.45184, 38.50154, 38.5511, 38.60051, 38.64976, 38.69886, 
    38.74781, 38.7966, 38.84525, 38.89374, 38.94207, 38.99025, 39.03827, 
    39.08614, 39.13385, 39.18141, 39.22881, 39.27605, 39.32313, 39.37006, 
    39.41682, 39.46343, 39.50988, 39.55616, 39.60229, 39.64825, 39.69405, 
    39.7397, 39.78517, 39.83049, 39.87564, 39.92063, 39.96545, 40.01011, 
    40.0546, 40.09893, 40.14309, 40.18708, 40.23091, 40.27457, 40.31806, 
    40.36138, 40.40453, 40.44751, 40.49033, 40.53297, 40.57544, 40.61774, 
    40.65987, 40.70183, 40.74361, 40.78522, 40.82666, 40.86793, 40.90902, 
    40.94993, 40.99067, 41.03123, 41.07161, 41.11182, 41.15186, 41.19171, 
    41.23138, 41.27088, 41.3102, 41.34934, 41.3883, 41.42707, 41.46567, 
    41.50409, 41.54232, 41.58037, 41.61824, 41.65593, 41.69343, 41.73075, 
    41.76788, 41.80483, 41.84159, 41.87817, 41.91457, 41.95077, 41.98679, 
    42.02262, 42.05826, 42.09372, 42.12898, 42.16405, 42.19894, 42.23364, 
    42.26814, 42.30246, 42.33658, 42.37051, 42.40425, 42.4378, 42.47115, 
    42.50431, 42.53728, 42.57005, 42.60263, 42.63501, 42.66719, 42.69918, 
    42.73098, 42.76257, 42.79397, 42.82518, 42.85618, 42.88699, 42.91759, 
    42.948, 42.97821, 43.00821, 43.03802, 43.06763, 43.09703, 43.12624, 
    43.15524, 43.18404, 43.21263, 43.24102, 43.26921, 43.2972, 43.32498, 
    43.35255, 43.37992, 43.40709, 43.43405, 43.46081, 43.48735, 43.51369, 
    43.53983, 43.56575, 43.59147, 43.61698, 43.64228, 43.66737, 43.69225, 
    43.71693, 43.74139, 43.76564, 43.78968, 43.81351, 43.83713, 43.86053, 
    43.88373, 43.90671, 43.92948, 43.95203, 43.97438, 43.99651, 44.01842, 
    44.04012, 44.06161, 44.08288, 44.10394, 44.12477, 44.1454, 44.16581, 
    44.186, 44.20597, 44.22573, 44.24527, 44.26459, 44.2837, 44.30258, 
    44.32125, 44.33969, 44.35793, 44.37594, 44.39373, 44.4113, 44.42865, 
    44.44578, 44.46269, 44.47938, 44.49585, 44.51209, 44.52811, 44.54392, 
    44.5595, 44.57486, 44.58999, 44.6049, 44.61959, 44.63406, 44.6483, 
    44.66232, 44.67612, 44.68969, 44.70304, 44.71616, 44.72906, 44.74173, 
    44.75418, 44.7664, 44.7784, 44.79017, 44.80171, 44.81303, 44.82413, 
    44.83499, 44.84563, 44.85604, 44.86623, 44.87619, 44.88593, 44.89543, 
    44.90471, 44.91376, 44.92258, 44.93117, 44.93954, 44.94768, 44.95559, 
    44.96327, 44.97072, 44.97794, 44.98494, 44.99171, 44.99824, 45.00455, 
    45.01063, 45.01648, 45.0221, 45.02749, 45.03265, 45.03759, 45.04229, 
    45.04676, 45.051, 45.05501, 45.0588, 45.06235, 45.06567, 45.06876, 
    45.07162, 45.07426, 45.07666, 45.07883, 45.08077, 45.08248, 45.08396, 
    45.08521, 45.08623, 45.08702, 45.08757, 45.0879, 45.088, 45.08787, 
    45.0875, 45.08691, 45.08608, 45.08503, 45.08374, 45.08223, 45.08048, 
    45.0785, 45.07629, 45.07386, 45.07119, 45.06829, 45.06516, 45.0618, 
    45.05821, 45.05439, 45.05035, 45.04607, 45.04156, 45.03682, 45.03185, 
    45.02665, 45.02122, 45.01557, 45.00969, 45.00357, 44.99722, 44.99065, 
    44.98385, 44.97682, 44.96956, 44.96207, 44.95435, 44.9464, 44.93823, 
    44.92983, 44.9212, 44.91234, 44.90326, 44.89394, 44.8844, 44.87463, 
    44.86464, 44.85442, 44.84396, 44.83329, 44.82239, 44.81126, 44.7999, 
    44.78832, 44.77652, 44.76448, 44.75222, 44.73974, 44.72703, 44.7141, 
    44.70094, 44.68756, 44.67395, 44.66012, 44.64606, 44.63179, 44.61729, 
    44.60256, 44.58761, 44.57244, 44.55705, 44.54143, 44.5256, 44.50954, 
    44.49326, 44.47675, 44.46003, 44.44308, 44.42592, 44.40854, 44.39093, 
    44.3731, 44.35506, 44.33679, 44.31831, 44.29961, 44.28069, 44.26155, 
    44.24219, 44.22262, 44.20283, 44.18282, 44.16259, 44.14215, 44.12149, 
    44.10062, 44.07953, 44.05822, 44.03671, 44.01497, 43.99302, 43.97086, 
    43.94848, 43.92589, 43.90309, 43.88007, 43.85685, 43.8334, 43.80975, 
    43.78589, 43.76182, 43.73753, 43.71304, 43.68833, 43.66341, 43.63829, 
    43.61296, 43.58742, 43.56166, 43.53571, 43.50954, 43.48317, 43.45659, 
    43.4298, 43.40281, 43.37561, 43.34821, 43.3206, 43.29279, 43.26477, 
    43.23655, 43.20812, 43.17949, 43.15066, 43.12163, 43.09239, 43.06296, 
    43.03332, 43.00348, 42.97344, 42.9432, 42.91276, 42.88213, 42.85129, 
    42.82025, 42.78902, 42.75759, 42.72596, 42.69414, 42.66212, 42.6299, 
    42.59749, 42.56488, 42.53208, 42.49908, 42.46589, 42.43251, 42.39893, 
    42.36516, 42.3312, 42.29704, 42.2627, 42.22816, 42.19344, 42.15852, 
    42.12341, 42.08812, 42.05264, 42.01696, 41.9811, 41.94506, 41.90882, 
    41.8724, 41.83579,
  37.78526, 37.83725, 37.8891, 37.9408, 37.99236, 38.04377, 38.09503, 
    38.14615, 38.19712, 38.24795, 38.29863, 38.34916, 38.39954, 38.44977, 
    38.49986, 38.54979, 38.59957, 38.6492, 38.69869, 38.74802, 38.7972, 
    38.84622, 38.89509, 38.94381, 38.99238, 39.04079, 39.08904, 39.13714, 
    39.18509, 39.23288, 39.28051, 39.32798, 39.3753, 39.42246, 39.46946, 
    39.5163, 39.56298, 39.6095, 39.65587, 39.70207, 39.74811, 39.79398, 
    39.8397, 39.88525, 39.93064, 39.97587, 40.02093, 40.06583, 40.11056, 
    40.15512, 40.19953, 40.24376, 40.28783, 40.33173, 40.37546, 40.41903, 
    40.46242, 40.50565, 40.5487, 40.59159, 40.6343, 40.67685, 40.71922, 
    40.76143, 40.80345, 40.84531, 40.88699, 40.9285, 40.96983, 41.01099, 
    41.05198, 41.09279, 41.13342, 41.17388, 41.21416, 41.25426, 41.29418, 
    41.33393, 41.37349, 41.41288, 41.45209, 41.49112, 41.52996, 41.56863, 
    41.60711, 41.64542, 41.68354, 41.72147, 41.75923, 41.79679, 41.83418, 
    41.87138, 41.9084, 41.94523, 41.98187, 42.01833, 42.0546, 42.09069, 
    42.12658, 42.16229, 42.19781, 42.23314, 42.26828, 42.30323, 42.33799, 
    42.37256, 42.40694, 42.44112, 42.47512, 42.50892, 42.54253, 42.57594, 
    42.60917, 42.64219, 42.67503, 42.70766, 42.74011, 42.77235, 42.80441, 
    42.83626, 42.86791, 42.89937, 42.93063, 42.9617, 42.99256, 43.02322, 
    43.05369, 43.08395, 43.11402, 43.14388, 43.17355, 43.20301, 43.23227, 
    43.26133, 43.29018, 43.31883, 43.34728, 43.37552, 43.40356, 43.4314, 
    43.45903, 43.48645, 43.51367, 43.54068, 43.56749, 43.59409, 43.62048, 
    43.64667, 43.67264, 43.69841, 43.72397, 43.74932, 43.77446, 43.79939, 
    43.82411, 43.84863, 43.87292, 43.89701, 43.92089, 43.94456, 43.96801, 
    43.99125, 44.01428, 44.03709, 44.05969, 44.08208, 44.10426, 44.12621, 
    44.14796, 44.16949, 44.1908, 44.2119, 44.23278, 44.25344, 44.2739, 
    44.29412, 44.31414, 44.33394, 44.35352, 44.37288, 44.39202, 44.41095, 
    44.42965, 44.44814, 44.46641, 44.48445, 44.50228, 44.51989, 44.53727, 
    44.55444, 44.57138, 44.5881, 44.60461, 44.62089, 44.63694, 44.65278, 
    44.66839, 44.68378, 44.69895, 44.71389, 44.72861, 44.74311, 44.75738, 
    44.77143, 44.78526, 44.79885, 44.81223, 44.82538, 44.8383, 44.851, 
    44.86348, 44.87572, 44.88774, 44.89954, 44.91111, 44.92245, 44.93357, 
    44.94446, 44.95512, 44.96556, 44.97577, 44.98574, 44.9955, 45.00502, 
    45.01432, 45.02339, 45.03223, 45.04084, 45.04922, 45.05738, 45.06531, 
    45.07301, 45.08047, 45.08771, 45.09472, 45.1015, 45.10806, 45.11438, 
    45.12047, 45.12633, 45.13196, 45.13736, 45.14254, 45.14748, 45.15219, 
    45.15667, 45.16092, 45.16494, 45.16874, 45.17229, 45.17562, 45.17872, 
    45.18159, 45.18423, 45.18663, 45.18881, 45.19075, 45.19247, 45.19395, 
    45.1952, 45.19622, 45.19701, 45.19757, 45.1979, 45.198, 45.19786, 
    45.1975, 45.1969, 45.19608, 45.19502, 45.19373, 45.19221, 45.19046, 
    45.18848, 45.18627, 45.18383, 45.18115, 45.17825, 45.17511, 45.17175, 
    45.16815, 45.16432, 45.16027, 45.15598, 45.15146, 45.14671, 45.14173, 
    45.13652, 45.13108, 45.12542, 45.11952, 45.11339, 45.10703, 45.10044, 
    45.09363, 45.08658, 45.07931, 45.0718, 45.06407, 45.05611, 45.04792, 
    45.03949, 45.03085, 45.02197, 45.01286, 45.00353, 44.99397, 44.98418, 
    44.97417, 44.96392, 44.95345, 44.94275, 44.93183, 44.92067, 44.9093, 
    44.89769, 44.88586, 44.8738, 44.86152, 44.84901, 44.83627, 44.82331, 
    44.81013, 44.79672, 44.78308, 44.76922, 44.75514, 44.74083, 44.7263, 
    44.71154, 44.69656, 44.68136, 44.66594, 44.65029, 44.63442, 44.61833, 
    44.60201, 44.58548, 44.56872, 44.55174, 44.53454, 44.51712, 44.49947, 
    44.48161, 44.46353, 44.44523, 44.42671, 44.40797, 44.38901, 44.36983, 
    44.35044, 44.33082, 44.31099, 44.29094, 44.27068, 44.25019, 44.22949, 
    44.20858, 44.18744, 44.1661, 44.14453, 44.12275, 44.10076, 44.07855, 
    44.05613, 44.0335, 44.01065, 43.98759, 43.96431, 43.94083, 43.91713, 
    43.89322, 43.86909, 43.84476, 43.82022, 43.79546, 43.7705, 43.74532, 
    43.71994, 43.69435, 43.66855, 43.64254, 43.61632, 43.5899, 43.56326, 
    43.53643, 43.50938, 43.48213, 43.45467, 43.42701, 43.39914, 43.37107, 
    43.34279, 43.31431, 43.28563, 43.25674, 43.22765, 43.19836, 43.16887, 
    43.13918, 43.10928, 43.07918, 43.04889, 43.01839, 42.98769, 42.95679, 
    42.9257, 42.89441, 42.86292, 42.83123, 42.79935, 42.76727, 42.73499, 
    42.70251, 42.66985, 42.63698, 42.60392, 42.57067, 42.53722, 42.50359, 
    42.46975, 42.43573, 42.40151, 42.3671, 42.3325, 42.29771, 42.26273, 
    42.22756, 42.1922, 42.15665, 42.12091, 42.08499, 42.04888, 42.01258, 
    41.97609, 41.93941,
  37.88202, 37.93408, 37.986, 38.03778, 38.08942, 38.14091, 38.19225, 
    38.24345, 38.29449, 38.3454, 38.39616, 38.44676, 38.49722, 38.54753, 
    38.59769, 38.64771, 38.69756, 38.74727, 38.79683, 38.84624, 38.8955, 
    38.9446, 38.99355, 39.04234, 39.09098, 39.13947, 39.18781, 39.23598, 
    39.284, 39.33187, 39.37957, 39.42712, 39.47452, 39.52176, 39.56883, 
    39.61575, 39.66251, 39.7091, 39.75554, 39.80182, 39.84793, 39.89388, 
    39.93967, 39.9853, 40.03077, 40.07607, 40.1212, 40.16618, 40.21098, 
    40.25562, 40.3001, 40.34441, 40.38855, 40.43252, 40.47633, 40.51997, 
    40.56343, 40.60673, 40.64986, 40.69282, 40.73561, 40.77822, 40.82067, 
    40.86295, 40.90505, 40.94698, 40.98873, 41.03031, 41.07172, 41.11295, 
    41.154, 41.19488, 41.23559, 41.27612, 41.31646, 41.35664, 41.39663, 
    41.43645, 41.47608, 41.51554, 41.55482, 41.59391, 41.63283, 41.67156, 
    41.71012, 41.74849, 41.78667, 41.82468, 41.8625, 41.90014, 41.93759, 
    41.97486, 42.01194, 42.04884, 42.08555, 42.12207, 42.15841, 42.19456, 
    42.23052, 42.2663, 42.30188, 42.33728, 42.37248, 42.4075, 42.44232, 
    42.47696, 42.51139, 42.54565, 42.5797, 42.61357, 42.64724, 42.68072, 
    42.714, 42.74709, 42.77999, 42.81268, 42.84519, 42.87749, 42.90961, 
    42.94152, 42.97324, 43.00476, 43.03608, 43.0672, 43.09812, 43.12885, 
    43.15937, 43.18969, 43.21981, 43.24973, 43.27945, 43.30897, 43.33829, 
    43.3674, 43.39631, 43.42502, 43.45352, 43.48182, 43.50991, 43.5378, 
    43.56549, 43.59297, 43.62024, 43.6473, 43.67416, 43.70081, 43.72726, 
    43.75349, 43.77952, 43.80534, 43.83095, 43.85635, 43.88154, 43.90652, 
    43.93129, 43.95585, 43.9802, 44.00434, 44.02826, 44.05198, 44.07547, 
    44.09876, 44.12183, 44.1447, 44.16734, 44.18977, 44.21199, 44.234, 
    44.25578, 44.27736, 44.29871, 44.31985, 44.34078, 44.36148, 44.38198, 
    44.40225, 44.42231, 44.44214, 44.46176, 44.48116, 44.50034, 44.51931, 
    44.53805, 44.55658, 44.57488, 44.59296, 44.61083, 44.62847, 44.64589, 
    44.66309, 44.68007, 44.69683, 44.71336, 44.72968, 44.74577, 44.76164, 
    44.77728, 44.79271, 44.8079, 44.82288, 44.83763, 44.85215, 44.86646, 
    44.88054, 44.89439, 44.90802, 44.92142, 44.93459, 44.94755, 44.96027, 
    44.97277, 44.98505, 44.99709, 45.00891, 45.02051, 45.03187, 45.04301, 
    45.05392, 45.06461, 45.07507, 45.0853, 45.0953, 45.10507, 45.11462, 
    45.12393, 45.13302, 45.14188, 45.15051, 45.15891, 45.16708, 45.17503, 
    45.18274, 45.19022, 45.19748, 45.2045, 45.2113, 45.21786, 45.2242, 
    45.2303, 45.23618, 45.24182, 45.24723, 45.25242, 45.25737, 45.26209, 
    45.26658, 45.27084, 45.27487, 45.27867, 45.28224, 45.28558, 45.28868, 
    45.29155, 45.2942, 45.29661, 45.29879, 45.30074, 45.30246, 45.30394, 
    45.3052, 45.30622, 45.30701, 45.30757, 45.3079, 45.308, 45.30787, 
    45.3075, 45.3069, 45.30608, 45.30502, 45.30372, 45.3022, 45.30045, 
    45.29846, 45.29624, 45.2938, 45.29111, 45.2882, 45.28506, 45.28169, 
    45.27809, 45.27425, 45.27019, 45.26589, 45.26136, 45.2566, 45.25161, 
    45.2464, 45.24094, 45.23526, 45.22935, 45.22321, 45.21684, 45.21024, 
    45.20341, 45.19635, 45.18906, 45.18153, 45.17379, 45.16581, 45.1576, 
    45.14916, 45.14049, 45.1316, 45.12247, 45.11312, 45.10354, 45.09373, 
    45.08369, 45.07343, 45.06293, 45.05222, 45.04126, 45.03009, 45.01869, 
    45.00706, 44.9952, 44.98312, 44.97081, 44.95827, 44.94551, 44.93253, 
    44.91931, 44.90587, 44.89221, 44.87832, 44.86421, 44.84987, 44.83531, 
    44.82052, 44.80551, 44.79028, 44.77482, 44.75914, 44.74324, 44.72711, 
    44.71077, 44.69419, 44.6774, 44.66039, 44.64315, 44.62569, 44.60802, 
    44.59012, 44.572, 44.55366, 44.5351, 44.51632, 44.49733, 44.47811, 
    44.45867, 44.43902, 44.41915, 44.39906, 44.37875, 44.35822, 44.33748, 
    44.31652, 44.29535, 44.27396, 44.25235, 44.23053, 44.20849, 44.18624, 
    44.16377, 44.14109, 44.1182, 44.09509, 44.07177, 44.04824, 44.02449, 
    44.00053, 43.97636, 43.95198, 43.92739, 43.90258, 43.87757, 43.85235, 
    43.82691, 43.80127, 43.77542, 43.74936, 43.72309, 43.69661, 43.66993, 
    43.64304, 43.61594, 43.58863, 43.56112, 43.53341, 43.50549, 43.47736, 
    43.44903, 43.42049, 43.39175, 43.36281, 43.33366, 43.30432, 43.27477, 
    43.24501, 43.21506, 43.18491, 43.15455, 43.124, 43.09324, 43.06229, 
    43.03114, 42.99978, 42.96824, 42.93649, 42.90454, 42.8724, 42.84006, 
    42.80753, 42.7748, 42.74187, 42.70875, 42.67543, 42.64193, 42.60822, 
    42.57433, 42.54024, 42.50596, 42.47149, 42.43682, 42.40197, 42.36692, 
    42.33169, 42.29626, 42.26065, 42.22485, 42.18886, 42.15268, 42.11631, 
    42.07976, 42.04301,
  37.97873, 38.03087, 38.08287, 38.13473, 38.18644, 38.23801, 38.28943, 
    38.3407, 38.39183, 38.44281, 38.49364, 38.54433, 38.59487, 38.64526, 
    38.6955, 38.74558, 38.79552, 38.84531, 38.89494, 38.94443, 38.99376, 
    39.04294, 39.09196, 39.14084, 39.18956, 39.23812, 39.28653, 39.33479, 
    39.38288, 39.43082, 39.47861, 39.52623, 39.5737, 39.62102, 39.66817, 
    39.71516, 39.76199, 39.80867, 39.85518, 39.90153, 39.94772, 39.99375, 
    40.03962, 40.08532, 40.13086, 40.17624, 40.22145, 40.26649, 40.31137, 
    40.35609, 40.40064, 40.44502, 40.48923, 40.53328, 40.57716, 40.62088, 
    40.66442, 40.70779, 40.75099, 40.79403, 40.83689, 40.87958, 40.9221, 
    40.96444, 41.00661, 41.04861, 41.09044, 41.1321, 41.17357, 41.21487, 
    41.256, 41.29695, 41.33773, 41.37833, 41.41875, 41.45899, 41.49905, 
    41.53894, 41.57865, 41.61817, 41.65752, 41.69669, 41.73567, 41.77448, 
    41.8131, 41.85154, 41.88979, 41.92786, 41.96576, 42.00346, 42.04098, 
    42.07832, 42.11547, 42.15243, 42.18921, 42.2258, 42.2622, 42.29842, 
    42.33445, 42.37029, 42.40593, 42.44139, 42.47666, 42.51174, 42.54663, 
    42.58133, 42.61583, 42.65015, 42.68427, 42.7182, 42.75193, 42.78547, 
    42.81882, 42.85197, 42.88493, 42.91769, 42.95025, 42.98262, 43.01479, 
    43.04677, 43.07854, 43.11012, 43.1415, 43.17268, 43.20367, 43.23445, 
    43.26503, 43.29541, 43.32559, 43.35557, 43.38535, 43.41492, 43.44429, 
    43.47346, 43.50243, 43.53119, 43.55975, 43.5881, 43.61625, 43.6442, 
    43.67194, 43.69947, 43.72679, 43.75391, 43.78082, 43.80753, 43.83402, 
    43.86031, 43.88639, 43.91226, 43.93792, 43.96337, 43.98861, 44.01364, 
    44.03846, 44.06307, 44.08747, 44.11165, 44.13562, 44.15938, 44.18293, 
    44.20626, 44.22939, 44.25229, 44.27498, 44.29746, 44.31972, 44.34177, 
    44.3636, 44.38522, 44.40662, 44.4278, 44.44877, 44.46952, 44.49005, 
    44.51036, 44.53046, 44.55034, 44.57, 44.58944, 44.60866, 44.62766, 
    44.64644, 44.665, 44.68335, 44.70147, 44.71937, 44.73705, 44.75451, 
    44.77174, 44.78876, 44.80555, 44.82212, 44.83847, 44.85459, 44.87049, 
    44.88617, 44.90162, 44.91685, 44.93186, 44.94664, 44.9612, 44.97553, 
    44.98964, 45.00352, 45.01717, 45.0306, 45.04381, 45.05679, 45.06954, 
    45.08207, 45.09436, 45.10643, 45.11828, 45.1299, 45.14129, 45.15245, 
    45.16339, 45.1741, 45.18457, 45.19482, 45.20485, 45.21464, 45.22421, 
    45.23354, 45.24265, 45.25153, 45.26017, 45.26859, 45.27678, 45.28474, 
    45.29247, 45.29997, 45.30724, 45.31428, 45.32109, 45.32767, 45.33402, 
    45.34014, 45.34602, 45.35168, 45.35711, 45.3623, 45.36726, 45.37199, 
    45.3765, 45.38076, 45.3848, 45.38861, 45.39219, 45.39553, 45.39864, 
    45.40152, 45.40417, 45.40659, 45.40877, 45.41072, 45.41245, 45.41393, 
    45.41519, 45.41622, 45.41701, 45.41757, 45.4179, 45.418, 45.41787, 
    45.4175, 45.4169, 45.41607, 45.41501, 45.41372, 45.41219, 45.41043, 
    45.40844, 45.40622, 45.40377, 45.40108, 45.39816, 45.39502, 45.39164, 
    45.38802, 45.38418, 45.3801, 45.3758, 45.37126, 45.36649, 45.36149, 
    45.35626, 45.3508, 45.34511, 45.33918, 45.33303, 45.32664, 45.32003, 
    45.31319, 45.30611, 45.2988, 45.29127, 45.2835, 45.27551, 45.26728, 
    45.25882, 45.25014, 45.24122, 45.23208, 45.22271, 45.21311, 45.20328, 
    45.19322, 45.18293, 45.17242, 45.16167, 45.1507, 45.1395, 45.12807, 
    45.11642, 45.10454, 45.09243, 45.0801, 45.06754, 45.05475, 45.04173, 
    45.02849, 45.01503, 45.00134, 44.98742, 44.97327, 44.95891, 44.94432, 
    44.9295, 44.91446, 44.89919, 44.8837, 44.86799, 44.85205, 44.8359, 
    44.81951, 44.80291, 44.78608, 44.76903, 44.75176, 44.73427, 44.71655, 
    44.69862, 44.68046, 44.66209, 44.64349, 44.62467, 44.60563, 44.58638, 
    44.5669, 44.54721, 44.5273, 44.50716, 44.48682, 44.46625, 44.44547, 
    44.42447, 44.40325, 44.38181, 44.36016, 44.3383, 44.31622, 44.29392, 
    44.27141, 44.24868, 44.22574, 44.20259, 44.17922, 44.15564, 44.13184, 
    44.10784, 44.08362, 44.05919, 44.03455, 44.0097, 43.98463, 43.95936, 
    43.93388, 43.90818, 43.88228, 43.85617, 43.82985, 43.80332, 43.77658, 
    43.74963, 43.72248, 43.69513, 43.66756, 43.63979, 43.61182, 43.58363, 
    43.55525, 43.52666, 43.49786, 43.46886, 43.43966, 43.41026, 43.38065, 
    43.35084, 43.32083, 43.29062, 43.2602, 43.22959, 43.19878, 43.16776, 
    43.13655, 43.10514, 43.07353, 43.04172, 43.00972, 42.97752, 42.94511, 
    42.91252, 42.87973, 42.84674, 42.81356, 42.78018, 42.74661, 42.71284, 
    42.67889, 42.64473, 42.61039, 42.57586, 42.54113, 42.50621, 42.4711, 
    42.4358, 42.40031, 42.36463, 42.32876, 42.2927, 42.25645, 42.22002, 
    42.1834, 42.1466,
  38.0754, 38.12762, 38.1797, 38.23164, 38.28343, 38.33507, 38.38657, 
    38.43792, 38.48913, 38.54019, 38.5911, 38.64186, 38.69248, 38.74294, 
    38.79326, 38.84343, 38.89344, 38.94331, 38.99302, 39.04258, 39.09199, 
    39.14125, 39.19035, 39.2393, 39.2881, 39.33674, 39.38522, 39.43356, 
    39.48173, 39.52975, 39.57761, 39.62531, 39.67286, 39.72025, 39.76748, 
    39.81454, 39.86145, 39.9082, 39.95479, 40.00122, 40.04749, 40.09359, 
    40.13953, 40.18531, 40.23092, 40.27637, 40.32166, 40.36678, 40.41174, 
    40.45653, 40.50115, 40.54561, 40.5899, 40.63402, 40.67797, 40.72176, 
    40.76537, 40.80882, 40.8521, 40.8952, 40.93814, 40.9809, 41.02349, 
    41.06591, 41.10815, 41.15023, 41.19213, 41.23385, 41.2754, 41.31678, 
    41.35798, 41.399, 41.43984, 41.48051, 41.521, 41.56132, 41.60145, 
    41.64141, 41.68119, 41.72078, 41.7602, 41.79943, 41.83849, 41.87736, 
    41.91605, 41.95456, 41.99289, 42.03103, 42.06898, 42.10676, 42.14435, 
    42.18175, 42.21897, 42.256, 42.29284, 42.3295, 42.36597, 42.40225, 
    42.43835, 42.47425, 42.50996, 42.54549, 42.58083, 42.61597, 42.65092, 
    42.68568, 42.72026, 42.75463, 42.78882, 42.82281, 42.85661, 42.89021, 
    42.92362, 42.95683, 42.98985, 43.02267, 43.0553, 43.08773, 43.11996, 
    43.152, 43.18383, 43.21547, 43.24691, 43.27815, 43.30919, 43.34003, 
    43.37067, 43.40112, 43.43135, 43.46139, 43.49123, 43.52085, 43.55029, 
    43.57951, 43.60854, 43.63735, 43.66597, 43.69437, 43.72258, 43.75058, 
    43.77837, 43.80595, 43.83334, 43.86051, 43.88747, 43.91423, 43.94078, 
    43.96711, 43.99324, 44.01917, 44.04488, 44.07038, 44.09567, 44.12075, 
    44.14562, 44.17028, 44.19472, 44.21895, 44.24297, 44.26678, 44.29037, 
    44.31376, 44.33693, 44.35987, 44.38261, 44.40514, 44.42744, 44.44954, 
    44.47141, 44.49307, 44.51451, 44.53574, 44.55675, 44.57754, 44.59812, 
    44.61847, 44.63861, 44.65853, 44.67823, 44.69771, 44.71697, 44.73601, 
    44.75483, 44.77343, 44.79181, 44.80997, 44.82791, 44.84562, 44.86312, 
    44.88039, 44.89744, 44.91426, 44.93087, 44.94725, 44.96341, 44.97934, 
    44.99505, 45.01054, 45.02579, 45.04083, 45.05564, 45.07023, 45.08459, 
    45.09873, 45.11264, 45.12633, 45.13979, 45.15302, 45.16602, 45.1788, 
    45.19135, 45.20368, 45.21578, 45.22765, 45.23929, 45.2507, 45.26189, 
    45.27285, 45.28358, 45.29408, 45.30435, 45.3144, 45.32421, 45.33379, 
    45.34315, 45.35228, 45.36118, 45.36984, 45.37828, 45.38649, 45.39446, 
    45.40221, 45.40972, 45.41701, 45.42406, 45.43089, 45.43748, 45.44384, 
    45.44997, 45.45587, 45.46154, 45.46698, 45.47218, 45.47715, 45.4819, 
    45.48641, 45.49068, 45.49473, 45.49855, 45.50213, 45.50548, 45.5086, 
    45.51149, 45.51414, 45.51656, 45.51875, 45.52071, 45.52243, 45.52393, 
    45.52518, 45.52621, 45.52701, 45.52757, 45.5279, 45.528, 45.52787, 
    45.5275, 45.5269, 45.52607, 45.525, 45.5237, 45.52217, 45.52041, 
    45.51842, 45.51619, 45.51373, 45.51104, 45.50812, 45.50497, 45.50158, 
    45.49796, 45.49411, 45.49002, 45.48571, 45.48116, 45.47638, 45.47137, 
    45.46613, 45.46066, 45.45495, 45.44902, 45.44285, 45.43645, 45.42982, 
    45.42296, 45.41587, 45.40855, 45.401, 45.39322, 45.3852, 45.37696, 
    45.36848, 45.35978, 45.35085, 45.34169, 45.33229, 45.32267, 45.31282, 
    45.30274, 45.29243, 45.28189, 45.27113, 45.26014, 45.24891, 45.23746, 
    45.22578, 45.21388, 45.20174, 45.18938, 45.1768, 45.16398, 45.15094, 
    45.13767, 45.12418, 45.11045, 45.09651, 45.08234, 45.06794, 45.05332, 
    45.03847, 45.0234, 45.0081, 44.99258, 44.97683, 44.96087, 44.94467, 
    44.92826, 44.91162, 44.89476, 44.87767, 44.86036, 44.84283, 44.82508, 
    44.80711, 44.78892, 44.7705, 44.75187, 44.73301, 44.71394, 44.69464, 
    44.67513, 44.65539, 44.63544, 44.61527, 44.59488, 44.57427, 44.55344, 
    44.5324, 44.51114, 44.48966, 44.46797, 44.44606, 44.42393, 44.40159, 
    44.37903, 44.35626, 44.33327, 44.31007, 44.28666, 44.26303, 44.23919, 
    44.21513, 44.19087, 44.16639, 44.1417, 44.11679, 44.09168, 44.06636, 
    44.04082, 44.01508, 43.98912, 43.96296, 43.93659, 43.91001, 43.88322, 
    43.85622, 43.82902, 43.80161, 43.77399, 43.74616, 43.71813, 43.6899, 
    43.66145, 43.63281, 43.60396, 43.5749, 43.54564, 43.51618, 43.48652, 
    43.45665, 43.42658, 43.39631, 43.36584, 43.33517, 43.3043, 43.27322, 
    43.24195, 43.21048, 43.17881, 43.14694, 43.11488, 43.08261, 43.05015, 
    43.01749, 42.98464, 42.95159, 42.91835, 42.88491, 42.85127, 42.81744, 
    42.78342, 42.74921, 42.7148, 42.6802, 42.64541, 42.61042, 42.57525, 
    42.53988, 42.50433, 42.46858, 42.43265, 42.39653, 42.36021, 42.32372, 
    42.28703, 42.25015,
  38.17204, 38.22434, 38.2765, 38.32851, 38.38038, 38.4321, 38.48368, 
    38.53511, 38.5864, 38.63753, 38.68852, 38.73936, 38.79005, 38.8406, 
    38.89099, 38.94123, 38.99133, 39.04127, 39.09106, 39.1407, 39.19019, 
    39.23952, 39.2887, 39.33773, 39.3866, 39.43532, 39.48388, 39.53229, 
    39.58054, 39.62864, 39.67657, 39.72435, 39.77198, 39.81944, 39.86674, 
    39.91389, 39.96088, 40.0077, 40.05437, 40.10087, 40.14721, 40.19339, 
    40.23941, 40.28526, 40.33096, 40.37648, 40.42184, 40.46704, 40.51207, 
    40.55693, 40.60163, 40.64616, 40.69053, 40.73472, 40.77875, 40.82261, 
    40.8663, 40.90982, 40.95317, 40.99635, 41.03936, 41.0822, 41.12486, 
    41.16735, 41.20967, 41.25182, 41.29379, 41.33558, 41.3772, 41.41865, 
    41.45992, 41.50101, 41.54193, 41.58267, 41.62324, 41.66362, 41.70383, 
    41.74385, 41.7837, 41.82337, 41.86285, 41.90216, 41.94128, 41.98022, 
    42.01899, 42.05756, 42.09596, 42.13417, 42.1722, 42.21003, 42.24769, 
    42.28516, 42.32245, 42.35955, 42.39646, 42.43318, 42.46972, 42.50607, 
    42.54222, 42.5782, 42.61398, 42.64957, 42.68497, 42.72018, 42.7552, 
    42.79002, 42.82466, 42.8591, 42.89334, 42.9274, 42.96126, 42.99493, 
    43.0284, 43.06168, 43.09476, 43.12764, 43.16033, 43.19282, 43.22511, 
    43.25721, 43.28911, 43.32081, 43.35231, 43.38361, 43.41471, 43.44561, 
    43.47631, 43.50681, 43.5371, 43.5672, 43.59709, 43.62678, 43.65626, 
    43.68555, 43.71463, 43.7435, 43.77217, 43.80063, 43.82889, 43.85695, 
    43.88479, 43.91243, 43.93987, 43.96709, 43.99411, 44.02092, 44.04752, 
    44.07391, 44.10009, 44.12606, 44.15182, 44.17738, 44.20272, 44.22785, 
    44.25277, 44.27747, 44.30197, 44.32625, 44.35032, 44.37417, 44.39781, 
    44.42124, 44.44445, 44.46745, 44.49024, 44.51281, 44.53516, 44.55729, 
    44.57922, 44.60092, 44.62241, 44.64367, 44.66473, 44.68556, 44.70618, 
    44.72657, 44.74675, 44.76671, 44.78645, 44.80597, 44.82527, 44.84435, 
    44.86321, 44.88185, 44.90027, 44.91846, 44.93644, 44.95419, 44.97172, 
    44.98903, 45.00611, 45.02297, 45.03961, 45.05603, 45.07222, 45.08818, 
    45.10393, 45.11945, 45.13474, 45.14981, 45.16465, 45.17927, 45.19366, 
    45.20782, 45.22176, 45.23548, 45.24896, 45.26222, 45.27526, 45.28806, 
    45.30064, 45.31299, 45.32512, 45.33701, 45.34868, 45.36012, 45.37133, 
    45.38231, 45.39306, 45.40358, 45.41388, 45.42394, 45.43378, 45.44338, 
    45.45276, 45.4619, 45.47082, 45.4795, 45.48796, 45.49618, 45.50418, 
    45.51194, 45.51947, 45.52677, 45.53384, 45.54068, 45.54729, 45.55366, 
    45.55981, 45.56572, 45.5714, 45.57685, 45.58206, 45.58705, 45.5918, 
    45.59632, 45.60061, 45.60466, 45.60848, 45.61208, 45.61543, 45.61856, 
    45.62145, 45.62411, 45.62654, 45.62873, 45.63069, 45.63242, 45.63391, 
    45.63518, 45.63621, 45.637, 45.63757, 45.6379, 45.638, 45.63786, 45.6375, 
    45.63689, 45.63606, 45.63499, 45.63369, 45.63216, 45.6304, 45.6284, 
    45.62617, 45.6237, 45.62101, 45.61808, 45.61492, 45.61152, 45.60789, 
    45.60403, 45.59995, 45.59562, 45.59106, 45.58627, 45.58125, 45.576, 
    45.57051, 45.5648, 45.55885, 45.55267, 45.54626, 45.53961, 45.53274, 
    45.52563, 45.5183, 45.51073, 45.50293, 45.4949, 45.48664, 45.47815, 
    45.46943, 45.46047, 45.45129, 45.44188, 45.43224, 45.42236, 45.41226, 
    45.40193, 45.39137, 45.38058, 45.36957, 45.35832, 45.34685, 45.33514, 
    45.32321, 45.31105, 45.29867, 45.28605, 45.27321, 45.26014, 45.24685, 
    45.23332, 45.21957, 45.2056, 45.1914, 45.17697, 45.16232, 45.14744, 
    45.13233, 45.117, 45.10145, 45.08567, 45.06967, 45.05344, 45.03699, 
    45.02032, 45.00342, 44.98631, 44.96896, 44.9514, 44.93361, 44.9156, 
    44.89737, 44.87892, 44.86024, 44.84135, 44.82224, 44.8029, 44.78334, 
    44.76357, 44.74358, 44.72336, 44.70293, 44.68228, 44.66141, 44.64032, 
    44.61902, 44.5975, 44.57576, 44.55381, 44.53164, 44.50925, 44.48665, 
    44.46383, 44.4408, 44.41755, 44.39409, 44.37041, 44.34652, 44.32242, 
    44.29811, 44.27358, 44.24884, 44.22388, 44.19872, 44.17335, 44.14776, 
    44.12197, 44.09596, 44.06975, 44.04332, 44.01669, 43.98985, 43.9628, 
    43.93554, 43.90807, 43.8804, 43.85252, 43.82444, 43.79614, 43.76765, 
    43.73895, 43.71004, 43.68093, 43.65161, 43.62209, 43.59237, 43.56245, 
    43.53232, 43.502, 43.47146, 43.44073, 43.4098, 43.37867, 43.34734, 
    43.31581, 43.28408, 43.25215, 43.22002, 43.18769, 43.15517, 43.12245, 
    43.08954, 43.05643, 43.02312, 42.98962, 42.95592, 42.92203, 42.88794, 
    42.85366, 42.81919, 42.78453, 42.74967, 42.71462, 42.67938, 42.64395, 
    42.60833, 42.57252, 42.53652, 42.50033, 42.46395, 42.42738, 42.39063, 
    42.35369,
  38.26864, 38.32102, 38.37325, 38.42535, 38.47729, 38.52909, 38.58075, 
    38.63226, 38.68362, 38.73484, 38.7859, 38.83682, 38.88759, 38.93821, 
    38.98869, 39.03901, 39.08918, 39.1392, 39.18907, 39.23878, 39.28835, 
    39.33776, 39.38702, 39.43612, 39.48507, 39.53387, 39.58251, 39.63099, 
    39.67932, 39.72749, 39.77551, 39.82336, 39.87106, 39.91861, 39.96599, 
    40.01321, 40.06027, 40.10717, 40.15392, 40.20049, 40.24691, 40.29317, 
    40.33926, 40.38519, 40.43095, 40.47655, 40.52199, 40.56726, 40.61237, 
    40.65731, 40.70208, 40.74669, 40.79113, 40.8354, 40.8795, 40.92344, 
    40.9672, 41.01079, 41.05422, 41.09747, 41.14055, 41.18346, 41.2262, 
    41.26876, 41.31115, 41.35337, 41.39542, 41.43729, 41.47898, 41.5205, 
    41.56184, 41.60301, 41.644, 41.68481, 41.72544, 41.7659, 41.80618, 
    41.84627, 41.88619, 41.92593, 41.96548, 42.00486, 42.04405, 42.08307, 
    42.12189, 42.16054, 42.19901, 42.23729, 42.27538, 42.31329, 42.35101, 
    42.38855, 42.4259, 42.46307, 42.50005, 42.53684, 42.57344, 42.60986, 
    42.64608, 42.68212, 42.71797, 42.75362, 42.78909, 42.82437, 42.85945, 
    42.89434, 42.92904, 42.96354, 42.99786, 43.03197, 43.0659, 43.09963, 
    43.13316, 43.1665, 43.19965, 43.23259, 43.26534, 43.29789, 43.33025, 
    43.36241, 43.39436, 43.42612, 43.45768, 43.48904, 43.5202, 43.55116, 
    43.58192, 43.61248, 43.64283, 43.67299, 43.70293, 43.73268, 43.76223, 
    43.79156, 43.8207, 43.84963, 43.87836, 43.90688, 43.93519, 43.9633, 
    43.9912, 44.01889, 44.04638, 44.07366, 44.10073, 44.12759, 44.15424, 
    44.18069, 44.20692, 44.23295, 44.25876, 44.28436, 44.30975, 44.33493, 
    44.3599, 44.38466, 44.4092, 44.43353, 44.45765, 44.48155, 44.50524, 
    44.52872, 44.55198, 44.57502, 44.59785, 44.62046, 44.64286, 44.66504, 
    44.68701, 44.70876, 44.73029, 44.7516, 44.77269, 44.79357, 44.81423, 
    44.83467, 44.85489, 44.87489, 44.89467, 44.91423, 44.93357, 44.95269, 
    44.97158, 44.99026, 45.00872, 45.02695, 45.04496, 45.06275, 45.08032, 
    45.09766, 45.11478, 45.13168, 45.14835, 45.1648, 45.18102, 45.19703, 
    45.2128, 45.22835, 45.24368, 45.25877, 45.27365, 45.2883, 45.30272, 
    45.31691, 45.33088, 45.34462, 45.35814, 45.37143, 45.38449, 45.39732, 
    45.40993, 45.4223, 45.43445, 45.44637, 45.45806, 45.46952, 45.48076, 
    45.49176, 45.50254, 45.51308, 45.5234, 45.53349, 45.54334, 45.55297, 
    45.56236, 45.57153, 45.58046, 45.58916, 45.59764, 45.60588, 45.61389, 
    45.62167, 45.62922, 45.63654, 45.64362, 45.65047, 45.65709, 45.66348, 
    45.66964, 45.67556, 45.68126, 45.68671, 45.69194, 45.69694, 45.7017, 
    45.70623, 45.71053, 45.71459, 45.71842, 45.72202, 45.72538, 45.72852, 
    45.73141, 45.73408, 45.73651, 45.73871, 45.74068, 45.74241, 45.74391, 
    45.74517, 45.7462, 45.74701, 45.74757, 45.7479, 45.748, 45.74786, 
    45.74749, 45.74689, 45.74606, 45.74499, 45.74369, 45.74215, 45.74038, 
    45.73838, 45.73614, 45.73367, 45.73097, 45.72803, 45.72487, 45.72147, 
    45.71783, 45.71396, 45.70986, 45.70553, 45.70096, 45.69616, 45.69113, 
    45.68587, 45.68037, 45.67464, 45.66868, 45.66249, 45.65606, 45.6494, 
    45.64251, 45.63539, 45.62804, 45.62046, 45.61264, 45.60459, 45.59631, 
    45.58781, 45.57906, 45.5701, 45.56089, 45.55146, 45.5418, 45.53191, 
    45.52178, 45.51143, 45.50085, 45.49004, 45.479, 45.46773, 45.45623, 
    45.4445, 45.43254, 45.42036, 45.40795, 45.39531, 45.38244, 45.36934, 
    45.35602, 45.34246, 45.32869, 45.31468, 45.30045, 45.286, 45.27131, 
    45.2564, 45.24126, 45.22591, 45.21032, 45.19451, 45.17847, 45.16221, 
    45.14573, 45.12902, 45.11209, 45.09493, 45.07755, 45.05995, 45.04213, 
    45.02408, 45.00581, 44.98732, 44.96861, 44.94968, 44.93052, 44.91115, 
    44.89156, 44.87174, 44.8517, 44.83145, 44.81097, 44.79028, 44.76937, 
    44.74824, 44.72689, 44.70533, 44.68355, 44.66155, 44.63933, 44.6169, 
    44.59425, 44.57139, 44.54831, 44.52502, 44.50151, 44.47778, 44.45385, 
    44.4297, 44.40533, 44.38076, 44.35597, 44.33097, 44.30575, 44.28033, 
    44.25469, 44.22884, 44.20279, 44.17652, 44.15004, 44.12336, 44.09646, 
    44.06936, 44.04205, 44.01453, 43.9868, 43.95887, 43.93073, 43.90238, 
    43.87383, 43.84507, 43.8161, 43.78694, 43.75756, 43.72799, 43.69821, 
    43.66823, 43.63805, 43.60766, 43.57707, 43.54628, 43.51529, 43.4841, 
    43.45271, 43.42111, 43.38932, 43.35733, 43.32515, 43.29276, 43.26017, 
    43.22739, 43.19442, 43.16124, 43.12787, 43.09431, 43.06055, 43.02659, 
    42.99244, 42.9581, 42.92356, 42.88883, 42.85391, 42.8188, 42.78349, 
    42.748, 42.71231, 42.67643, 42.64037, 42.60411, 42.56767, 42.53103, 
    42.49421, 42.4572,
  38.3652, 38.41766, 38.46997, 38.52214, 38.57417, 38.62605, 38.67778, 
    38.72937, 38.78081, 38.8321, 38.88325, 38.93425, 38.9851, 39.03579, 
    39.08634, 39.13675, 39.18699, 39.23709, 39.28704, 39.33683, 39.38647, 
    39.43596, 39.4853, 39.53448, 39.58351, 39.63238, 39.6811, 39.72966, 
    39.77807, 39.82632, 39.87441, 39.92234, 39.97012, 40.01773, 40.06519, 
    40.11249, 40.15963, 40.20661, 40.25343, 40.30008, 40.34658, 40.39291, 
    40.43908, 40.48508, 40.53092, 40.5766, 40.62211, 40.66746, 40.71264, 
    40.75766, 40.80251, 40.84719, 40.8917, 40.93605, 40.98022, 41.02423, 
    41.06807, 41.11174, 41.15524, 41.19856, 41.24171, 41.2847, 41.32751, 
    41.37015, 41.41261, 41.4549, 41.49702, 41.53896, 41.58073, 41.62232, 
    41.66373, 41.70497, 41.74603, 41.78692, 41.82762, 41.86815, 41.9085, 
    41.94867, 41.98866, 42.02846, 42.06809, 42.10754, 42.1468, 42.18588, 
    42.22478, 42.2635, 42.30203, 42.34038, 42.37854, 42.41652, 42.45431, 
    42.49192, 42.52934, 42.56657, 42.60362, 42.64048, 42.67715, 42.71363, 
    42.74992, 42.78603, 42.82194, 42.85766, 42.89319, 42.92853, 42.96368, 
    42.99864, 43.0334, 43.06797, 43.10235, 43.13653, 43.17052, 43.20431, 
    43.23791, 43.27131, 43.30452, 43.33752, 43.37034, 43.40295, 43.43537, 
    43.46759, 43.4996, 43.53143, 43.56305, 43.59446, 43.62568, 43.6567, 
    43.68752, 43.71814, 43.74855, 43.77876, 43.80877, 43.83857, 43.86818, 
    43.89757, 43.92676, 43.95575, 43.98453, 44.01311, 44.04148, 44.06964, 
    44.0976, 44.12534, 44.15289, 44.18022, 44.20734, 44.23426, 44.26096, 
    44.28746, 44.31374, 44.33982, 44.36568, 44.39134, 44.41678, 44.44201, 
    44.46703, 44.49183, 44.51643, 44.54081, 44.56497, 44.58892, 44.61266, 
    44.63618, 44.65949, 44.68258, 44.70546, 44.72812, 44.75056, 44.77279, 
    44.7948, 44.81659, 44.83816, 44.85952, 44.88065, 44.90157, 44.92228, 
    44.94275, 44.96302, 44.98306, 45.00288, 45.02248, 45.04186, 45.06102, 
    45.07995, 45.09867, 45.11716, 45.13543, 45.15348, 45.17131, 45.18891, 
    45.20629, 45.22345, 45.24038, 45.25708, 45.27357, 45.28983, 45.30586, 
    45.32167, 45.33725, 45.35261, 45.36774, 45.38264, 45.39732, 45.41177, 
    45.426, 45.44, 45.45377, 45.46731, 45.48063, 45.49372, 45.50658, 
    45.51921, 45.53161, 45.54379, 45.55573, 45.56745, 45.57893, 45.59019, 
    45.60122, 45.61201, 45.62259, 45.63292, 45.64303, 45.6529, 45.66255, 
    45.67197, 45.68115, 45.69011, 45.69883, 45.70732, 45.71558, 45.72361, 
    45.7314, 45.73896, 45.7463, 45.7534, 45.76027, 45.7669, 45.7733, 
    45.77947, 45.78541, 45.79111, 45.79659, 45.80182, 45.80683, 45.8116, 
    45.81614, 45.82045, 45.82452, 45.82836, 45.83196, 45.83533, 45.83847, 
    45.84138, 45.84405, 45.84649, 45.84869, 45.85066, 45.8524, 45.8539, 
    45.85517, 45.8562, 45.857, 45.85757, 45.8579, 45.858, 45.85786, 45.85749, 
    45.85689, 45.85605, 45.85498, 45.85368, 45.85214, 45.85036, 45.84836, 
    45.84612, 45.84364, 45.84093, 45.83799, 45.83482, 45.83141, 45.82777, 
    45.82389, 45.81978, 45.81544, 45.81086, 45.80605, 45.80101, 45.79573, 
    45.79023, 45.78448, 45.77851, 45.7723, 45.76587, 45.75919, 45.75229, 
    45.74515, 45.73779, 45.73018, 45.72235, 45.71429, 45.70599, 45.69746, 
    45.68871, 45.67971, 45.67049, 45.66104, 45.65136, 45.64145, 45.6313, 
    45.62093, 45.61032, 45.59949, 45.58842, 45.57713, 45.56561, 45.55386, 
    45.54187, 45.52966, 45.51722, 45.50456, 45.49166, 45.47854, 45.46519, 
    45.45161, 45.4378, 45.42376, 45.4095, 45.39502, 45.3803, 45.36536, 
    45.35019, 45.3348, 45.31918, 45.30334, 45.28727, 45.27097, 45.25446, 
    45.23771, 45.22075, 45.20356, 45.18614, 45.1685, 45.15064, 45.13256, 
    45.11425, 45.09572, 45.07697, 45.058, 45.03881, 45.01939, 44.99976, 
    44.9799, 44.95983, 44.93953, 44.91901, 44.89828, 44.87733, 44.85615, 
    44.83476, 44.81315, 44.79133, 44.76928, 44.74702, 44.72454, 44.70185, 
    44.67894, 44.65582, 44.63247, 44.60892, 44.58515, 44.56116, 44.53696, 
    44.51255, 44.48792, 44.46309, 44.43803, 44.41277, 44.38729, 44.36161, 
    44.33571, 44.3096, 44.28328, 44.25675, 44.23001, 44.20306, 44.17591, 
    44.14854, 44.12097, 44.09319, 44.0652, 44.037, 44.0086, 43.97999, 
    43.95118, 43.92216, 43.89293, 43.86351, 43.83387, 43.80404, 43.77399, 
    43.74375, 43.71331, 43.68266, 43.65181, 43.62076, 43.58951, 43.55806, 
    43.52641, 43.49455, 43.4625, 43.43025, 43.3978, 43.36516, 43.33232, 
    43.29928, 43.26604, 43.23261, 43.19898, 43.16515, 43.13113, 43.09692, 
    43.06252, 43.02792, 42.99312, 42.95813, 42.92295, 42.88758, 42.85202, 
    42.81627, 42.78033, 42.74419, 42.70787, 42.67136, 42.63466, 42.59777, 
    42.5607,
  38.46172, 38.51426, 38.56665, 38.6189, 38.67101, 38.72296, 38.77478, 
    38.82644, 38.87796, 38.92933, 38.98056, 39.03163, 39.08256, 39.13334, 
    39.18397, 39.23444, 39.28477, 39.33495, 39.38497, 39.43484, 39.48457, 
    39.53413, 39.58355, 39.6328, 39.68191, 39.73086, 39.77966, 39.8283, 
    39.87678, 39.92511, 39.97327, 40.02129, 40.06914, 40.11683, 40.16437, 
    40.21175, 40.25896, 40.30602, 40.35291, 40.39964, 40.44621, 40.49262, 
    40.53886, 40.58495, 40.63086, 40.67661, 40.7222, 40.76762, 40.81288, 
    40.85797, 40.9029, 40.94765, 40.99224, 41.03666, 41.08091, 41.125, 
    41.16891, 41.21265, 41.25622, 41.29962, 41.34285, 41.38591, 41.42879, 
    41.4715, 41.51404, 41.55641, 41.5986, 41.64061, 41.68245, 41.72411, 
    41.7656, 41.80691, 41.84805, 41.889, 41.92978, 41.97038, 42.0108, 
    42.05103, 42.09109, 42.13097, 42.17067, 42.21019, 42.24952, 42.28867, 
    42.32764, 42.36643, 42.40503, 42.44345, 42.48168, 42.51973, 42.55759, 
    42.59526, 42.63275, 42.67006, 42.70717, 42.74409, 42.78083, 42.81738, 
    42.85374, 42.88991, 42.92589, 42.96168, 42.99728, 43.03268, 43.06789, 
    43.10292, 43.13774, 43.17238, 43.20682, 43.24107, 43.27512, 43.30898, 
    43.34264, 43.3761, 43.40937, 43.44244, 43.47532, 43.50799, 43.54047, 
    43.57275, 43.60483, 43.63671, 43.66839, 43.69987, 43.73115, 43.76223, 
    43.79311, 43.82378, 43.85425, 43.88452, 43.91459, 43.94445, 43.97411, 
    44.00356, 44.03281, 44.06186, 44.09069, 44.11932, 44.14775, 44.17596, 
    44.20398, 44.23178, 44.25938, 44.28676, 44.31394, 44.34091, 44.36767, 
    44.39421, 44.42056, 44.44668, 44.4726, 44.4983, 44.5238, 44.54908, 
    44.57414, 44.599, 44.62364, 44.64807, 44.67228, 44.69628, 44.72007, 
    44.74364, 44.76699, 44.79013, 44.81305, 44.83576, 44.85825, 44.88052, 
    44.90257, 44.92441, 44.94603, 44.96743, 44.98861, 45.00957, 45.03031, 
    45.05083, 45.07114, 45.09122, 45.11108, 45.13072, 45.15014, 45.16934, 
    45.18832, 45.20707, 45.2256, 45.24391, 45.262, 45.27986, 45.2975, 
    45.31491, 45.3321, 45.34907, 45.36581, 45.38233, 45.39862, 45.41469, 
    45.43053, 45.44615, 45.46154, 45.4767, 45.49163, 45.50634, 45.52083, 
    45.53508, 45.54911, 45.56291, 45.57648, 45.58982, 45.60294, 45.61583, 
    45.62849, 45.64091, 45.65311, 45.66508, 45.67683, 45.68834, 45.69962, 
    45.71067, 45.72149, 45.73208, 45.74244, 45.75257, 45.76247, 45.77213, 
    45.78157, 45.79078, 45.79975, 45.80849, 45.817, 45.82527, 45.83332, 
    45.84113, 45.84871, 45.85606, 45.86317, 45.87005, 45.87671, 45.88312, 
    45.8893, 45.89525, 45.90097, 45.90645, 45.9117, 45.91672, 45.9215, 
    45.92605, 45.93037, 45.93445, 45.93829, 45.94191, 45.94529, 45.94843, 
    45.95134, 45.95402, 45.95646, 45.95867, 45.96064, 45.96238, 45.96389, 
    45.96516, 45.9662, 45.967, 45.96757, 45.9679, 45.968, 45.96786, 45.96749, 
    45.96689, 45.96605, 45.96498, 45.96367, 45.96212, 45.96035, 45.95834, 
    45.95609, 45.95361, 45.9509, 45.94795, 45.94477, 45.94135, 45.9377, 
    45.93382, 45.9297, 45.92535, 45.92076, 45.91594, 45.91089, 45.9056, 
    45.90008, 45.89433, 45.88834, 45.88212, 45.87567, 45.86898, 45.86206, 
    45.85491, 45.84753, 45.83991, 45.83206, 45.82398, 45.81567, 45.80712, 
    45.79834, 45.78933, 45.78009, 45.77062, 45.76092, 45.75098, 45.74082, 
    45.73042, 45.7198, 45.70894, 45.69785, 45.68653, 45.67498, 45.66321, 
    45.6512, 45.63897, 45.6265, 45.6138, 45.60088, 45.58773, 45.57435, 
    45.56074, 45.54691, 45.53284, 45.51855, 45.50403, 45.48929, 45.47432, 
    45.45912, 45.44369, 45.42804, 45.41216, 45.39606, 45.37973, 45.36318, 
    45.3464, 45.3294, 45.31217, 45.29472, 45.27705, 45.25915, 45.24103, 
    45.22268, 45.20412, 45.18533, 45.16632, 45.14708, 45.12763, 45.10795, 
    45.08806, 45.06794, 45.0476, 45.02705, 45.00627, 44.98527, 44.96405, 
    44.94262, 44.92097, 44.8991, 44.87701, 44.8547, 44.83218, 44.80944, 
    44.78648, 44.76331, 44.73992, 44.71632, 44.6925, 44.66846, 44.64422, 
    44.61976, 44.59508, 44.57019, 44.54509, 44.51978, 44.49425, 44.46851, 
    44.44256, 44.4164, 44.39003, 44.36345, 44.33665, 44.30965, 44.28244, 
    44.25502, 44.2274, 44.19956, 44.17152, 44.14326, 44.11481, 44.08614, 
    44.05727, 44.0282, 43.99892, 43.96943, 43.93974, 43.90984, 43.87975, 
    43.84945, 43.81894, 43.78823, 43.75732, 43.72622, 43.6949, 43.66339, 
    43.63168, 43.59977, 43.56765, 43.53534, 43.50283, 43.47013, 43.43722, 
    43.40412, 43.37082, 43.33732, 43.30363, 43.26974, 43.23566, 43.20139, 
    43.16691, 43.13225, 43.09739, 43.06234, 43.02709, 42.99166, 42.95603, 
    42.92021, 42.8842, 42.848, 42.81161, 42.77503, 42.73827, 42.70131, 
    42.66417,
  38.5582, 38.61082, 38.66329, 38.71562, 38.7678, 38.81984, 38.87173, 
    38.92348, 38.97507, 39.02652, 39.07783, 39.12898, 39.17999, 39.23084, 
    39.28155, 39.33211, 39.38251, 39.43277, 39.48287, 39.53282, 39.58262, 
    39.63227, 39.68176, 39.73109, 39.78028, 39.82931, 39.87818, 39.9269, 
    39.97546, 40.02386, 40.07211, 40.1202, 40.16813, 40.2159, 40.26351, 
    40.31096, 40.35825, 40.40539, 40.45236, 40.49916, 40.54581, 40.5923, 
    40.63862, 40.68478, 40.73077, 40.7766, 40.82226, 40.86776, 40.91309, 
    40.95826, 41.00326, 41.04809, 41.09275, 41.13725, 41.18157, 41.22573, 
    41.26972, 41.31353, 41.35718, 41.40066, 41.44396, 41.48709, 41.53005, 
    41.57283, 41.61544, 41.65788, 41.70015, 41.74223, 41.78415, 41.82588, 
    41.86744, 41.90882, 41.95003, 41.99106, 42.03191, 42.07257, 42.11307, 
    42.15338, 42.19351, 42.23346, 42.27323, 42.31281, 42.35222, 42.39144, 
    42.43048, 42.46933, 42.50801, 42.54649, 42.58479, 42.62291, 42.66084, 
    42.69859, 42.73614, 42.77351, 42.8107, 42.84769, 42.88449, 42.92111, 
    42.95753, 42.99377, 43.02982, 43.06567, 43.10133, 43.13681, 43.17208, 
    43.20717, 43.24207, 43.27676, 43.31127, 43.34558, 43.3797, 43.41362, 
    43.44734, 43.48087, 43.5142, 43.54734, 43.58027, 43.61301, 43.64555, 
    43.67789, 43.71003, 43.74197, 43.77372, 43.80526, 43.8366, 43.86774, 
    43.89867, 43.92941, 43.95994, 43.99026, 44.02039, 44.05031, 44.08002, 
    44.10954, 44.13884, 44.16794, 44.19684, 44.22552, 44.25401, 44.28228, 
    44.31034, 44.3382, 44.36585, 44.3933, 44.42052, 44.44755, 44.47436, 
    44.50096, 44.52735, 44.55353, 44.5795, 44.60526, 44.6308, 44.65613, 
    44.68125, 44.70615, 44.73085, 44.75532, 44.77958, 44.80363, 44.82747, 
    44.85108, 44.87449, 44.89767, 44.92064, 44.94339, 44.96592, 44.98824, 
    45.01034, 45.03222, 45.05388, 45.07533, 45.09655, 45.11756, 45.13834, 
    45.15891, 45.17925, 45.19938, 45.21928, 45.23896, 45.25842, 45.27766, 
    45.29667, 45.31546, 45.33403, 45.35238, 45.3705, 45.3884, 45.40608, 
    45.42353, 45.44076, 45.45776, 45.47454, 45.49109, 45.50742, 45.52352, 
    45.53939, 45.55504, 45.57046, 45.58566, 45.60062, 45.61536, 45.62988, 
    45.64416, 45.65822, 45.67205, 45.68565, 45.69902, 45.71216, 45.72508, 
    45.73776, 45.75022, 45.76244, 45.77444, 45.78621, 45.79774, 45.80904, 
    45.82012, 45.83096, 45.84158, 45.85196, 45.86211, 45.87203, 45.88171, 
    45.89117, 45.90039, 45.90939, 45.91814, 45.92667, 45.93497, 45.94303, 
    45.95086, 45.95845, 45.96582, 45.97295, 45.97984, 45.98651, 45.99294, 
    45.99913, 46.0051, 46.01083, 46.01632, 46.02158, 46.02661, 46.0314, 
    46.03596, 46.04028, 46.04438, 46.04823, 46.05185, 46.05524, 46.05839, 
    46.06131, 46.06399, 46.06644, 46.06865, 46.07063, 46.07237, 46.07388, 
    46.07515, 46.07619, 46.077, 46.07757, 46.0779, 46.078, 46.07786, 
    46.07749, 46.07689, 46.07605, 46.07497, 46.07366, 46.07211, 46.07033, 
    46.06832, 46.06607, 46.06358, 46.06086, 46.05791, 46.05472, 46.05129, 
    46.04763, 46.04374, 46.03962, 46.03526, 46.03066, 46.02583, 46.02076, 
    46.01547, 46.00993, 46.00417, 45.99817, 45.99194, 45.98547, 45.97877, 
    45.97184, 45.96467, 45.95727, 45.94963, 45.94177, 45.93367, 45.92534, 
    45.91677, 45.90798, 45.89895, 45.88969, 45.8802, 45.87048, 45.86052, 
    45.85033, 45.83991, 45.82927, 45.81838, 45.80727, 45.79593, 45.78436, 
    45.77256, 45.76052, 45.74826, 45.73577, 45.72305, 45.7101, 45.69692, 
    45.68351, 45.66988, 45.65601, 45.64192, 45.62759, 45.61305, 45.59827, 
    45.58327, 45.56804, 45.55258, 45.5369, 45.52098, 45.50485, 45.48849, 
    45.4719, 45.45509, 45.43805, 45.42078, 45.4033, 45.38559, 45.36765, 
    45.34949, 45.33111, 45.31251, 45.29368, 45.27463, 45.25536, 45.23586, 
    45.21614, 45.19621, 45.17605, 45.15567, 45.13507, 45.11425, 45.09321, 
    45.07195, 45.05047, 45.02877, 45.00686, 44.98473, 44.96238, 44.9398, 
    44.91702, 44.89402, 44.8708, 44.84736, 44.82371, 44.79984, 44.77576, 
    44.75146, 44.72695, 44.70223, 44.67729, 44.65214, 44.62677, 44.6012, 
    44.57541, 44.5494, 44.52319, 44.49677, 44.47013, 44.44329, 44.41623, 
    44.38897, 44.36149, 44.33381, 44.30592, 44.27782, 44.24952, 44.221, 
    44.19228, 44.16335, 44.13422, 44.10488, 44.07534, 44.04559, 44.01564, 
    43.98548, 43.95512, 43.92456, 43.89379, 43.86282, 43.83165, 43.80028, 
    43.76871, 43.73693, 43.70496, 43.67279, 43.64042, 43.60785, 43.57508, 
    43.54211, 43.50894, 43.47558, 43.44202, 43.40826, 43.37431, 43.34017, 
    43.30582, 43.27129, 43.23656, 43.20164, 43.16652, 43.13121, 43.09571, 
    43.06001, 43.02413, 42.98805, 42.95179, 42.91533, 42.87868, 42.84185, 
    42.80482, 42.76761,
  38.65465, 38.70734, 38.7599, 38.8123, 38.86456, 38.91668, 38.96865, 
    39.02047, 39.07215, 39.12368, 39.17506, 39.2263, 39.27738, 39.32832, 
    39.3791, 39.42973, 39.48022, 39.53055, 39.58073, 39.63076, 39.68064, 
    39.73036, 39.77993, 39.82935, 39.87861, 39.92772, 39.97667, 40.02546, 
    40.0741, 40.12258, 40.17091, 40.21907, 40.26708, 40.31493, 40.36262, 
    40.41014, 40.45752, 40.50473, 40.55177, 40.59866, 40.64538, 40.69194, 
    40.73834, 40.78457, 40.83064, 40.87655, 40.92229, 40.96786, 41.01327, 
    41.05851, 41.10358, 41.14849, 41.19323, 41.2378, 41.2822, 41.32644, 
    41.3705, 41.41439, 41.45811, 41.50166, 41.54504, 41.58824, 41.63128, 
    41.67413, 41.71682, 41.75933, 41.80167, 41.84383, 41.88581, 41.92762, 
    41.96925, 42.01071, 42.05199, 42.09309, 42.13401, 42.17475, 42.21531, 
    42.2557, 42.2959, 42.33592, 42.37576, 42.41542, 42.45489, 42.49418, 
    42.53329, 42.57222, 42.61096, 42.64951, 42.68789, 42.72607, 42.76407, 
    42.80188, 42.83951, 42.87695, 42.9142, 42.95126, 42.98813, 43.02481, 
    43.06131, 43.09761, 43.13372, 43.16965, 43.20538, 43.24091, 43.27626, 
    43.31141, 43.34637, 43.38113, 43.4157, 43.45008, 43.48426, 43.51824, 
    43.55203, 43.58562, 43.61902, 43.65221, 43.68521, 43.71801, 43.75062, 
    43.78302, 43.81522, 43.84723, 43.87903, 43.91063, 43.94203, 43.97323, 
    44.00422, 44.03502, 44.06561, 44.09599, 44.12618, 44.15615, 44.18593, 
    44.2155, 44.24486, 44.27402, 44.30297, 44.33171, 44.36025, 44.38858, 
    44.4167, 44.44461, 44.47232, 44.49981, 44.5271, 44.55417, 44.58104, 
    44.60769, 44.63414, 44.66037, 44.68639, 44.7122, 44.73779, 44.76317, 
    44.78834, 44.8133, 44.83804, 44.86256, 44.88688, 44.91097, 44.93485, 
    44.95852, 44.98197, 45.0052, 45.02821, 45.05101, 45.07359, 45.09595, 
    45.1181, 45.14003, 45.16173, 45.18322, 45.20449, 45.22554, 45.24636, 
    45.26697, 45.28736, 45.30752, 45.32747, 45.34719, 45.36669, 45.38597, 
    45.40502, 45.42385, 45.44246, 45.46085, 45.47901, 45.49694, 45.51466, 
    45.53214, 45.54941, 45.56644, 45.58326, 45.59984, 45.6162, 45.63234, 
    45.64825, 45.66393, 45.67938, 45.69461, 45.70961, 45.72438, 45.73892, 
    45.75324, 45.76732, 45.78118, 45.79481, 45.80821, 45.82138, 45.83432, 
    45.84703, 45.85952, 45.87177, 45.88379, 45.89558, 45.90714, 45.91847, 
    45.92957, 45.94043, 45.95107, 45.96148, 45.97165, 45.98159, 45.99129, 
    46.00077, 46.01001, 46.01902, 46.0278, 46.03635, 46.04466, 46.05274, 
    46.06059, 46.0682, 46.07558, 46.08272, 46.08963, 46.09631, 46.10275, 
    46.10896, 46.11494, 46.12068, 46.12619, 46.13146, 46.1365, 46.1413, 
    46.14587, 46.1502, 46.1543, 46.15816, 46.1618, 46.16519, 46.16835, 
    46.17127, 46.17396, 46.17641, 46.17863, 46.18061, 46.18236, 46.18387, 
    46.18515, 46.18619, 46.187, 46.18756, 46.1879, 46.188, 46.18786, 
    46.18749, 46.18688, 46.18604, 46.18496, 46.18365, 46.1821, 46.18032, 
    46.1783, 46.17604, 46.17355, 46.17083, 46.16786, 46.16467, 46.16124, 
    46.15757, 46.15367, 46.14953, 46.14516, 46.14056, 46.13572, 46.13064, 
    46.12533, 46.11979, 46.11401, 46.108, 46.10175, 46.09527, 46.08855, 
    46.08161, 46.07442, 46.06701, 46.05936, 46.05148, 46.04336, 46.03501, 
    46.02643, 46.01762, 46.00857, 45.99929, 45.98977, 45.98003, 45.97005, 
    45.95984, 45.9494, 45.93873, 45.92783, 45.91669, 45.90533, 45.89373, 
    45.8819, 45.86985, 45.85756, 45.84504, 45.83229, 45.81931, 45.80611, 
    45.79267, 45.779, 45.76511, 45.75099, 45.73664, 45.72206, 45.70725, 
    45.69221, 45.67695, 45.66146, 45.64574, 45.6298, 45.61363, 45.59724, 
    45.58061, 45.56377, 45.54669, 45.52939, 45.51187, 45.49412, 45.47615, 
    45.45795, 45.43953, 45.42089, 45.40202, 45.38293, 45.36362, 45.34408, 
    45.32433, 45.30435, 45.28415, 45.26373, 45.24308, 45.22222, 45.20114, 
    45.17984, 45.15831, 45.13657, 45.11461, 45.09243, 45.07004, 45.04742, 
    45.02459, 45.00154, 44.97827, 44.95479, 44.93109, 44.90718, 44.88305, 
    44.8587, 44.83414, 44.80936, 44.78437, 44.75917, 44.73376, 44.70813, 
    44.68229, 44.65623, 44.62997, 44.60349, 44.57681, 44.5499, 44.5228, 
    44.49548, 44.46795, 44.44021, 44.41227, 44.38411, 44.35575, 44.32718, 
    44.2984, 44.26942, 44.24023, 44.21083, 44.18123, 44.15143, 44.12142, 
    44.0912, 44.06078, 44.03016, 43.99933, 43.96831, 43.93708, 43.90564, 
    43.87401, 43.84217, 43.81014, 43.77791, 43.74547, 43.71284, 43.68001, 
    43.64698, 43.61375, 43.58032, 43.5467, 43.51288, 43.47887, 43.44465, 
    43.41025, 43.37565, 43.34085, 43.30586, 43.27068, 43.23531, 43.19974, 
    43.16397, 43.12803, 43.09188, 43.05555, 43.01902, 42.98231, 42.94541, 
    42.90832, 42.87104,
  38.75106, 38.80383, 38.85646, 38.90895, 38.96129, 39.01348, 39.06553, 
    39.11744, 39.16919, 39.2208, 39.27226, 39.32357, 39.37473, 39.42575, 
    39.47661, 39.52732, 39.57789, 39.6283, 39.67856, 39.72867, 39.77862, 
    39.82842, 39.87807, 39.92757, 39.97691, 40.02609, 40.07512, 40.12399, 
    40.17271, 40.22127, 40.26967, 40.31791, 40.366, 40.41392, 40.46169, 
    40.5093, 40.55674, 40.60403, 40.65115, 40.69812, 40.74492, 40.79155, 
    40.83803, 40.88434, 40.93048, 40.97647, 41.02228, 41.06793, 41.11342, 
    41.15873, 41.20388, 41.24887, 41.29368, 41.33833, 41.3828, 41.42711, 
    41.47125, 41.51522, 41.55901, 41.60263, 41.64609, 41.68937, 41.73247, 
    41.77541, 41.81816, 41.86075, 41.90316, 41.9454, 41.98745, 42.02934, 
    42.07104, 42.11257, 42.15392, 42.19509, 42.23608, 42.2769, 42.31753, 
    42.35799, 42.39826, 42.43835, 42.47826, 42.51799, 42.55754, 42.5969, 
    42.63608, 42.67508, 42.71389, 42.75251, 42.79095, 42.82921, 42.86728, 
    42.90516, 42.94285, 42.98036, 43.01768, 43.05481, 43.09175, 43.1285, 
    43.16506, 43.20143, 43.23761, 43.2736, 43.30939, 43.345, 43.38041, 
    43.41563, 43.45065, 43.48548, 43.52011, 43.55455, 43.5888, 43.62285, 
    43.6567, 43.69036, 43.72382, 43.75708, 43.79014, 43.823, 43.85566, 
    43.88813, 43.92039, 43.95246, 43.98432, 44.01598, 44.04744, 44.0787, 
    44.10976, 44.14061, 44.17126, 44.20171, 44.23195, 44.26199, 44.29182, 
    44.32145, 44.35086, 44.38008, 44.40909, 44.43789, 44.46648, 44.49487, 
    44.52304, 44.55101, 44.57877, 44.60632, 44.63366, 44.66079, 44.68771, 
    44.71441, 44.74091, 44.7672, 44.79327, 44.81913, 44.84477, 44.8702, 
    44.89542, 44.92043, 44.94522, 44.9698, 44.99416, 45.0183, 45.04223, 
    45.06594, 45.08944, 45.11272, 45.13578, 45.15863, 45.18126, 45.20366, 
    45.22585, 45.24782, 45.26957, 45.29111, 45.31242, 45.33351, 45.35438, 
    45.37503, 45.39546, 45.41566, 45.43565, 45.45541, 45.47495, 45.49427, 
    45.51336, 45.53223, 45.55088, 45.56931, 45.5875, 45.60548, 45.62323, 
    45.64075, 45.65805, 45.67513, 45.69197, 45.70859, 45.72499, 45.74115, 
    45.7571, 45.77281, 45.7883, 45.80355, 45.81859, 45.83339, 45.84796, 
    45.86231, 45.87643, 45.89031, 45.90397, 45.9174, 45.9306, 45.94357, 
    45.95631, 45.96881, 45.98109, 45.99314, 46.00496, 46.01654, 46.02789, 
    46.03901, 46.0499, 46.06056, 46.07099, 46.08118, 46.09114, 46.10087, 
    46.11037, 46.11963, 46.12866, 46.13746, 46.14602, 46.15435, 46.16245, 
    46.17031, 46.17794, 46.18533, 46.19249, 46.19942, 46.20611, 46.21257, 
    46.2188, 46.22478, 46.23054, 46.23605, 46.24134, 46.24639, 46.2512, 
    46.25578, 46.26012, 46.26423, 46.2681, 46.27174, 46.27514, 46.27831, 
    46.28123, 46.28393, 46.28639, 46.28861, 46.2906, 46.29235, 46.29387, 
    46.29514, 46.29618, 46.29699, 46.29757, 46.2979, 46.298, 46.29786, 
    46.29749, 46.29688, 46.29604, 46.29496, 46.29364, 46.29209, 46.2903, 
    46.28828, 46.28601, 46.28352, 46.28079, 46.27782, 46.27462, 46.27118, 
    46.26751, 46.2636, 46.25945, 46.25507, 46.25045, 46.24561, 46.24052, 
    46.2352, 46.22964, 46.22385, 46.21783, 46.21157, 46.20507, 46.19834, 
    46.19138, 46.18418, 46.17675, 46.16908, 46.16118, 46.15305, 46.14468, 
    46.13608, 46.12725, 46.11818, 46.10888, 46.09935, 46.08958, 46.07959, 
    46.06936, 46.05889, 46.0482, 46.03727, 46.02611, 46.01472, 46.0031, 
    45.99125, 45.97916, 45.96685, 45.95431, 45.94153, 45.92852, 45.91529, 
    45.90182, 45.88813, 45.87421, 45.86005, 45.84567, 45.83106, 45.81622, 
    45.80116, 45.78586, 45.77034, 45.75459, 45.73861, 45.72241, 45.70598, 
    45.68932, 45.67244, 45.65533, 45.63799, 45.62043, 45.60265, 45.58464, 
    45.56641, 45.54795, 45.52926, 45.51036, 45.49123, 45.47187, 45.4523, 
    45.4325, 45.41248, 45.39224, 45.37178, 45.35109, 45.33019, 45.30906, 
    45.28772, 45.26615, 45.24436, 45.22236, 45.20013, 45.17769, 45.15503, 
    45.13215, 45.10905, 45.08574, 45.06221, 45.03846, 45.0145, 44.99032, 
    44.96592, 44.94131, 44.91649, 44.89145, 44.8662, 44.84073, 44.81505, 
    44.78916, 44.76305, 44.73673, 44.71021, 44.68346, 44.65651, 44.62935, 
    44.60197, 44.57439, 44.5466, 44.5186, 44.49039, 44.46197, 44.43335, 
    44.40451, 44.37547, 44.34623, 44.31677, 44.28711, 44.25725, 44.22718, 
    44.19691, 44.16643, 44.13575, 44.10486, 44.07377, 44.04248, 44.01099, 
    43.97929, 43.9474, 43.9153, 43.88301, 43.85051, 43.81781, 43.78492, 
    43.75183, 43.71854, 43.68505, 43.65136, 43.61748, 43.5834, 43.54912, 
    43.51465, 43.47998, 43.44513, 43.41007, 43.37482, 43.33938, 43.30375, 
    43.26792, 43.2319, 43.19569, 43.15929, 43.1227, 43.08592, 43.04895, 
    43.01179, 42.97444,
  38.84742, 38.90028, 38.95298, 39.00555, 39.05797, 39.11024, 39.16237, 
    39.21436, 39.26619, 39.31788, 39.36942, 39.42081, 39.47205, 39.52314, 
    39.57409, 39.62488, 39.67552, 39.72601, 39.77635, 39.82653, 39.87657, 
    39.92645, 39.97617, 40.02575, 40.07516, 40.12443, 40.17353, 40.22248, 
    40.27128, 40.31992, 40.3684, 40.41672, 40.46488, 40.51289, 40.56073, 
    40.60841, 40.65594, 40.7033, 40.7505, 40.79754, 40.84442, 40.89113, 
    40.93768, 40.98407, 41.0303, 41.07635, 41.12225, 41.16797, 41.21353, 
    41.25893, 41.30415, 41.34921, 41.3941, 41.43882, 41.48338, 41.52776, 
    41.57197, 41.61601, 41.65988, 41.70358, 41.74711, 41.79046, 41.83364, 
    41.87665, 41.91948, 41.96214, 42.00462, 42.04693, 42.08907, 42.13102, 
    42.1728, 42.2144, 42.25582, 42.29707, 42.33813, 42.37902, 42.41973, 
    42.46025, 42.5006, 42.54076, 42.58074, 42.62054, 42.66016, 42.69959, 
    42.73884, 42.77791, 42.81679, 42.85549, 42.894, 42.93232, 42.97046, 
    43.00841, 43.04617, 43.08375, 43.12114, 43.15833, 43.19534, 43.23216, 
    43.26879, 43.30523, 43.34148, 43.37753, 43.41339, 43.44906, 43.48454, 
    43.51982, 43.55491, 43.58981, 43.62451, 43.65901, 43.69332, 43.72744, 
    43.76135, 43.79507, 43.82859, 43.86192, 43.89504, 43.92797, 43.96069, 
    43.99322, 44.02555, 44.05767, 44.0896, 44.12132, 44.15284, 44.18416, 
    44.21528, 44.24619, 44.2769, 44.30741, 44.33771, 44.3678, 44.39769, 
    44.42738, 44.45686, 44.48613, 44.51519, 44.54405, 44.5727, 44.60114, 
    44.62937, 44.65739, 44.68521, 44.71281, 44.74021, 44.76739, 44.79436, 
    44.82113, 44.84767, 44.87401, 44.90014, 44.92604, 44.95174, 44.97723, 
    45.00249, 45.02755, 45.05239, 45.07702, 45.10143, 45.12562, 45.1496, 
    45.17336, 45.19691, 45.22023, 45.24334, 45.26624, 45.28891, 45.31136, 
    45.3336, 45.35561, 45.37741, 45.39898, 45.42034, 45.44147, 45.46239, 
    45.48308, 45.50355, 45.5238, 45.54382, 45.56363, 45.58321, 45.60257, 
    45.6217, 45.64061, 45.65929, 45.67776, 45.696, 45.714, 45.73179, 
    45.74936, 45.76669, 45.7838, 45.80068, 45.81734, 45.83377, 45.84997, 
    45.86594, 45.88169, 45.89721, 45.9125, 45.92756, 45.94239, 45.957, 
    45.97138, 45.98552, 45.99944, 46.01313, 46.02658, 46.03981, 46.05281, 
    46.06557, 46.07811, 46.09041, 46.10249, 46.11433, 46.12593, 46.13731, 
    46.14846, 46.15937, 46.17005, 46.1805, 46.19072, 46.2007, 46.21045, 
    46.21996, 46.22925, 46.2383, 46.24711, 46.2557, 46.26404, 46.27216, 
    46.28004, 46.28768, 46.29509, 46.30227, 46.30921, 46.31591, 46.32239, 
    46.32862, 46.33463, 46.34039, 46.34592, 46.35122, 46.35627, 46.3611, 
    46.36569, 46.37004, 46.37416, 46.37804, 46.38168, 46.38509, 46.38826, 
    46.3912, 46.3939, 46.39636, 46.39859, 46.40058, 46.40234, 46.40385, 
    46.40514, 46.40618, 46.40699, 46.40756, 46.4079, 46.408, 46.40786, 
    46.40749, 46.40688, 46.40603, 46.40495, 46.40363, 46.40207, 46.40028, 
    46.39825, 46.39599, 46.39349, 46.39075, 46.38778, 46.38457, 46.38112, 
    46.37744, 46.37352, 46.36937, 46.36498, 46.36035, 46.35549, 46.3504, 
    46.34506, 46.33949, 46.33369, 46.32765, 46.32138, 46.31487, 46.30812, 
    46.30115, 46.29393, 46.28649, 46.2788, 46.27089, 46.26274, 46.25435, 
    46.24573, 46.23688, 46.22779, 46.21848, 46.20892, 46.19913, 46.18911, 
    46.17886, 46.16838, 46.15766, 46.14671, 46.13553, 46.12411, 46.11247, 
    46.10059, 46.08848, 46.07614, 46.06357, 46.05077, 46.03773, 46.02447, 
    46.01098, 45.99725, 45.9833, 45.96912, 45.9547, 45.94006, 45.92519, 
    45.9101, 45.89477, 45.87922, 45.86343, 45.84742, 45.83118, 45.81472, 
    45.79803, 45.78111, 45.76396, 45.74659, 45.72899, 45.71117, 45.69312, 
    45.67485, 45.65635, 45.63763, 45.61869, 45.59952, 45.58012, 45.56051, 
    45.54067, 45.52061, 45.50032, 45.47982, 45.45909, 45.43814, 45.41697, 
    45.39558, 45.37397, 45.35214, 45.33009, 45.30782, 45.28534, 45.26263, 
    45.2397, 45.21656, 45.1932, 45.16962, 45.14582, 45.12181, 45.09758, 
    45.07314, 45.04848, 45.0236, 44.99851, 44.97321, 44.94769, 44.92196, 
    44.89602, 44.86986, 44.84349, 44.81691, 44.79011, 44.7631, 44.73589, 
    44.70846, 44.68082, 44.65298, 44.62492, 44.59665, 44.56818, 44.5395, 
    44.51061, 44.48151, 44.45221, 44.4227, 44.39298, 44.36306, 44.33293, 
    44.30259, 44.27206, 44.24131, 44.21037, 44.17922, 44.14787, 44.11632, 
    44.08456, 44.0526, 44.02045, 43.98809, 43.95553, 43.92277, 43.88981, 
    43.85666, 43.8233, 43.78975, 43.756, 43.72205, 43.68791, 43.65357, 
    43.61903, 43.5843, 43.54937, 43.51426, 43.47894, 43.44343, 43.40773, 
    43.37184, 43.33575, 43.29948, 43.26301, 43.22635, 43.1895, 43.15246, 
    43.11523, 43.07782,
  38.94375, 38.99668, 39.04947, 39.10212, 39.15461, 39.20697, 39.25918, 
    39.31124, 39.36315, 39.41492, 39.46654, 39.51801, 39.56933, 39.6205, 
    39.67152, 39.72239, 39.77311, 39.82368, 39.8741, 39.92437, 39.97448, 
    40.02444, 40.07424, 40.12389, 40.17339, 40.22273, 40.27192, 40.32095, 
    40.36982, 40.41853, 40.46709, 40.51549, 40.56373, 40.61181, 40.65973, 
    40.7075, 40.7551, 40.80254, 40.84982, 40.89693, 40.94389, 40.99068, 
    41.03731, 41.08377, 41.13007, 41.17621, 41.22218, 41.26798, 41.31361, 
    41.35909, 41.40439, 41.44952, 41.49449, 41.53929, 41.58392, 41.62837, 
    41.67266, 41.71678, 41.76072, 41.8045, 41.8481, 41.89153, 41.93478, 
    41.97786, 42.02077, 42.0635, 42.10606, 42.14844, 42.19065, 42.23268, 
    42.27453, 42.3162, 42.3577, 42.39902, 42.44016, 42.48111, 42.52189, 
    42.56249, 42.60291, 42.64314, 42.6832, 42.72307, 42.76276, 42.80226, 
    42.84158, 42.88072, 42.91967, 42.95844, 42.99702, 43.03541, 43.07362, 
    43.11164, 43.14947, 43.18711, 43.22457, 43.26184, 43.29892, 43.3358, 
    43.3725, 43.409, 43.44532, 43.48144, 43.51737, 43.5531, 43.58865, 43.624, 
    43.65915, 43.69411, 43.72888, 43.76345, 43.79782, 43.832, 43.86598, 
    43.89977, 43.93335, 43.96674, 43.99993, 44.03292, 44.0657, 44.09829, 
    44.13068, 44.16287, 44.19486, 44.22664, 44.25822, 44.2896, 44.32078, 
    44.35175, 44.38252, 44.41309, 44.44345, 44.4736, 44.50355, 44.53329, 
    44.56283, 44.59216, 44.62128, 44.6502, 44.6789, 44.7074, 44.73569, 
    44.76376, 44.79163, 44.81929, 44.84674, 44.87398, 44.901, 44.92782, 
    44.95442, 44.98081, 45.00699, 45.03295, 45.0587, 45.08424, 45.10956, 
    45.13466, 45.15955, 45.18423, 45.20869, 45.23293, 45.25696, 45.28077, 
    45.30436, 45.32774, 45.35089, 45.37383, 45.39655, 45.41905, 45.44133, 
    45.46339, 45.48523, 45.50685, 45.52825, 45.54943, 45.57038, 45.59112, 
    45.61163, 45.63192, 45.65199, 45.67184, 45.69146, 45.71086, 45.73003, 
    45.74898, 45.7677, 45.78621, 45.80448, 45.82253, 45.84035, 45.85795, 
    45.87532, 45.89247, 45.90939, 45.92607, 45.94254, 45.95877, 45.97478, 
    45.99057, 46.00611, 46.02144, 46.03653, 46.0514, 46.06604, 46.08044, 
    46.09462, 46.10856, 46.12228, 46.13577, 46.14902, 46.16204, 46.17484, 
    46.1874, 46.19973, 46.21183, 46.22369, 46.23533, 46.24673, 46.2579, 
    46.26884, 46.27954, 46.29001, 46.30025, 46.31025, 46.32002, 46.32956, 
    46.33886, 46.34793, 46.35677, 46.36536, 46.37373, 46.38186, 46.38976, 
    46.39742, 46.40485, 46.41204, 46.41899, 46.42572, 46.4322, 46.43845, 
    46.44447, 46.45024, 46.45579, 46.46109, 46.46616, 46.471, 46.4756, 
    46.47996, 46.48409, 46.48797, 46.49163, 46.49504, 46.49822, 46.50116, 
    46.50387, 46.50634, 46.50857, 46.51057, 46.51233, 46.51385, 46.51513, 
    46.51618, 46.51699, 46.51756, 46.5179, 46.518, 46.51786, 46.51749, 
    46.51688, 46.51603, 46.51494, 46.51362, 46.51206, 46.51027, 46.50823, 
    46.50596, 46.50346, 46.50071, 46.49773, 46.49451, 46.49106, 46.48737, 
    46.48345, 46.47928, 46.47488, 46.47025, 46.46538, 46.46027, 46.45493, 
    46.44934, 46.44353, 46.43748, 46.43119, 46.42467, 46.41791, 46.41092, 
    46.40369, 46.39622, 46.38853, 46.38059, 46.37243, 46.36402, 46.35538, 
    46.34651, 46.33741, 46.32806, 46.31849, 46.30869, 46.29865, 46.28837, 
    46.27786, 46.26712, 46.25615, 46.24494, 46.2335, 46.22183, 46.20993, 
    46.1978, 46.18543, 46.17283, 46.16, 46.14694, 46.13365, 46.12012, 
    46.10637, 46.09239, 46.07818, 46.06374, 46.04906, 46.03416, 46.01903, 
    46.00367, 45.98808, 45.97227, 45.95622, 45.93995, 45.92345, 45.90672, 
    45.88977, 45.87259, 45.85518, 45.83755, 45.81969, 45.8016, 45.78329, 
    45.76476, 45.74599, 45.72701, 45.7078, 45.68837, 45.66871, 45.64883, 
    45.62873, 45.6084, 45.58786, 45.56709, 45.54609, 45.52488, 45.50344, 
    45.48179, 45.45992, 45.43782, 45.4155, 45.39297, 45.37022, 45.34724, 
    45.32405, 45.30064, 45.27702, 45.25317, 45.22911, 45.20483, 45.18034, 
    45.15563, 45.13071, 45.10557, 45.08021, 45.05464, 45.02886, 45.00286, 
    44.97665, 44.95023, 44.92359, 44.89674, 44.86969, 44.84241, 44.81493, 
    44.78724, 44.75934, 44.73122, 44.7029, 44.67437, 44.64563, 44.61669, 
    44.58753, 44.55817, 44.5286, 44.49883, 44.46885, 44.43866, 44.40827, 
    44.37767, 44.34687, 44.31586, 44.28465, 44.25324, 44.22163, 44.18981, 
    44.15779, 44.12557, 44.09315, 44.06053, 44.02771, 43.99469, 43.96147, 
    43.92805, 43.89444, 43.86062, 43.82661, 43.7924, 43.758, 43.7234, 
    43.6886, 43.65361, 43.61842, 43.58304, 43.54747, 43.5117, 43.47574, 
    43.43959, 43.40324, 43.36671, 43.32998, 43.29306, 43.25595, 43.21866, 
    43.18118,
  39.04004, 39.09305, 39.14592, 39.19864, 39.25122, 39.30365, 39.35594, 
    39.40808, 39.46008, 39.51192, 39.56362, 39.61517, 39.66657, 39.71782, 
    39.76892, 39.81987, 39.87067, 39.92132, 39.97182, 40.02216, 40.07235, 
    40.12239, 40.17227, 40.222, 40.27158, 40.321, 40.37026, 40.41937, 
    40.46832, 40.51711, 40.56575, 40.61423, 40.66254, 40.7107, 40.75871, 
    40.80655, 40.85423, 40.90174, 40.9491, 40.99629, 41.04332, 41.09019, 
    41.1369, 41.18344, 41.22982, 41.27603, 41.32207, 41.36795, 41.41367, 
    41.45921, 41.50459, 41.5498, 41.59484, 41.63972, 41.68442, 41.72895, 
    41.77332, 41.81751, 41.86153, 41.90538, 41.94906, 41.99256, 42.03589, 
    42.07905, 42.12203, 42.16484, 42.20747, 42.24992, 42.29221, 42.33431, 
    42.37623, 42.41798, 42.45955, 42.50094, 42.54215, 42.58318, 42.62403, 
    42.6647, 42.70519, 42.7455, 42.78563, 42.82557, 42.86533, 42.9049, 
    42.9443, 42.98351, 43.02253, 43.06136, 43.10001, 43.13848, 43.17675, 
    43.21484, 43.25275, 43.29046, 43.32798, 43.36532, 43.40247, 43.43942, 
    43.47618, 43.51276, 43.54914, 43.58533, 43.62133, 43.65713, 43.69274, 
    43.72815, 43.76337, 43.7984, 43.83323, 43.86787, 43.90231, 43.93655, 
    43.9706, 44.00444, 44.03809, 44.07154, 44.10479, 44.13785, 44.1707, 
    44.20335, 44.2358, 44.26805, 44.3001, 44.33195, 44.36359, 44.39503, 
    44.42627, 44.4573, 44.48813, 44.51875, 44.54917, 44.57939, 44.60939, 
    44.63919, 44.66879, 44.69818, 44.72736, 44.75632, 44.78509, 44.81364, 
    44.84199, 44.87012, 44.89804, 44.92576, 44.95326, 44.98056, 45.00764, 
    45.0345, 45.06116, 45.0876, 45.11383, 45.13985, 45.16565, 45.19123, 
    45.21661, 45.24176, 45.2667, 45.29143, 45.31594, 45.34023, 45.36431, 
    45.38816, 45.41181, 45.43523, 45.45843, 45.48142, 45.50418, 45.52673, 
    45.54906, 45.57116, 45.59305, 45.61471, 45.63615, 45.65738, 45.67838, 
    45.69915, 45.71971, 45.74004, 45.76015, 45.78004, 45.7997, 45.81914, 
    45.83835, 45.85734, 45.87611, 45.89465, 45.91296, 45.93105, 45.94891, 
    45.96654, 45.98395, 46.00113, 46.01809, 46.03481, 46.05131, 46.06758, 
    46.08362, 46.09943, 46.11502, 46.13037, 46.1455, 46.1604, 46.17506, 
    46.1895, 46.20371, 46.21769, 46.23143, 46.24495, 46.25823, 46.27128, 
    46.2841, 46.29669, 46.30904, 46.32117, 46.33306, 46.34472, 46.35614, 
    46.36734, 46.3783, 46.38902, 46.39952, 46.40978, 46.4198, 46.4296, 
    46.43915, 46.44847, 46.45756, 46.46642, 46.47504, 46.48342, 46.49157, 
    46.49948, 46.50716, 46.5146, 46.52181, 46.52878, 46.53551, 46.54202, 
    46.54828, 46.55431, 46.5601, 46.56565, 46.57097, 46.57605, 46.58089, 
    46.5855, 46.58987, 46.59401, 46.59791, 46.60157, 46.60499, 46.60818, 
    46.61113, 46.61384, 46.61631, 46.61855, 46.62055, 46.62231, 46.62384, 
    46.62513, 46.62617, 46.62699, 46.62756, 46.6279, 46.628, 46.62786, 
    46.62749, 46.62687, 46.62602, 46.62494, 46.62361, 46.62205, 46.62025, 
    46.61821, 46.61594, 46.61343, 46.61068, 46.60769, 46.60447, 46.60101, 
    46.59731, 46.59337, 46.5892, 46.58479, 46.58015, 46.57526, 46.57014, 
    46.56479, 46.5592, 46.55337, 46.5473, 46.541, 46.53447, 46.52769, 
    46.52068, 46.51344, 46.50596, 46.49825, 46.4903, 46.48211, 46.47369, 
    46.46503, 46.45614, 46.44701, 46.43766, 46.42806, 46.41823, 46.40817, 
    46.39787, 46.38734, 46.37658, 46.36558, 46.35435, 46.34289, 46.3312, 
    46.31927, 46.30711, 46.29471, 46.28209, 46.26923, 46.25614, 46.24282, 
    46.22927, 46.21549, 46.20148, 46.18723, 46.17276, 46.15806, 46.14312, 
    46.12796, 46.11257, 46.09695, 46.0811, 46.06502, 46.04871, 46.03218, 
    46.01542, 45.99843, 45.98121, 45.96377, 45.94609, 45.9282, 45.91008, 
    45.89173, 45.87315, 45.85435, 45.83533, 45.81608, 45.7966, 45.77691, 
    45.75699, 45.73684, 45.71647, 45.69588, 45.67507, 45.65403, 45.63278, 
    45.6113, 45.5896, 45.56768, 45.54554, 45.52318, 45.5006, 45.47779, 
    45.45478, 45.43154, 45.40808, 45.38441, 45.36052, 45.3364, 45.31208, 
    45.28753, 45.26278, 45.2378, 45.21261, 45.1872, 45.16158, 45.13575, 
    45.1097, 45.08343, 45.05696, 45.03027, 45.00336, 44.97625, 44.94893, 
    44.92139, 44.89364, 44.86568, 44.83752, 44.80914, 44.78055, 44.75176, 
    44.72275, 44.69354, 44.66412, 44.63449, 44.60466, 44.57462, 44.54437, 
    44.51392, 44.48326, 44.4524, 44.42134, 44.39007, 44.3586, 44.32692, 
    44.29504, 44.26296, 44.23068, 44.1982, 44.16552, 44.13263, 44.09955, 
    44.06627, 44.03278, 43.9991, 43.96522, 43.93115, 43.89687, 43.8624, 
    43.82774, 43.79287, 43.75782, 43.72256, 43.68712, 43.65148, 43.61564, 
    43.57962, 43.5434, 43.50698, 43.47038, 43.43359, 43.3966, 43.35942, 
    43.32206, 43.28451,
  39.13628, 39.18938, 39.24232, 39.29513, 39.34779, 39.4003, 39.45267, 
    39.50489, 39.55696, 39.60889, 39.66066, 39.71229, 39.76377, 39.8151, 
    39.86628, 39.91731, 39.96819, 40.01892, 40.06949, 40.11992, 40.17019, 
    40.2203, 40.27027, 40.32008, 40.36973, 40.41923, 40.46857, 40.51775, 
    40.56678, 40.61566, 40.66437, 40.71293, 40.76133, 40.80956, 40.85764, 
    40.90556, 40.95332, 41.00091, 41.04835, 41.09562, 41.14273, 41.18967, 
    41.23646, 41.28307, 41.32953, 41.37582, 41.42194, 41.4679, 41.51369, 
    41.55931, 41.60476, 41.65005, 41.69517, 41.74012, 41.7849, 41.82951, 
    41.87395, 41.91822, 41.96231, 42.00624, 42.04999, 42.09357, 42.13697, 
    42.1802, 42.22326, 42.26614, 42.30885, 42.35138, 42.39373, 42.43591, 
    42.47791, 42.51973, 42.56137, 42.60283, 42.64412, 42.68522, 42.72615, 
    42.76689, 42.80745, 42.84783, 42.88803, 42.92804, 42.96787, 43.00752, 
    43.04699, 43.08626, 43.12535, 43.16426, 43.20298, 43.24152, 43.27987, 
    43.31802, 43.356, 43.39378, 43.43137, 43.46878, 43.50599, 43.54301, 
    43.57985, 43.61649, 43.65294, 43.68919, 43.72526, 43.76113, 43.79681, 
    43.83229, 43.86758, 43.90267, 43.93756, 43.97227, 44.00677, 44.04108, 
    44.07519, 44.1091, 44.14281, 44.17633, 44.20964, 44.24276, 44.27567, 
    44.30839, 44.3409, 44.37321, 44.40532, 44.43723, 44.46894, 44.50044, 
    44.53174, 44.56283, 44.59372, 44.6244, 44.65488, 44.68515, 44.71522, 
    44.74508, 44.77473, 44.80418, 44.83342, 44.86244, 44.89126, 44.91987, 
    44.94827, 44.97646, 45.00444, 45.03222, 45.05977, 45.08712, 45.11425, 
    45.14117, 45.16788, 45.19438, 45.22066, 45.24673, 45.27258, 45.29822, 
    45.32365, 45.34885, 45.37384, 45.39862, 45.42318, 45.44752, 45.47165, 
    45.49555, 45.51924, 45.54271, 45.56596, 45.589, 45.61181, 45.6344, 
    45.65677, 45.67892, 45.70086, 45.72256, 45.74405, 45.76532, 45.78636, 
    45.80718, 45.82778, 45.84816, 45.86831, 45.88823, 45.90794, 45.92741, 
    45.94667, 45.9657, 45.9845, 46.00308, 46.02143, 46.03955, 46.05745, 
    46.07513, 46.09257, 46.10979, 46.12678, 46.14354, 46.16007, 46.17638, 
    46.19246, 46.2083, 46.22392, 46.23931, 46.25446, 46.26939, 46.28409, 
    46.29856, 46.31279, 46.3268, 46.34058, 46.35412, 46.36743, 46.38051, 
    46.39336, 46.40597, 46.41835, 46.43051, 46.44242, 46.45411, 46.46556, 
    46.47678, 46.48776, 46.49851, 46.50903, 46.51931, 46.52935, 46.53917, 
    46.54874, 46.55809, 46.56719, 46.57607, 46.58471, 46.59311, 46.60127, 
    46.6092, 46.6169, 46.62436, 46.63158, 46.63857, 46.64532, 46.65183, 
    46.65811, 46.66415, 46.66995, 46.67552, 46.68085, 46.68594, 46.69079, 
    46.69541, 46.69979, 46.70394, 46.70784, 46.71151, 46.71494, 46.71814, 
    46.72109, 46.72381, 46.72629, 46.72853, 46.73053, 46.7323, 46.73383, 
    46.73512, 46.73617, 46.73698, 46.73756, 46.7379, 46.738, 46.73786, 
    46.73748, 46.73687, 46.73602, 46.73493, 46.7336, 46.73204, 46.73023, 
    46.72819, 46.72591, 46.72339, 46.72064, 46.71764, 46.71441, 46.71095, 
    46.70724, 46.7033, 46.69912, 46.6947, 46.69004, 46.68515, 46.68002, 
    46.67465, 46.66905, 46.66321, 46.65713, 46.65081, 46.64426, 46.63748, 
    46.63045, 46.62319, 46.6157, 46.60796, 46.59999, 46.59179, 46.58335, 
    46.57468, 46.56577, 46.55662, 46.54725, 46.53763, 46.52778, 46.5177, 
    46.50738, 46.49682, 46.48604, 46.47502, 46.46376, 46.45227, 46.44055, 
    46.4286, 46.41641, 46.40399, 46.39134, 46.37846, 46.36534, 46.35199, 
    46.33841, 46.3246, 46.31056, 46.29628, 46.28178, 46.26705, 46.25208, 
    46.23689, 46.22146, 46.20581, 46.18993, 46.17381, 46.15747, 46.1409, 
    46.12411, 46.10708, 46.08983, 46.07235, 46.05464, 46.03671, 46.01854, 
    46.00016, 45.98154, 45.9627, 45.94364, 45.92435, 45.90483, 45.8851, 
    45.86514, 45.84495, 45.82454, 45.80391, 45.78305, 45.76197, 45.74067, 
    45.71915, 45.6974, 45.67543, 45.65325, 45.63084, 45.60822, 45.58537, 
    45.5623, 45.53901, 45.51551, 45.49179, 45.46785, 45.44369, 45.41931, 
    45.39471, 45.36991, 45.34488, 45.31964, 45.29418, 45.26851, 45.24262, 
    45.21652, 45.1902, 45.16367, 45.13693, 45.10997, 45.08281, 45.05543, 
    45.02784, 45.00003, 44.97202, 44.94379, 44.91536, 44.88672, 44.85786, 
    44.8288, 44.79953, 44.77006, 44.74037, 44.71048, 44.68038, 44.65007, 
    44.61956, 44.58885, 44.55793, 44.5268, 44.49547, 44.46394, 44.4322, 
    44.40026, 44.36812, 44.33577, 44.30323, 44.27048, 44.23753, 44.20439, 
    44.17104, 44.13749, 44.10375, 44.06981, 44.03566, 44.00133, 43.96679, 
    43.93206, 43.89713, 43.86201, 43.82669, 43.79118, 43.75547, 43.71957, 
    43.68347, 43.64719, 43.61071, 43.57404, 43.53717, 43.50012, 43.46287, 
    43.42544, 43.38782,
  39.23249, 39.28566, 39.33869, 39.39157, 39.44431, 39.49691, 39.54935, 
    39.60165, 39.6538, 39.70581, 39.75767, 39.80938, 39.86094, 39.91235, 
    39.9636, 40.01471, 40.06567, 40.11648, 40.16713, 40.21764, 40.26799, 
    40.31818, 40.36822, 40.41811, 40.46784, 40.51742, 40.56684, 40.61611, 
    40.66521, 40.71416, 40.76296, 40.81159, 40.86007, 40.90839, 40.95654, 
    41.00454, 41.05237, 41.10005, 41.14756, 41.19491, 41.2421, 41.28912, 
    41.33598, 41.38268, 41.42921, 41.47557, 41.52177, 41.56781, 41.61367, 
    41.65937, 41.70491, 41.75027, 41.79546, 41.84049, 41.88535, 41.93003, 
    41.97454, 42.01889, 42.06306, 42.10706, 42.15089, 42.19454, 42.23802, 
    42.28133, 42.32446, 42.36742, 42.4102, 42.4528, 42.49523, 42.53748, 
    42.57956, 42.62145, 42.66317, 42.7047, 42.74606, 42.78724, 42.82823, 
    42.86905, 42.90968, 42.95013, 42.99041, 43.03049, 43.07039, 43.11012, 
    43.14965, 43.189, 43.22816, 43.26714, 43.30593, 43.34454, 43.38295, 
    43.42118, 43.45922, 43.49708, 43.53474, 43.57221, 43.6095, 43.64659, 
    43.68349, 43.7202, 43.75671, 43.79304, 43.82917, 43.86511, 43.90085, 
    43.9364, 43.97176, 44.00692, 44.04188, 44.07664, 44.11121, 44.14559, 
    44.17976, 44.21374, 44.24752, 44.28109, 44.31447, 44.34765, 44.38063, 
    44.41341, 44.44598, 44.47836, 44.51053, 44.5425, 44.57427, 44.60583, 
    44.63719, 44.66834, 44.69929, 44.73004, 44.76057, 44.79091, 44.82103, 
    44.85095, 44.88066, 44.91016, 44.93946, 44.96854, 44.99742, 45.02609, 
    45.05455, 45.08279, 45.11083, 45.13865, 45.16627, 45.19367, 45.22086, 
    45.24783, 45.2746, 45.30114, 45.32748, 45.3536, 45.37951, 45.4052, 
    45.43067, 45.45593, 45.48097, 45.5058, 45.53041, 45.5548, 45.57898, 
    45.60293, 45.62667, 45.65018, 45.67348, 45.69656, 45.71942, 45.74206, 
    45.76448, 45.78668, 45.80865, 45.83041, 45.85194, 45.87325, 45.89434, 
    45.9152, 45.93584, 45.95626, 45.97645, 45.99642, 46.01617, 46.03569, 
    46.05498, 46.07405, 46.09289, 46.11151, 46.1299, 46.14806, 46.166, 
    46.18371, 46.20119, 46.21844, 46.23547, 46.25226, 46.26883, 46.28517, 
    46.30128, 46.31716, 46.33281, 46.34823, 46.36342, 46.37838, 46.39311, 
    46.40761, 46.42188, 46.43591, 46.44972, 46.46329, 46.47663, 46.48974, 
    46.50261, 46.51525, 46.52766, 46.53984, 46.55178, 46.56349, 46.57497, 
    46.58621, 46.59722, 46.60799, 46.61853, 46.62883, 46.6389, 46.64874, 
    46.65833, 46.66769, 46.67682, 46.68571, 46.69437, 46.70279, 46.71098, 
    46.71892, 46.72663, 46.73411, 46.74135, 46.74835, 46.75512, 46.76164, 
    46.76793, 46.77399, 46.7798, 46.78538, 46.79072, 46.79583, 46.80069, 
    46.80532, 46.80971, 46.81386, 46.81778, 46.82145, 46.82489, 46.82809, 
    46.83105, 46.83377, 46.83626, 46.83851, 46.84052, 46.84229, 46.84382, 
    46.84511, 46.84616, 46.84698, 46.84756, 46.8479, 46.848, 46.84786, 
    46.84748, 46.84687, 46.84602, 46.84492, 46.84359, 46.84202, 46.84021, 
    46.83817, 46.83588, 46.83336, 46.8306, 46.8276, 46.82436, 46.82089, 
    46.81717, 46.81322, 46.80903, 46.8046, 46.79994, 46.79503, 46.78989, 
    46.78452, 46.7789, 46.77304, 46.76695, 46.76062, 46.75406, 46.74726, 
    46.74022, 46.73294, 46.72543, 46.71768, 46.7097, 46.70147, 46.69302, 
    46.68432, 46.6754, 46.66623, 46.65683, 46.64719, 46.63732, 46.62722, 
    46.61687, 46.6063, 46.59549, 46.58445, 46.57317, 46.56166, 46.54991, 
    46.53793, 46.52572, 46.51327, 46.50059, 46.48768, 46.47454, 46.46116, 
    46.44755, 46.43371, 46.41964, 46.40533, 46.3908, 46.37603, 46.36104, 
    46.34581, 46.33035, 46.31467, 46.29875, 46.2826, 46.26623, 46.24962, 
    46.23279, 46.21573, 46.19844, 46.18092, 46.16317, 46.1452, 46.127, 
    46.10858, 46.08992, 46.07105, 46.05194, 46.03261, 46.01306, 45.99328, 
    45.97327, 45.95304, 45.93259, 45.91191, 45.89102, 45.8699, 45.84855, 
    45.82698, 45.80519, 45.78318, 45.76095, 45.73849, 45.71582, 45.69293, 
    45.66982, 45.64648, 45.62293, 45.59916, 45.57516, 45.55096, 45.52653, 
    45.50189, 45.47703, 45.45195, 45.42665, 45.40115, 45.37542, 45.34948, 
    45.32333, 45.29696, 45.27038, 45.24358, 45.21657, 45.18935, 45.16191, 
    45.13427, 45.10641, 45.07834, 45.05006, 45.02157, 44.99287, 44.96396, 
    44.93484, 44.90551, 44.87598, 44.84623, 44.81628, 44.78612, 44.75576, 
    44.72519, 44.69441, 44.66343, 44.63224, 44.60085, 44.56926, 44.53746, 
    44.50546, 44.47325, 44.44085, 44.40824, 44.37543, 44.34242, 44.30921, 
    44.27579, 44.24218, 44.20838, 44.17437, 44.14016, 44.10576, 44.07116, 
    44.03636, 44.00137, 43.96618, 43.93079, 43.89521, 43.85944, 43.82347, 
    43.78731, 43.75095, 43.71441, 43.67767, 43.64073, 43.60361, 43.5663, 
    43.52879, 43.4911,
  39.32866, 39.38191, 39.43502, 39.48798, 39.5408, 39.59347, 39.646, 
    39.69838, 39.75061, 39.8027, 39.85463, 39.90642, 39.95806, 40.00955, 
    40.06089, 40.11208, 40.16312, 40.214, 40.26474, 40.31532, 40.36575, 
    40.41602, 40.46614, 40.51611, 40.56592, 40.61558, 40.66508, 40.71442, 
    40.76361, 40.81264, 40.86151, 40.91022, 40.95878, 41.00717, 41.05541, 
    41.10348, 41.15139, 41.19915, 41.24674, 41.29417, 41.34143, 41.38853, 
    41.43547, 41.48224, 41.52885, 41.57529, 41.62157, 41.66768, 41.71363, 
    41.7594, 41.80501, 41.85045, 41.89573, 41.94083, 41.98576, 42.03052, 
    42.07511, 42.11953, 42.16378, 42.20786, 42.25176, 42.29549, 42.33904, 
    42.38243, 42.42563, 42.46866, 42.51152, 42.5542, 42.5967, 42.63903, 
    42.68117, 42.72314, 42.76493, 42.80654, 42.84797, 42.88922, 42.93029, 
    42.97118, 43.01189, 43.05241, 43.09275, 43.13291, 43.17289, 43.21268, 
    43.25229, 43.29171, 43.33094, 43.36999, 43.40885, 43.44753, 43.48602, 
    43.52431, 43.56243, 43.60035, 43.63808, 43.67562, 43.71297, 43.75014, 
    43.78711, 43.82388, 43.86047, 43.89686, 43.93306, 43.96907, 44.00488, 
    44.04049, 44.07591, 44.11114, 44.14617, 44.181, 44.21564, 44.25008, 
    44.28431, 44.31836, 44.3522, 44.38584, 44.41928, 44.45253, 44.48557, 
    44.51841, 44.55105, 44.58348, 44.61572, 44.64775, 44.67958, 44.7112, 
    44.74263, 44.77384, 44.80485, 44.83566, 44.86625, 44.89664, 44.92683, 
    44.95681, 44.98658, 45.01614, 45.04549, 45.07463, 45.10357, 45.13229, 
    45.1608, 45.18911, 45.2172, 45.24508, 45.27275, 45.30021, 45.32745, 
    45.35448, 45.38129, 45.4079, 45.43428, 45.46046, 45.48642, 45.51216, 
    45.53769, 45.563, 45.58809, 45.61297, 45.63763, 45.66207, 45.68629, 
    45.7103, 45.73408, 45.75765, 45.78099, 45.80412, 45.82703, 45.84972, 
    45.87218, 45.89442, 45.91644, 45.93824, 45.95982, 45.98117, 46.0023, 
    46.02321, 46.0439, 46.06436, 46.08459, 46.1046, 46.12439, 46.14395, 
    46.16328, 46.18239, 46.20127, 46.21993, 46.23836, 46.25656, 46.27453, 
    46.29228, 46.3098, 46.32709, 46.34415, 46.36098, 46.37759, 46.39396, 
    46.4101, 46.42602, 46.4417, 46.45716, 46.47238, 46.48737, 46.50213, 
    46.51666, 46.53096, 46.54502, 46.55886, 46.57246, 46.58583, 46.59896, 
    46.61187, 46.62453, 46.63697, 46.64917, 46.66114, 46.67287, 46.68438, 
    46.69564, 46.70667, 46.71747, 46.72803, 46.73835, 46.74845, 46.7583, 
    46.76792, 46.7773, 46.78645, 46.79536, 46.80404, 46.81248, 46.82068, 
    46.82864, 46.83637, 46.84386, 46.85112, 46.85813, 46.86491, 46.87145, 
    46.87776, 46.88382, 46.88965, 46.89524, 46.9006, 46.90571, 46.91059, 
    46.91523, 46.91962, 46.92379, 46.92771, 46.9314, 46.93484, 46.93805, 
    46.94102, 46.94374, 46.94624, 46.94849, 46.9505, 46.95227, 46.95381, 
    46.9551, 46.95616, 46.95698, 46.95756, 46.9579, 46.958, 46.95786, 
    46.95749, 46.95687, 46.95601, 46.95492, 46.95358, 46.95201, 46.9502, 
    46.94815, 46.94586, 46.94333, 46.94056, 46.93756, 46.93431, 46.93083, 
    46.9271, 46.92315, 46.91895, 46.91451, 46.90983, 46.90492, 46.89977, 
    46.89437, 46.88875, 46.88288, 46.87678, 46.87043, 46.86385, 46.85704, 
    46.84998, 46.84269, 46.83516, 46.8274, 46.8194, 46.81116, 46.80268, 
    46.79397, 46.78502, 46.77584, 46.76641, 46.75676, 46.74686, 46.73674, 
    46.72638, 46.71578, 46.70494, 46.69387, 46.68257, 46.67104, 46.65926, 
    46.64726, 46.63502, 46.62255, 46.60984, 46.5969, 46.58373, 46.57032, 
    46.55669, 46.54282, 46.52871, 46.51438, 46.49981, 46.48502, 46.46999, 
    46.45473, 46.43924, 46.42352, 46.40757, 46.39138, 46.37497, 46.35833, 
    46.34146, 46.32437, 46.30704, 46.28949, 46.27171, 46.2537, 46.23546, 
    46.217, 46.1983, 46.17938, 46.16024, 46.14087, 46.12127, 46.10145, 
    46.08141, 46.06113, 46.04064, 46.01992, 45.99898, 45.97781, 45.95642, 
    45.93481, 45.91298, 45.89092, 45.86864, 45.84614, 45.82342, 45.80048, 
    45.77732, 45.75394, 45.73034, 45.70651, 45.68248, 45.65822, 45.63374, 
    45.60905, 45.58414, 45.55901, 45.53366, 45.5081, 45.48233, 45.45633, 
    45.43013, 45.40371, 45.37707, 45.35022, 45.32315, 45.29588, 45.26839, 
    45.24068, 45.21277, 45.18465, 45.15631, 45.12776, 45.099, 45.07004, 
    45.04086, 45.01147, 44.98188, 44.95208, 44.92207, 44.89185, 44.86143, 
    44.8308, 44.79996, 44.76892, 44.73767, 44.70621, 44.67456, 44.6427, 
    44.61063, 44.57837, 44.5459, 44.51323, 44.48035, 44.44728, 44.41401, 
    44.38053, 44.34686, 44.31298, 44.27891, 44.24464, 44.21017, 44.1755, 
    44.14064, 44.10558, 44.07032, 44.03487, 43.99923, 43.96338, 43.92735, 
    43.89112, 43.85469, 43.81808, 43.78127, 43.74427, 43.70708, 43.6697, 
    43.63213, 43.59436,
  39.42478, 39.47812, 39.5313, 39.58435, 39.63725, 39.69, 39.7426, 39.79506, 
    39.84738, 39.89954, 39.95156, 40.00343, 40.05515, 40.10672, 40.15813, 
    40.2094, 40.26052, 40.31149, 40.3623, 40.41296, 40.46347, 40.51382, 
    40.56403, 40.61407, 40.66396, 40.7137, 40.76328, 40.8127, 40.86197, 
    40.91108, 40.96003, 41.00882, 41.05745, 41.10592, 41.15424, 41.20239, 
    41.25038, 41.29821, 41.34588, 41.39339, 41.44073, 41.48791, 41.53493, 
    41.58178, 41.62846, 41.67498, 41.72134, 41.76753, 41.81355, 41.8594, 
    41.90509, 41.95061, 41.99596, 42.04113, 42.08614, 42.13098, 42.17565, 
    42.22015, 42.26447, 42.30862, 42.3526, 42.3964, 42.44004, 42.48349, 
    42.52678, 42.56988, 42.61281, 42.65556, 42.69814, 42.74054, 42.78276, 
    42.82481, 42.86667, 42.90835, 42.94986, 42.99118, 43.03233, 43.07329, 
    43.11407, 43.15466, 43.19508, 43.23531, 43.27536, 43.31522, 43.3549, 
    43.39439, 43.4337, 43.47282, 43.51175, 43.5505, 43.58905, 43.62743, 
    43.66561, 43.7036, 43.7414, 43.77901, 43.81643, 43.85366, 43.8907, 
    43.92755, 43.9642, 44.00066, 44.03693, 44.073, 44.10888, 44.14457, 
    44.18005, 44.21534, 44.25044, 44.28534, 44.32004, 44.35454, 44.38885, 
    44.42295, 44.45686, 44.49057, 44.52407, 44.55738, 44.59049, 44.62339, 
    44.65609, 44.68859, 44.72089, 44.75299, 44.78488, 44.81656, 44.84805, 
    44.87932, 44.91039, 44.94125, 44.97191, 45.00237, 45.03261, 45.06264, 
    45.09247, 45.12209, 45.1515, 45.18071, 45.2097, 45.23848, 45.26705, 
    45.29541, 45.32356, 45.35149, 45.37922, 45.40673, 45.43403, 45.46111, 
    45.48798, 45.51464, 45.54108, 45.56731, 45.59332, 45.61911, 45.64469, 
    45.67005, 45.6952, 45.72013, 45.74483, 45.76933, 45.7936, 45.81765, 
    45.84149, 45.8651, 45.8885, 45.91167, 45.93463, 45.95736, 45.97987, 
    46.00216, 46.02423, 46.04607, 46.06769, 46.08909, 46.11027, 46.13122, 
    46.15194, 46.17245, 46.19272, 46.21278, 46.2326, 46.2522, 46.27158, 
    46.29073, 46.30965, 46.32835, 46.34681, 46.36505, 46.38306, 46.40085, 
    46.4184, 46.43573, 46.45283, 46.4697, 46.48634, 46.50274, 46.51892, 
    46.53487, 46.55059, 46.56607, 46.58133, 46.59636, 46.61115, 46.62571, 
    46.64003, 46.65413, 46.668, 46.68163, 46.69502, 46.70818, 46.72112, 
    46.73381, 46.74627, 46.7585, 46.7705, 46.78226, 46.79378, 46.80507, 
    46.81613, 46.82695, 46.83753, 46.84788, 46.85799, 46.86787, 46.87751, 
    46.88691, 46.89608, 46.90501, 46.9137, 46.92216, 46.93038, 46.93836, 
    46.94611, 46.95361, 46.96088, 46.96791, 46.97471, 46.98127, 46.98758, 
    46.99366, 46.9995, 47.00511, 47.01047, 47.0156, 47.02048, 47.02513, 
    47.02954, 47.03371, 47.03764, 47.04134, 47.04479, 47.048, 47.05098, 
    47.05371, 47.05621, 47.05847, 47.06049, 47.06226, 47.0638, 47.0651, 
    47.06616, 47.06698, 47.06756, 47.0679, 47.068, 47.06786, 47.06748, 
    47.06686, 47.06601, 47.06491, 47.06357, 47.062, 47.06018, 47.05812, 
    47.05583, 47.0533, 47.05053, 47.04751, 47.04426, 47.04077, 47.03704, 
    47.03307, 47.02886, 47.02441, 47.01973, 47.0148, 47.00964, 47.00424, 
    46.9986, 46.99272, 46.9866, 46.98024, 46.97365, 46.96682, 46.95975, 
    46.95244, 46.9449, 46.93711, 46.92909, 46.92084, 46.91234, 46.90361, 
    46.89464, 46.88544, 46.876, 46.86632, 46.85641, 46.84626, 46.83587, 
    46.82525, 46.81439, 46.8033, 46.79197, 46.78041, 46.76862, 46.75658, 
    46.74432, 46.73182, 46.71909, 46.70612, 46.69292, 46.67949, 46.66582, 
    46.65192, 46.63778, 46.62342, 46.60882, 46.59399, 46.57893, 46.56364, 
    46.54812, 46.53236, 46.51638, 46.50016, 46.48372, 46.46704, 46.45014, 
    46.43301, 46.41564, 46.39805, 46.38023, 46.36218, 46.34391, 46.32541, 
    46.30667, 46.28772, 46.26853, 46.24912, 46.22948, 46.20962, 46.18953, 
    46.16922, 46.14868, 46.12792, 46.10693, 46.08572, 46.06429, 46.04263, 
    46.02075, 45.99865, 45.97632, 45.95378, 45.93101, 45.90802, 45.88481, 
    45.86138, 45.83773, 45.81386, 45.78978, 45.76547, 45.74094, 45.7162, 
    45.69123, 45.66605, 45.64066, 45.61505, 45.58922, 45.56317, 45.53691, 
    45.51044, 45.48375, 45.45684, 45.42972, 45.40239, 45.37485, 45.34709, 
    45.31912, 45.29094, 45.26254, 45.23394, 45.20512, 45.1761, 45.14687, 
    45.11742, 45.08777, 45.05791, 45.02784, 44.99756, 44.96708, 44.93639, 
    44.90549, 44.87439, 44.84308, 44.81157, 44.77985, 44.74792, 44.7158, 
    44.68347, 44.65094, 44.6182, 44.58527, 44.55213, 44.51879, 44.48525, 
    44.45151, 44.41757, 44.38343, 44.3491, 44.31456, 44.27983, 44.2449, 
    44.20977, 44.17445, 44.13893, 44.10322, 44.06731, 44.0312, 43.99491, 
    43.95842, 43.92173, 43.88486, 43.84779, 43.81053, 43.77308, 43.73543, 
    43.6976,
  39.52087, 39.57428, 39.62755, 39.68067, 39.73365, 39.78648, 39.83917, 
    39.89171, 39.9441, 39.99635, 40.04844, 40.10039, 40.15219, 40.20384, 
    40.25534, 40.30669, 40.35789, 40.40893, 40.45982, 40.51057, 40.56115, 
    40.61159, 40.66187, 40.71199, 40.76197, 40.81178, 40.86144, 40.91094, 
    40.96029, 41.00948, 41.05851, 41.10738, 41.15609, 41.20464, 41.25303, 
    41.30127, 41.34933, 41.39724, 41.44499, 41.49258, 41.54, 41.58725, 
    41.63435, 41.68128, 41.72804, 41.77464, 41.82107, 41.86734, 41.91344, 
    41.95937, 42.00513, 42.05073, 42.09615, 42.14141, 42.18649, 42.23141, 
    42.27615, 42.32072, 42.36512, 42.40935, 42.45341, 42.49729, 42.541, 
    42.58453, 42.62788, 42.67107, 42.71407, 42.7569, 42.79955, 42.84203, 
    42.88432, 42.92644, 42.96838, 43.01014, 43.05172, 43.09311, 43.13433, 
    43.17537, 43.21622, 43.25689, 43.29737, 43.33768, 43.3778, 43.41773, 
    43.45748, 43.49705, 43.53643, 43.57562, 43.61462, 43.65344, 43.69207, 
    43.73051, 43.76876, 43.80682, 43.8447, 43.88238, 43.91987, 43.95716, 
    43.99427, 44.03119, 44.06791, 44.10444, 44.14077, 44.17691, 44.21286, 
    44.24861, 44.28417, 44.31953, 44.35469, 44.38965, 44.42442, 44.45899, 
    44.49336, 44.52753, 44.5615, 44.59528, 44.62885, 44.66222, 44.69539, 
    44.72836, 44.76112, 44.79369, 44.82605, 44.8582, 44.89016, 44.9219, 
    44.95345, 44.98478, 45.01591, 45.04684, 45.07756, 45.10807, 45.13837, 
    45.16847, 45.19836, 45.22803, 45.2575, 45.28676, 45.31581, 45.34465, 
    45.37328, 45.4017, 45.4299, 45.45789, 45.48567, 45.51324, 45.54059, 
    45.56773, 45.59466, 45.62137, 45.64786, 45.67414, 45.70021, 45.72605, 
    45.75168, 45.7771, 45.80229, 45.82727, 45.85203, 45.87657, 45.90089, 
    45.925, 45.94888, 45.97255, 45.99599, 46.01921, 46.04221, 46.06499, 
    46.08755, 46.10989, 46.132, 46.15389, 46.17556, 46.197, 46.21822, 
    46.23921, 46.25998, 46.28053, 46.30085, 46.32094, 46.34081, 46.36045, 
    46.37987, 46.39906, 46.41802, 46.43676, 46.45526, 46.47354, 46.49159, 
    46.50941, 46.527, 46.54437, 46.5615, 46.57841, 46.59508, 46.61152, 
    46.62774, 46.64372, 46.65947, 46.67499, 46.69028, 46.70533, 46.72016, 
    46.73475, 46.74911, 46.76323, 46.77713, 46.79079, 46.80421, 46.81741, 
    46.83036, 46.84309, 46.85558, 46.86783, 46.87985, 46.89164, 46.90319, 
    46.9145, 46.92558, 46.93642, 46.94703, 46.9574, 46.96753, 46.97743, 
    46.98709, 46.99651, 47.0057, 47.01465, 47.02337, 47.03184, 47.04008, 
    47.04808, 47.05584, 47.06336, 47.07065, 47.07769, 47.0845, 47.09108, 
    47.09741, 47.1035, 47.10935, 47.11497, 47.12035, 47.12548, 47.13038, 
    47.13504, 47.13946, 47.14364, 47.14758, 47.15128, 47.15474, 47.15796, 
    47.16094, 47.16368, 47.16618, 47.16845, 47.17047, 47.17225, 47.17379, 
    47.17509, 47.17616, 47.17698, 47.17756, 47.1779, 47.178, 47.17786, 
    47.17748, 47.17686, 47.176, 47.1749, 47.17356, 47.17198, 47.17016, 
    47.16811, 47.16581, 47.16327, 47.16048, 47.15747, 47.15421, 47.15071, 
    47.14697, 47.14299, 47.13877, 47.13432, 47.12962, 47.12469, 47.11951, 
    47.1141, 47.10844, 47.10255, 47.09642, 47.09005, 47.08344, 47.0766, 
    47.06951, 47.06219, 47.05463, 47.04683, 47.03879, 47.03051, 47.022, 
    47.01325, 47.00426, 46.99504, 46.98558, 46.97588, 46.96595, 46.95577, 
    46.94537, 46.93472, 46.92384, 46.91272, 46.90137, 46.88979, 46.87796, 
    46.86591, 46.85361, 46.84109, 46.82833, 46.81533, 46.8021, 46.78864, 
    46.77494, 46.76101, 46.74685, 46.73246, 46.71783, 46.70297, 46.68787, 
    46.67255, 46.65699, 46.6412, 46.62519, 46.60894, 46.59246, 46.57575, 
    46.55881, 46.54164, 46.52424, 46.50661, 46.48875, 46.47066, 46.45235, 
    46.43381, 46.41504, 46.39604, 46.37681, 46.35736, 46.33768, 46.31778, 
    46.29765, 46.27729, 46.25671, 46.23591, 46.21488, 46.19362, 46.17214, 
    46.15044, 46.12852, 46.10637, 46.084, 46.06141, 46.03859, 46.01555, 
    45.99229, 45.96882, 45.94512, 45.9212, 45.89706, 45.87271, 45.84813, 
    45.82333, 45.79832, 45.77309, 45.74764, 45.72198, 45.6961, 45.67, 
    45.64368, 45.61716, 45.59041, 45.56345, 45.53628, 45.50889, 45.48129, 
    45.45348, 45.42545, 45.39722, 45.36877, 45.3401, 45.31123, 45.28215, 
    45.25286, 45.22335, 45.19364, 45.16372, 45.13359, 45.10326, 45.07271, 
    45.04196, 45.011, 44.97984, 44.94847, 44.91689, 44.88511, 44.85313, 
    44.82094, 44.78855, 44.75595, 44.72316, 44.69016, 44.65696, 44.62355, 
    44.58995, 44.55614, 44.52214, 44.48794, 44.45353, 44.41893, 44.38414, 
    44.34914, 44.31395, 44.27856, 44.24297, 44.20719, 44.17121, 44.13504, 
    44.09867, 44.06211, 44.02536, 43.98842, 43.95128, 43.91395, 43.87643, 
    43.83872, 43.80082,
  39.61691, 39.6704, 39.72375, 39.77695, 39.83001, 39.88293, 39.9357, 
    39.98832, 40.04079, 40.09311, 40.14529, 40.19732, 40.2492, 40.30093, 
    40.35251, 40.40393, 40.45521, 40.50634, 40.55731, 40.60814, 40.6588, 
    40.70932, 40.75967, 40.80988, 40.85993, 40.90982, 40.95956, 41.00915, 
    41.05857, 41.10784, 41.15695, 41.2059, 41.25469, 41.30332, 41.35179, 
    41.4001, 41.44825, 41.49624, 41.54406, 41.59173, 41.63923, 41.68657, 
    41.73373, 41.78074, 41.82759, 41.87426, 41.92077, 41.96712, 42.01329, 
    42.0593, 42.10514, 42.15081, 42.19632, 42.24165, 42.28681, 42.3318, 
    42.37663, 42.42127, 42.46575, 42.51006, 42.55418, 42.59814, 42.64193, 
    42.68553, 42.72897, 42.77222, 42.8153, 42.85821, 42.90094, 42.94349, 
    42.98586, 43.02805, 43.07006, 43.11189, 43.15355, 43.19501, 43.23631, 
    43.27741, 43.31834, 43.35909, 43.39964, 43.44002, 43.48021, 43.52022, 
    43.56004, 43.59968, 43.63913, 43.67839, 43.71747, 43.75636, 43.79506, 
    43.83357, 43.87189, 43.91002, 43.94796, 43.98572, 44.02328, 44.06065, 
    44.09782, 44.13481, 44.1716, 44.20819, 44.2446, 44.28081, 44.31682, 
    44.35264, 44.38826, 44.42369, 44.45892, 44.49395, 44.52878, 44.56342, 
    44.59785, 44.63209, 44.66613, 44.69997, 44.7336, 44.76704, 44.80027, 
    44.8333, 44.86613, 44.89876, 44.93118, 44.9634, 44.99541, 45.02723, 
    45.05883, 45.09023, 45.12142, 45.15241, 45.18319, 45.21376, 45.24412, 
    45.27428, 45.30422, 45.33396, 45.36349, 45.39281, 45.42191, 45.45081, 
    45.4795, 45.50797, 45.53623, 45.56428, 45.59211, 45.61974, 45.64714, 
    45.67434, 45.70132, 45.72808, 45.75463, 45.78096, 45.80708, 45.83298, 
    45.85866, 45.88413, 45.90938, 45.93441, 45.95922, 45.98381, 46.00818, 
    46.03233, 46.05627, 46.07998, 46.10347, 46.12674, 46.14979, 46.17262, 
    46.19522, 46.21761, 46.23976, 46.2617, 46.28341, 46.3049, 46.32616, 
    46.3472, 46.36802, 46.3886, 46.40897, 46.4291, 46.44901, 46.4687, 
    46.48815, 46.50738, 46.52638, 46.54516, 46.56371, 46.58202, 46.60011, 
    46.61797, 46.6356, 46.653, 46.67017, 46.68711, 46.70382, 46.7203, 
    46.73655, 46.75256, 46.76834, 46.7839, 46.79922, 46.81431, 46.82916, 
    46.84378, 46.85818, 46.87233, 46.88625, 46.89994, 46.9134, 46.92662, 
    46.93961, 46.95236, 46.96487, 46.97715, 46.9892, 47.00101, 47.01258, 
    47.02393, 47.03503, 47.04589, 47.05652, 47.06692, 47.07707, 47.08699, 
    47.09667, 47.10612, 47.11533, 47.12429, 47.13303, 47.14152, 47.14978, 
    47.15779, 47.16557, 47.17311, 47.18041, 47.18748, 47.1943, 47.20089, 
    47.20723, 47.21334, 47.2192, 47.22483, 47.23022, 47.23537, 47.24028, 
    47.24495, 47.24937, 47.25356, 47.25751, 47.26122, 47.26469, 47.26792, 
    47.2709, 47.27365, 47.27616, 47.27842, 47.28045, 47.28224, 47.28378, 
    47.28509, 47.28615, 47.28697, 47.28756, 47.2879, 47.288, 47.28786, 
    47.28748, 47.28686, 47.286, 47.2849, 47.28355, 47.28197, 47.28015, 
    47.27808, 47.27578, 47.27323, 47.27045, 47.26742, 47.26416, 47.26065, 
    47.2569, 47.25291, 47.24869, 47.24422, 47.23951, 47.23457, 47.22938, 
    47.22396, 47.21829, 47.21239, 47.20624, 47.19986, 47.19324, 47.18637, 
    47.17928, 47.17194, 47.16436, 47.15654, 47.14849, 47.14019, 47.13166, 
    47.12289, 47.11388, 47.10464, 47.09516, 47.08544, 47.07548, 47.06529, 
    47.05486, 47.04419, 47.03329, 47.02215, 47.01077, 46.99916, 46.98731, 
    46.97523, 46.96291, 46.95036, 46.93757, 46.92455, 46.91129, 46.89779, 
    46.88407, 46.87011, 46.85592, 46.84149, 46.82683, 46.81194, 46.79681, 
    46.78145, 46.76587, 46.75004, 46.73399, 46.7177, 46.70119, 46.68444, 
    46.66747, 46.65026, 46.63282, 46.61516, 46.59726, 46.57914, 46.56079, 
    46.5422, 46.52339, 46.50436, 46.48509, 46.4656, 46.44588, 46.42593, 
    46.40576, 46.38536, 46.36474, 46.34389, 46.32281, 46.30151, 46.27999, 
    46.25824, 46.23627, 46.21408, 46.19166, 46.16902, 46.14616, 46.12308, 
    46.09977, 46.07624, 46.0525, 46.02853, 46.00434, 45.97993, 45.95531, 
    45.93046, 45.9054, 45.88012, 45.85461, 45.8289, 45.80296, 45.77681, 
    45.75045, 45.72386, 45.69706, 45.67005, 45.64282, 45.61538, 45.58773, 
    45.55986, 45.53177, 45.50348, 45.47497, 45.44625, 45.41732, 45.38818, 
    45.35883, 45.32927, 45.2995, 45.26952, 45.23933, 45.20893, 45.17833, 
    45.14752, 45.1165, 45.08527, 45.05384, 45.02221, 44.99036, 44.95832, 
    44.92607, 44.89361, 44.86095, 44.82809, 44.79503, 44.76176, 44.72829, 
    44.69463, 44.66076, 44.62669, 44.59242, 44.55795, 44.52328, 44.48842, 
    44.45336, 44.4181, 44.38264, 44.34699, 44.31114, 44.27509, 44.23885, 
    44.20242, 44.16579, 44.12897, 44.09196, 44.05475, 44.01735, 43.97976, 
    43.94197, 43.904,
  39.71291, 39.76648, 39.81991, 39.8732, 39.92634, 39.97933, 40.03218, 
    40.08488, 40.13743, 40.18984, 40.2421, 40.2942, 40.34616, 40.39798, 
    40.44963, 40.50114, 40.5525, 40.60371, 40.65476, 40.70566, 40.75641, 
    40.807, 40.85744, 40.90773, 40.95786, 41.00784, 41.05765, 41.10732, 
    41.15682, 41.20617, 41.25535, 41.30438, 41.35325, 41.40196, 41.45051, 
    41.4989, 41.54713, 41.5952, 41.6431, 41.69085, 41.73842, 41.78584, 
    41.83309, 41.88017, 41.92709, 41.97385, 42.02044, 42.06686, 42.11311, 
    42.1592, 42.20512, 42.25087, 42.29645, 42.34186, 42.3871, 42.43217, 
    42.47707, 42.52179, 42.56635, 42.61073, 42.65493, 42.69897, 42.74282, 
    42.78651, 42.83002, 42.87335, 42.91651, 42.95948, 43.00229, 43.04491, 
    43.08736, 43.12962, 43.17171, 43.21362, 43.25534, 43.29689, 43.33825, 
    43.37944, 43.42044, 43.46125, 43.50189, 43.54234, 43.5826, 43.62268, 
    43.66257, 43.70229, 43.74181, 43.78114, 43.82029, 43.85925, 43.89802, 
    43.9366, 43.97499, 44.0132, 44.05121, 44.08904, 44.12666, 44.1641, 
    44.20135, 44.2384, 44.27526, 44.31193, 44.3484, 44.38468, 44.42076, 
    44.45665, 44.49234, 44.52783, 44.56313, 44.59822, 44.63312, 44.66782, 
    44.70233, 44.73663, 44.77073, 44.80463, 44.83834, 44.87184, 44.90513, 
    44.93823, 44.97112, 45.00381, 45.0363, 45.06858, 45.10066, 45.13253, 
    45.1642, 45.19566, 45.22691, 45.25796, 45.2888, 45.31943, 45.34985, 
    45.38007, 45.41008, 45.43987, 45.46946, 45.49884, 45.528, 45.55695, 
    45.5857, 45.61423, 45.64254, 45.67065, 45.69854, 45.72622, 45.75368, 
    45.78093, 45.80796, 45.83479, 45.86139, 45.88778, 45.91394, 45.9399, 
    45.96563, 45.99115, 46.01645, 46.04153, 46.06639, 46.09103, 46.11546, 
    46.13966, 46.16364, 46.1874, 46.21095, 46.23426, 46.25736, 46.28023, 
    46.30288, 46.32531, 46.34752, 46.3695, 46.39126, 46.41279, 46.4341, 
    46.45518, 46.47604, 46.49667, 46.51707, 46.53725, 46.55721, 46.57693, 
    46.59643, 46.6157, 46.63474, 46.65355, 46.67214, 46.69049, 46.70862, 
    46.72652, 46.74419, 46.76162, 46.77883, 46.79581, 46.81255, 46.82907, 
    46.84535, 46.8614, 46.87722, 46.8928, 46.90816, 46.92328, 46.93816, 
    46.95282, 46.96724, 46.98143, 46.99538, 47.0091, 47.02258, 47.03583, 
    47.04885, 47.06163, 47.07417, 47.08648, 47.09855, 47.11039, 47.12198, 
    47.13335, 47.14447, 47.15536, 47.16602, 47.17643, 47.18661, 47.19655, 
    47.20625, 47.21572, 47.22495, 47.23394, 47.24269, 47.2512, 47.25947, 
    47.26751, 47.2753, 47.28286, 47.29018, 47.29726, 47.30409, 47.31069, 
    47.31705, 47.32317, 47.32905, 47.33469, 47.34009, 47.34525, 47.35017, 
    47.35485, 47.35929, 47.36349, 47.36744, 47.37116, 47.37464, 47.37787, 
    47.38087, 47.38362, 47.38613, 47.3884, 47.39043, 47.39222, 47.39377, 
    47.39508, 47.39614, 47.39697, 47.39756, 47.3979, 47.398, 47.39786, 
    47.39748, 47.39686, 47.39599, 47.39489, 47.39354, 47.39196, 47.39013, 
    47.38806, 47.38575, 47.3832, 47.38041, 47.37738, 47.3741, 47.37059, 
    47.36683, 47.36284, 47.3586, 47.35413, 47.34941, 47.34445, 47.33925, 
    47.33382, 47.32814, 47.32222, 47.31606, 47.30967, 47.30303, 47.29615, 
    47.28904, 47.28168, 47.27409, 47.26625, 47.25818, 47.24987, 47.24132, 
    47.23253, 47.2235, 47.21424, 47.20473, 47.195, 47.18502, 47.1748, 
    47.16435, 47.15366, 47.14273, 47.13157, 47.12017, 47.10853, 47.09665, 
    47.08455, 47.0722, 47.05962, 47.0468, 47.03375, 47.02047, 47.00694, 
    46.99319, 46.9792, 46.96497, 46.95052, 46.93583, 46.9209, 46.90574, 
    46.89035, 46.87473, 46.85888, 46.84279, 46.82647, 46.80992, 46.79314, 
    46.77612, 46.75888, 46.74141, 46.72371, 46.70577, 46.68761, 46.66922, 
    46.65059, 46.63174, 46.61267, 46.59336, 46.57383, 46.55407, 46.53408, 
    46.51386, 46.49342, 46.47275, 46.45186, 46.43074, 46.4094, 46.38783, 
    46.36604, 46.34402, 46.32178, 46.29932, 46.27663, 46.25372, 46.23059, 
    46.20723, 46.18366, 46.15986, 46.13585, 46.11161, 46.08715, 46.06247, 
    46.03758, 46.01246, 45.98713, 45.96157, 45.93581, 45.90982, 45.88361, 
    45.85719, 45.83055, 45.8037, 45.77663, 45.74935, 45.72186, 45.69415, 
    45.66622, 45.63808, 45.60973, 45.58117, 45.55239, 45.5234, 45.4942, 
    45.46479, 45.43517, 45.40534, 45.37531, 45.34505, 45.3146, 45.28393, 
    45.25306, 45.22198, 45.19069, 45.1592, 45.1275, 45.0956, 45.06349, 
    45.03117, 44.99865, 44.96593, 44.93301, 44.89988, 44.86655, 44.83302, 
    44.79929, 44.76535, 44.73122, 44.69688, 44.66235, 44.62762, 44.59268, 
    44.55755, 44.52223, 44.4867, 44.45098, 44.41507, 44.37895, 44.34264, 
    44.30614, 44.26944, 44.23256, 44.19547, 44.15819, 44.12072, 44.08307, 
    44.04521, 44.00717,
  39.80887, 39.86252, 39.91603, 39.9694, 40.02262, 40.0757, 40.12862, 
    40.1814, 40.23404, 40.28653, 40.33886, 40.39105, 40.44309, 40.49498, 
    40.54672, 40.59831, 40.64975, 40.70103, 40.75217, 40.80315, 40.85398, 
    40.90466, 40.95517, 41.00554, 41.05575, 41.1058, 41.1557, 41.20544, 
    41.25503, 41.30445, 41.35372, 41.40283, 41.45178, 41.50057, 41.5492, 
    41.59767, 41.64598, 41.69412, 41.74211, 41.78993, 41.83759, 41.88508, 
    41.93241, 41.97957, 42.02657, 42.0734, 42.12007, 42.16657, 42.2129, 
    42.25907, 42.30506, 42.35089, 42.39655, 42.44204, 42.48735, 42.5325, 
    42.57747, 42.62228, 42.6669, 42.71136, 42.75565, 42.79976, 42.84369, 
    42.88745, 42.93104, 42.97445, 43.01768, 43.06073, 43.10361, 43.14631, 
    43.18883, 43.23117, 43.27333, 43.31532, 43.35712, 43.39874, 43.44017, 
    43.48143, 43.5225, 43.5634, 43.6041, 43.64463, 43.68496, 43.72512, 
    43.76508, 43.80486, 43.84446, 43.88387, 43.92308, 43.96212, 44.00096, 
    44.03961, 44.07808, 44.11635, 44.15443, 44.19233, 44.23003, 44.26754, 
    44.30485, 44.34197, 44.3789, 44.41564, 44.45218, 44.48853, 44.52467, 
    44.56063, 44.59639, 44.63195, 44.66731, 44.70248, 44.73744, 44.77221, 
    44.80678, 44.84115, 44.87532, 44.90928, 44.94305, 44.97662, 45.00998, 
    45.04314, 45.0761, 45.10885, 45.1414, 45.17374, 45.20588, 45.23782, 
    45.26955, 45.30107, 45.33238, 45.36349, 45.39439, 45.42509, 45.45557, 
    45.48584, 45.51591, 45.54576, 45.57541, 45.60485, 45.63407, 45.66308, 
    45.69188, 45.72047, 45.74884, 45.77701, 45.80495, 45.83269, 45.86021, 
    45.88751, 45.9146, 45.94147, 45.96813, 45.99457, 46.02079, 46.0468, 
    46.07259, 46.09816, 46.12351, 46.14864, 46.17356, 46.19825, 46.22272, 
    46.24697, 46.27101, 46.29482, 46.31841, 46.34177, 46.36492, 46.38784, 
    46.41054, 46.43301, 46.45527, 46.47729, 46.4991, 46.52067, 46.54203, 
    46.56315, 46.58405, 46.60473, 46.62518, 46.6454, 46.66539, 46.68516, 
    46.7047, 46.72401, 46.74309, 46.76194, 46.78057, 46.79897, 46.81713, 
    46.83506, 46.85277, 46.87024, 46.88749, 46.9045, 46.92128, 46.93783, 
    46.95415, 46.97023, 46.98608, 47.00171, 47.01709, 47.03225, 47.04716, 
    47.06185, 47.0763, 47.09052, 47.1045, 47.11825, 47.13176, 47.14504, 
    47.15808, 47.17089, 47.18346, 47.19579, 47.20789, 47.21975, 47.23138, 
    47.24277, 47.25392, 47.26483, 47.27551, 47.28595, 47.29615, 47.30611, 
    47.31583, 47.32532, 47.33457, 47.34357, 47.35234, 47.36088, 47.36917, 
    47.37722, 47.38503, 47.3926, 47.39994, 47.40703, 47.41389, 47.4205, 
    47.42688, 47.43301, 47.4389, 47.44455, 47.44996, 47.45514, 47.46006, 
    47.46476, 47.4692, 47.47341, 47.47738, 47.4811, 47.48458, 47.48783, 
    47.49083, 47.49359, 47.49611, 47.49838, 47.50042, 47.50221, 47.50377, 
    47.50507, 47.50614, 47.50697, 47.50755, 47.5079, 47.508, 47.50786, 
    47.50748, 47.50686, 47.50599, 47.50488, 47.50353, 47.50195, 47.50011, 
    47.49804, 47.49572, 47.49317, 47.49037, 47.48733, 47.48405, 47.48053, 
    47.47676, 47.47276, 47.46852, 47.46403, 47.4593, 47.45433, 47.44912, 
    47.44368, 47.43798, 47.43205, 47.42588, 47.41947, 47.41282, 47.40593, 
    47.3988, 47.39143, 47.38381, 47.37596, 47.36787, 47.35954, 47.35098, 
    47.34217, 47.33312, 47.32384, 47.31431, 47.30455, 47.29455, 47.28431, 
    47.27383, 47.26312, 47.25217, 47.24098, 47.22956, 47.2179, 47.20599, 
    47.19386, 47.18149, 47.16888, 47.15604, 47.14296, 47.12964, 47.11609, 
    47.10231, 47.08829, 47.07403, 47.05954, 47.04482, 47.02986, 47.01467, 
    46.99925, 46.98359, 46.9677, 46.95158, 46.93523, 46.91864, 46.90182, 
    46.88478, 46.8675, 46.84998, 46.83224, 46.81427, 46.79607, 46.77764, 
    46.75898, 46.74009, 46.72097, 46.70162, 46.68205, 46.66225, 46.64222, 
    46.62196, 46.60147, 46.58076, 46.55983, 46.53866, 46.51727, 46.49566, 
    46.47382, 46.45176, 46.42947, 46.40696, 46.38423, 46.36127, 46.33809, 
    46.31469, 46.29107, 46.26722, 46.24315, 46.21886, 46.19436, 46.16963, 
    46.14468, 46.11951, 46.09413, 46.06852, 46.0427, 46.01666, 45.9904, 
    45.96393, 45.93724, 45.91033, 45.88321, 45.85587, 45.82832, 45.80055, 
    45.77257, 45.74437, 45.71596, 45.68734, 45.65851, 45.62946, 45.6002, 
    45.57074, 45.54106, 45.51117, 45.48107, 45.45076, 45.42025, 45.38952, 
    45.35859, 45.32744, 45.2961, 45.26454, 45.23278, 45.20081, 45.16864, 
    45.13626, 45.10368, 45.0709, 45.03791, 45.00471, 44.97132, 44.93772, 
    44.90392, 44.86992, 44.83572, 44.80132, 44.76672, 44.73192, 44.69693, 
    44.66173, 44.62634, 44.59074, 44.55495, 44.51897, 44.48279, 44.44641, 
    44.40984, 44.37307, 44.33611, 44.29896, 44.26162, 44.22408, 44.18634, 
    44.14842, 44.11031,
  39.90479, 39.95852, 40.01211, 40.06556, 40.11886, 40.17202, 40.22503, 
    40.27789, 40.3306, 40.38317, 40.43559, 40.48786, 40.53998, 40.59195, 
    40.64377, 40.69544, 40.74696, 40.79832, 40.84954, 40.9006, 40.95151, 
    41.00227, 41.05286, 41.10331, 41.1536, 41.20374, 41.25371, 41.30354, 
    41.3532, 41.40271, 41.45205, 41.50124, 41.55027, 41.59914, 41.64785, 
    41.6964, 41.74479, 41.79301, 41.84107, 41.88897, 41.93671, 41.98428, 
    42.03169, 42.07893, 42.12601, 42.17292, 42.21967, 42.26625, 42.31266, 
    42.3589, 42.40497, 42.45088, 42.49661, 42.54218, 42.58757, 42.6328, 
    42.67785, 42.72273, 42.76744, 42.81197, 42.85633, 42.90052, 42.94453, 
    42.98837, 43.03203, 43.07551, 43.11882, 43.16195, 43.2049, 43.24768, 
    43.29027, 43.33269, 43.37493, 43.41698, 43.45886, 43.50055, 43.54207, 
    43.5834, 43.62455, 43.66551, 43.70629, 43.74689, 43.7873, 43.82752, 
    43.86756, 43.90742, 43.94708, 43.98656, 44.02586, 44.06496, 44.10387, 
    44.1426, 44.18113, 44.21948, 44.25763, 44.29559, 44.33337, 44.37094, 
    44.40833, 44.44552, 44.48252, 44.51933, 44.55593, 44.59235, 44.62857, 
    44.66459, 44.70042, 44.73604, 44.77147, 44.80671, 44.84174, 44.87658, 
    44.91121, 44.94564, 44.97988, 45.01391, 45.04774, 45.08138, 45.1148, 
    45.14803, 45.18105, 45.21386, 45.24648, 45.27888, 45.31109, 45.34309, 
    45.37488, 45.40646, 45.43784, 45.46901, 45.49997, 45.53072, 45.56127, 
    45.59161, 45.62173, 45.65165, 45.68135, 45.71085, 45.74013, 45.7692, 
    45.79805, 45.8267, 45.85513, 45.88335, 45.91135, 45.93914, 45.96672, 
    45.99408, 46.02122, 46.04815, 46.07486, 46.10136, 46.12763, 46.15369, 
    46.17953, 46.20515, 46.23056, 46.25574, 46.28071, 46.30545, 46.32998, 
    46.35428, 46.37836, 46.40222, 46.42586, 46.44927, 46.47247, 46.49543, 
    46.51818, 46.5407, 46.563, 46.58508, 46.60692, 46.62855, 46.64994, 
    46.67112, 46.69206, 46.71278, 46.73327, 46.75354, 46.77357, 46.79338, 
    46.81296, 46.83231, 46.85144, 46.87033, 46.88899, 46.90742, 46.92563, 
    46.9436, 46.96135, 46.97886, 46.99614, 47.01319, 47.03001, 47.04659, 
    47.06294, 47.07906, 47.09495, 47.1106, 47.12602, 47.1412, 47.15616, 
    47.17088, 47.18536, 47.19961, 47.21362, 47.2274, 47.24094, 47.25425, 
    47.26732, 47.28015, 47.29275, 47.30511, 47.31723, 47.32912, 47.34077, 
    47.35218, 47.36336, 47.3743, 47.385, 47.39546, 47.40568, 47.41566, 
    47.42541, 47.43492, 47.44419, 47.45321, 47.462, 47.47055, 47.47886, 
    47.48693, 47.49476, 47.50235, 47.5097, 47.51681, 47.52368, 47.53031, 
    47.5367, 47.54284, 47.54875, 47.55441, 47.55984, 47.56502, 47.56996, 
    47.57466, 47.57912, 47.58333, 47.58731, 47.59104, 47.59453, 47.59778, 
    47.60079, 47.60356, 47.60608, 47.60836, 47.6104, 47.6122, 47.61375, 
    47.61507, 47.61614, 47.61697, 47.61755, 47.6179, 47.618, 47.61786, 
    47.61748, 47.61685, 47.61599, 47.61488, 47.61353, 47.61193, 47.6101, 
    47.60802, 47.6057, 47.60313, 47.60033, 47.59729, 47.594, 47.59047, 
    47.5867, 47.58268, 47.57843, 47.57393, 47.56919, 47.56422, 47.55899, 
    47.55353, 47.54783, 47.54189, 47.5357, 47.52928, 47.52261, 47.5157, 
    47.50856, 47.50117, 47.49354, 47.48567, 47.47757, 47.46922, 47.46063, 
    47.4518, 47.44274, 47.43343, 47.42389, 47.4141, 47.40408, 47.39382, 
    47.38332, 47.37259, 47.36161, 47.3504, 47.33895, 47.32726, 47.31533, 
    47.30317, 47.29077, 47.27814, 47.26527, 47.25216, 47.23881, 47.22523, 
    47.21142, 47.19737, 47.18308, 47.16856, 47.15381, 47.13882, 47.1236, 
    47.10814, 47.09245, 47.07653, 47.06037, 47.04398, 47.02736, 47.01051, 
    46.99342, 46.9761, 46.95856, 46.94078, 46.92277, 46.90453, 46.88605, 
    46.86736, 46.84843, 46.82927, 46.80988, 46.79026, 46.77042, 46.75034, 
    46.73005, 46.70952, 46.68876, 46.66778, 46.64657, 46.62514, 46.60348, 
    46.5816, 46.55949, 46.53716, 46.5146, 46.49182, 46.46881, 46.44558, 
    46.42213, 46.39846, 46.37457, 46.35045, 46.32611, 46.30155, 46.27678, 
    46.25177, 46.22655, 46.20112, 46.17546, 46.14959, 46.12349, 46.09718, 
    46.07065, 46.04391, 46.01694, 45.98977, 45.96237, 45.93476, 45.90694, 
    45.8789, 45.85065, 45.82218, 45.7935, 45.76461, 45.73551, 45.70619, 
    45.67667, 45.64693, 45.61698, 45.58682, 45.55645, 45.52588, 45.49509, 
    45.46409, 45.43289, 45.40148, 45.36986, 45.33804, 45.30601, 45.27377, 
    45.24133, 45.20869, 45.17584, 45.14278, 45.10953, 45.07607, 45.04241, 
    45.00854, 44.97448, 44.94021, 44.90575, 44.87108, 44.83621, 44.80115, 
    44.76588, 44.73042, 44.69476, 44.65891, 44.62285, 44.5866, 44.55016, 
    44.51352, 44.47668, 44.43965, 44.40243, 44.36501, 44.3274, 44.2896, 
    44.25161, 44.21342,
  40.00066, 40.05448, 40.10815, 40.16168, 40.21506, 40.2683, 40.32138, 
    40.37433, 40.42712, 40.47977, 40.53227, 40.58463, 40.63683, 40.68888, 
    40.74078, 40.79253, 40.84413, 40.89558, 40.94687, 40.99801, 41.049, 
    41.09984, 41.15052, 41.20104, 41.25142, 41.30163, 41.35169, 41.40159, 
    41.45133, 41.50092, 41.55035, 41.59961, 41.64872, 41.69767, 41.74646, 
    41.79509, 41.84356, 41.89186, 41.94, 41.98798, 42.0358, 42.08345, 
    42.13094, 42.17826, 42.22541, 42.27241, 42.31923, 42.36589, 42.41238, 
    42.45869, 42.50485, 42.55083, 42.59665, 42.64229, 42.68776, 42.73306, 
    42.77819, 42.82315, 42.86794, 42.91254, 42.95698, 43.00125, 43.04533, 
    43.08925, 43.13298, 43.17654, 43.21993, 43.26314, 43.30616, 43.34901, 
    43.39169, 43.43418, 43.47649, 43.51862, 43.56057, 43.60234, 43.64393, 
    43.68534, 43.72656, 43.7676, 43.80845, 43.84912, 43.8896, 43.9299, 
    43.97002, 44.00994, 44.04968, 44.08923, 44.1286, 44.16777, 44.20676, 
    44.24556, 44.28416, 44.32258, 44.36081, 44.39884, 44.43668, 44.47433, 
    44.51178, 44.54905, 44.58612, 44.62299, 44.65967, 44.69615, 44.73244, 
    44.76853, 44.80442, 44.84012, 44.87562, 44.91092, 44.94602, 44.98092, 
    45.01562, 45.05012, 45.08442, 45.11852, 45.15242, 45.18612, 45.2196, 
    45.2529, 45.28598, 45.31886, 45.35154, 45.38401, 45.41628, 45.44834, 
    45.48019, 45.51184, 45.54328, 45.57451, 45.60553, 45.63634, 45.66695, 
    45.69735, 45.72754, 45.75751, 45.78727, 45.81683, 45.84617, 45.8753, 
    45.90421, 45.93291, 45.9614, 45.98968, 46.01774, 46.04559, 46.07322, 
    46.10063, 46.12783, 46.15482, 46.18158, 46.20813, 46.23446, 46.26057, 
    46.28646, 46.31214, 46.3376, 46.36283, 46.38785, 46.41264, 46.43722, 
    46.46157, 46.4857, 46.50961, 46.5333, 46.55676, 46.58001, 46.60302, 
    46.62582, 46.64838, 46.67073, 46.69285, 46.71474, 46.73641, 46.75785, 
    46.77907, 46.80006, 46.82082, 46.84136, 46.86166, 46.88174, 46.90159, 
    46.92122, 46.94061, 46.95977, 46.97871, 46.99741, 47.01588, 47.03413, 
    47.05214, 47.06992, 47.08747, 47.10479, 47.12187, 47.13872, 47.15534, 
    47.17173, 47.18789, 47.2038, 47.21949, 47.23494, 47.25016, 47.26515, 
    47.2799, 47.29441, 47.30869, 47.32273, 47.33654, 47.35011, 47.36345, 
    47.37655, 47.38941, 47.40203, 47.41442, 47.42657, 47.43849, 47.45016, 
    47.4616, 47.4728, 47.48376, 47.49448, 47.50497, 47.51521, 47.52522, 
    47.53499, 47.54451, 47.5538, 47.56285, 47.57166, 47.58023, 47.58855, 
    47.59664, 47.60449, 47.6121, 47.61946, 47.62659, 47.63347, 47.64011, 
    47.64651, 47.65268, 47.6586, 47.66427, 47.66971, 47.6749, 47.67986, 
    47.68456, 47.68903, 47.69326, 47.69724, 47.70098, 47.70448, 47.70774, 
    47.71075, 47.71352, 47.71605, 47.71834, 47.72038, 47.72219, 47.72374, 
    47.72506, 47.72614, 47.72696, 47.72755, 47.7279, 47.728, 47.72786, 
    47.72747, 47.72685, 47.72598, 47.72487, 47.72351, 47.72192, 47.72008, 
    47.71799, 47.71567, 47.7131, 47.71029, 47.70724, 47.70395, 47.70041, 
    47.69663, 47.6926, 47.68834, 47.68383, 47.67908, 47.6741, 47.66887, 
    47.66339, 47.65768, 47.65172, 47.64552, 47.63908, 47.6324, 47.62548, 
    47.61831, 47.61091, 47.60326, 47.59538, 47.58725, 47.57889, 47.57028, 
    47.56144, 47.55235, 47.54303, 47.53346, 47.52365, 47.51361, 47.50333, 
    47.49281, 47.48204, 47.47105, 47.45981, 47.44833, 47.43662, 47.42467, 
    47.41248, 47.40005, 47.38739, 47.37449, 47.36135, 47.34798, 47.33437, 
    47.32053, 47.30645, 47.29213, 47.27758, 47.26279, 47.24777, 47.23252, 
    47.21703, 47.2013, 47.18534, 47.16916, 47.15273, 47.13607, 47.11918, 
    47.10206, 47.08471, 47.06712, 47.0493, 47.03125, 47.01298, 46.99446, 
    46.97573, 46.95676, 46.93756, 46.91813, 46.89847, 46.87858, 46.85847, 
    46.83812, 46.81755, 46.79675, 46.77573, 46.75448, 46.733, 46.7113, 
    46.68937, 46.66721, 46.64483, 46.62223, 46.5994, 46.57634, 46.55307, 
    46.52957, 46.50584, 46.4819, 46.45773, 46.43335, 46.40874, 46.38391, 
    46.35886, 46.33358, 46.30809, 46.28239, 46.25646, 46.23031, 46.20395, 
    46.17736, 46.15056, 46.12354, 46.09631, 46.06886, 46.04119, 46.01332, 
    45.98522, 45.95691, 45.92839, 45.89965, 45.8707, 45.84154, 45.81216, 
    45.78258, 45.75278, 45.72277, 45.69255, 45.66212, 45.63148, 45.60064, 
    45.56958, 45.53832, 45.50684, 45.47517, 45.44328, 45.41119, 45.37889, 
    45.34638, 45.31367, 45.28076, 45.24764, 45.21432, 45.1808, 45.14707, 
    45.11314, 45.07901, 45.04468, 45.01014, 44.97541, 44.94048, 44.90535, 
    44.87001, 44.83448, 44.79876, 44.76283, 44.72671, 44.69039, 44.65388, 
    44.61717, 44.58027, 44.54317, 44.50587, 44.46839, 44.43071, 44.39283, 
    44.35477, 44.31652,
  40.09649, 40.15039, 40.20414, 40.25775, 40.31121, 40.36453, 40.41771, 
    40.47073, 40.52361, 40.57634, 40.62892, 40.68135, 40.73363, 40.78576, 
    40.83775, 40.88958, 40.94126, 40.99279, 41.04416, 41.09538, 41.14645, 
    41.19737, 41.24813, 41.29874, 41.34919, 41.39948, 41.44962, 41.4996, 
    41.54943, 41.59909, 41.6486, 41.69795, 41.74714, 41.79617, 41.84504, 
    41.89375, 41.94229, 41.99068, 42.0389, 42.08696, 42.13485, 42.18258, 
    42.23015, 42.27755, 42.32479, 42.37185, 42.41876, 42.46549, 42.51206, 
    42.55846, 42.60469, 42.65075, 42.69664, 42.74236, 42.78791, 42.83329, 
    42.8785, 42.92354, 42.9684, 43.01309, 43.0576, 43.10194, 43.14611, 
    43.1901, 43.23391, 43.27755, 43.32101, 43.36429, 43.4074, 43.45033, 
    43.49307, 43.53564, 43.57803, 43.62023, 43.66226, 43.7041, 43.74577, 
    43.78724, 43.82854, 43.86965, 43.91058, 43.95132, 43.99188, 44.03226, 
    44.07244, 44.11244, 44.15226, 44.19188, 44.23132, 44.27057, 44.30962, 
    44.34849, 44.38717, 44.42566, 44.46395, 44.50206, 44.53997, 44.57769, 
    44.61522, 44.65255, 44.68969, 44.72663, 44.76338, 44.79993, 44.83628, 
    44.87244, 44.90841, 44.94417, 44.97974, 45.01511, 45.05027, 45.08524, 
    45.12001, 45.15458, 45.18895, 45.22311, 45.25707, 45.29083, 45.32439, 
    45.35775, 45.3909, 45.42384, 45.45658, 45.48912, 45.52145, 45.55357, 
    45.58549, 45.6172, 45.6487, 45.67999, 45.71107, 45.74195, 45.77262, 
    45.80307, 45.83332, 45.86336, 45.89318, 45.92279, 45.95219, 45.98138, 
    46.01035, 46.03912, 46.06766, 46.09599, 46.12411, 46.15202, 46.1797, 
    46.20717, 46.23443, 46.26147, 46.28828, 46.31489, 46.34127, 46.36744, 
    46.39339, 46.41911, 46.44462, 46.46991, 46.49498, 46.51982, 46.54445, 
    46.56886, 46.59304, 46.61699, 46.64073, 46.66425, 46.68753, 46.7106, 
    46.73344, 46.75606, 46.77845, 46.80061, 46.82256, 46.84427, 46.86576, 
    46.88702, 46.90805, 46.92886, 46.94944, 46.96978, 46.98991, 47.0098, 
    47.02946, 47.0489, 47.0681, 47.08707, 47.10582, 47.12433, 47.14262, 
    47.16066, 47.17848, 47.19607, 47.21342, 47.23055, 47.24744, 47.26409, 
    47.28051, 47.2967, 47.31266, 47.32838, 47.34386, 47.35912, 47.37413, 
    47.38892, 47.40346, 47.41777, 47.43184, 47.44568, 47.45928, 47.47265, 
    47.48577, 47.49866, 47.51132, 47.52374, 47.53591, 47.54785, 47.55955, 
    47.57101, 47.58224, 47.59322, 47.60397, 47.61448, 47.62474, 47.63477, 
    47.64456, 47.65411, 47.66342, 47.67249, 47.68131, 47.6899, 47.69825, 
    47.70635, 47.71422, 47.72184, 47.72922, 47.73636, 47.74326, 47.74992, 
    47.75634, 47.76251, 47.76844, 47.77413, 47.77958, 47.78478, 47.78975, 
    47.79447, 47.79895, 47.80318, 47.80717, 47.81092, 47.81443, 47.81769, 
    47.82071, 47.82349, 47.82603, 47.82832, 47.83037, 47.83217, 47.83374, 
    47.83505, 47.83613, 47.83696, 47.83755, 47.8379, 47.838, 47.83786, 
    47.83747, 47.83685, 47.83598, 47.83486, 47.8335, 47.83191, 47.83006, 
    47.82797, 47.82564, 47.82307, 47.82025, 47.81719, 47.81389, 47.81034, 
    47.80656, 47.80253, 47.79825, 47.79374, 47.78898, 47.78398, 47.77873, 
    47.77325, 47.76752, 47.76155, 47.75534, 47.74888, 47.74219, 47.73525, 
    47.72807, 47.72065, 47.71299, 47.70509, 47.69695, 47.68856, 47.67994, 
    47.67107, 47.66196, 47.65261, 47.64303, 47.6332, 47.62314, 47.61283, 
    47.60229, 47.5915, 47.58048, 47.56922, 47.55772, 47.54598, 47.534, 
    47.52179, 47.50933, 47.49664, 47.48372, 47.47055, 47.45715, 47.44351, 
    47.42963, 47.41552, 47.40118, 47.38659, 47.37177, 47.35672, 47.34143, 
    47.32591, 47.31015, 47.29416, 47.27793, 47.26147, 47.24478, 47.22786, 
    47.2107, 47.1933, 47.17568, 47.15783, 47.13974, 47.12142, 47.10287, 
    47.08409, 47.06508, 47.04584, 47.02637, 47.00667, 46.98674, 46.96658, 
    46.94619, 46.92558, 46.90474, 46.88367, 46.86237, 46.84085, 46.8191, 
    46.79712, 46.77492, 46.75249, 46.72984, 46.70697, 46.68386, 46.66054, 
    46.63699, 46.61322, 46.58923, 46.56501, 46.54057, 46.51591, 46.49103, 
    46.46593, 46.4406, 46.41506, 46.3893, 46.36332, 46.33712, 46.3107, 
    46.28406, 46.2572, 46.23013, 46.20284, 46.17534, 46.14762, 46.11968, 
    46.09153, 46.06316, 46.03458, 46.00578, 45.97678, 45.94756, 45.91812, 
    45.88848, 45.85862, 45.82855, 45.79827, 45.76778, 45.73708, 45.70617, 
    45.67506, 45.64373, 45.61219, 45.58045, 45.5485, 45.51635, 45.48399, 
    45.45142, 45.41864, 45.38567, 45.35248, 45.3191, 45.28551, 45.25171, 
    45.21772, 45.18352, 45.14912, 45.11452, 45.07972, 45.04472, 45.00953, 
    44.97412, 44.93853, 44.90273, 44.86674, 44.83055, 44.79416, 44.75758, 
    44.7208, 44.68382, 44.64666, 44.60929, 44.57174, 44.53399, 44.49604, 
    44.45791, 44.41958,
  40.19228, 40.24626, 40.30009, 40.35379, 40.40733, 40.46073, 40.51398, 
    40.56709, 40.62004, 40.67286, 40.72552, 40.77803, 40.83039, 40.88261, 
    40.93467, 40.98658, 41.03835, 41.08995, 41.14141, 41.19271, 41.24387, 
    41.29486, 41.3457, 41.39639, 41.44692, 41.4973, 41.54752, 41.59758, 
    41.64748, 41.69723, 41.74682, 41.79625, 41.84552, 41.89463, 41.94358, 
    41.99236, 42.04099, 42.08945, 42.13776, 42.18589, 42.23387, 42.28168, 
    42.32933, 42.3768, 42.42412, 42.47127, 42.51825, 42.56506, 42.61171, 
    42.65819, 42.7045, 42.75064, 42.79661, 42.84241, 42.88803, 42.93349, 
    42.97878, 43.02389, 43.06883, 43.1136, 43.15819, 43.20261, 43.24685, 
    43.29092, 43.33481, 43.37852, 43.42206, 43.46542, 43.5086, 43.5516, 
    43.59443, 43.63707, 43.67953, 43.72181, 43.76392, 43.80584, 43.84757, 
    43.88913, 43.9305, 43.97168, 44.01269, 44.0535, 44.09414, 44.13458, 
    44.17484, 44.21492, 44.2548, 44.2945, 44.33401, 44.37333, 44.41246, 
    44.4514, 44.49015, 44.52871, 44.56708, 44.60525, 44.64323, 44.68103, 
    44.71862, 44.75602, 44.79323, 44.83025, 44.86706, 44.90369, 44.94011, 
    44.97634, 45.01237, 45.0482, 45.08384, 45.11927, 45.15451, 45.18954, 
    45.22438, 45.25901, 45.29345, 45.32768, 45.36171, 45.39553, 45.42916, 
    45.46257, 45.49579, 45.5288, 45.56161, 45.5942, 45.6266, 45.65878, 
    45.69077, 45.72254, 45.7541, 45.78546, 45.8166, 45.84754, 45.87827, 
    45.90878, 45.93909, 45.96918, 45.99907, 46.02874, 46.0582, 46.08745, 
    46.11648, 46.1453, 46.1739, 46.20229, 46.23047, 46.25843, 46.28617, 
    46.3137, 46.34101, 46.3681, 46.39498, 46.42163, 46.44807, 46.47429, 
    46.50029, 46.52608, 46.55164, 46.57698, 46.6021, 46.627, 46.65167, 
    46.67612, 46.70036, 46.72437, 46.74815, 46.77171, 46.79505, 46.81816, 
    46.84106, 46.86372, 46.88616, 46.90837, 46.93036, 46.95212, 46.97365, 
    46.99496, 47.01603, 47.03688, 47.05751, 47.0779, 47.09806, 47.118, 
    47.1377, 47.15718, 47.17643, 47.19544, 47.21422, 47.23278, 47.2511, 
    47.26919, 47.28704, 47.30467, 47.32206, 47.33922, 47.35614, 47.37284, 
    47.38929, 47.40552, 47.42151, 47.43726, 47.45278, 47.46807, 47.48312, 
    47.49793, 47.5125, 47.52685, 47.54095, 47.55482, 47.56845, 47.58184, 
    47.595, 47.60792, 47.6206, 47.63304, 47.64524, 47.65721, 47.66894, 
    47.68043, 47.69167, 47.70268, 47.71346, 47.72398, 47.73428, 47.74432, 
    47.75414, 47.7637, 47.77303, 47.78212, 47.79097, 47.79957, 47.80794, 
    47.81606, 47.82394, 47.83158, 47.83898, 47.84614, 47.85305, 47.85973, 
    47.86615, 47.87234, 47.87829, 47.88399, 47.88945, 47.89466, 47.89964, 
    47.90437, 47.90886, 47.9131, 47.9171, 47.92086, 47.92438, 47.92765, 
    47.93068, 47.93346, 47.936, 47.9383, 47.94035, 47.94216, 47.94373, 
    47.94505, 47.94613, 47.94696, 47.94755, 47.9479, 47.948, 47.94786, 
    47.94747, 47.94684, 47.94597, 47.94485, 47.94349, 47.94189, 47.94004, 
    47.93795, 47.93562, 47.93304, 47.93021, 47.92715, 47.92384, 47.92028, 
    47.91649, 47.91245, 47.90816, 47.90364, 47.89887, 47.89386, 47.8886, 
    47.8831, 47.87736, 47.87138, 47.86515, 47.85868, 47.85197, 47.84502, 
    47.83783, 47.83039, 47.82271, 47.81479, 47.80663, 47.79823, 47.78959, 
    47.7807, 47.77157, 47.76221, 47.7526, 47.74275, 47.73266, 47.72234, 
    47.71177, 47.70096, 47.68991, 47.67862, 47.6671, 47.65533, 47.64333, 
    47.63109, 47.61861, 47.60589, 47.59293, 47.57974, 47.56631, 47.55264, 
    47.53873, 47.52459, 47.51022, 47.4956, 47.48075, 47.46566, 47.45034, 
    47.43478, 47.41899, 47.40297, 47.38671, 47.37021, 47.35348, 47.33652, 
    47.31932, 47.3019, 47.28423, 47.26634, 47.24821, 47.22986, 47.21127, 
    47.19245, 47.1734, 47.15411, 47.1346, 47.11486, 47.09489, 47.07469, 
    47.05426, 47.0336, 47.01271, 46.9916, 46.97026, 46.94869, 46.9269, 
    46.90487, 46.88262, 46.86015, 46.83745, 46.81453, 46.79137, 46.768, 
    46.7444, 46.72058, 46.69654, 46.67227, 46.64778, 46.62307, 46.59814, 
    46.57298, 46.54761, 46.52201, 46.4962, 46.47016, 46.44391, 46.41743, 
    46.39074, 46.36383, 46.3367, 46.30936, 46.2818, 46.25402, 46.22603, 
    46.19782, 46.1694, 46.14075, 46.1119, 46.08284, 46.05355, 46.02406, 
    45.99436, 45.96444, 45.93431, 45.90397, 45.87342, 45.84266, 45.81169, 
    45.78051, 45.74912, 45.71753, 45.68572, 45.65371, 45.62149, 45.58906, 
    45.55643, 45.52359, 45.49055, 45.4573, 45.42385, 45.3902, 45.35634, 
    45.32228, 45.28801, 45.25355, 45.21888, 45.18401, 45.14895, 45.11368, 
    45.07821, 45.04255, 45.00668, 44.97062, 44.93436, 44.8979, 44.86125, 
    44.82441, 44.78736, 44.75012, 44.71269, 44.67506, 44.63724, 44.59922, 
    44.56102, 44.52262,
  40.28803, 40.34209, 40.396, 40.44978, 40.5034, 40.55688, 40.61022, 40.6634, 
    40.71644, 40.76934, 40.82208, 40.87467, 40.92712, 40.97941, 41.03156, 
    41.08355, 41.1354, 41.18708, 41.23862, 41.29, 41.34124, 41.39231, 
    41.44324, 41.49401, 41.54462, 41.59507, 41.64537, 41.69552, 41.7455, 
    41.79533, 41.845, 41.89451, 41.94386, 41.99305, 42.04208, 42.09095, 
    42.13965, 42.18819, 42.23658, 42.28479, 42.33285, 42.38074, 42.42847, 
    42.47602, 42.52342, 42.57065, 42.61771, 42.6646, 42.71133, 42.75788, 
    42.80427, 42.85049, 42.89654, 42.94242, 42.98812, 43.03366, 43.07902, 
    43.12421, 43.16923, 43.21407, 43.25874, 43.30324, 43.34756, 43.3917, 
    43.43567, 43.47946, 43.52308, 43.56651, 43.60977, 43.65285, 43.69575, 
    43.73847, 43.78101, 43.82336, 43.86554, 43.90754, 43.94935, 43.99098, 
    44.03242, 44.07368, 44.11476, 44.15565, 44.19636, 44.23688, 44.27721, 
    44.31736, 44.35732, 44.39709, 44.43667, 44.47607, 44.51527, 44.55428, 
    44.5931, 44.63173, 44.67017, 44.70842, 44.74648, 44.78434, 44.822, 
    44.85948, 44.89676, 44.93384, 44.97073, 45.00742, 45.04391, 45.08021, 
    45.11631, 45.15221, 45.18791, 45.22342, 45.25872, 45.29382, 45.32873, 
    45.36343, 45.39793, 45.43222, 45.46632, 45.50021, 45.5339, 45.56739, 
    45.60067, 45.63374, 45.66661, 45.69927, 45.73173, 45.76398, 45.79602, 
    45.82786, 45.85949, 45.8909, 45.92211, 45.95311, 45.9839, 46.01448, 
    46.04485, 46.075, 46.10495, 46.13468, 46.1642, 46.1935, 46.22259, 
    46.25147, 46.28013, 46.30858, 46.33681, 46.36483, 46.39263, 46.42021, 
    46.44758, 46.47473, 46.50166, 46.52837, 46.55486, 46.58114, 46.60719, 
    46.63303, 46.65864, 46.68403, 46.7092, 46.73415, 46.75888, 46.78339, 
    46.80767, 46.83173, 46.85556, 46.87917, 46.90256, 46.92572, 46.94866, 
    46.97137, 46.99386, 47.01612, 47.03815, 47.05996, 47.08154, 47.10289, 
    47.12401, 47.14491, 47.16557, 47.186, 47.20621, 47.22619, 47.24594, 
    47.26545, 47.28474, 47.30379, 47.32262, 47.34121, 47.35957, 47.3777, 
    47.3956, 47.41326, 47.43069, 47.44788, 47.46485, 47.48158, 47.49807, 
    47.51433, 47.53035, 47.54614, 47.5617, 47.57701, 47.59209, 47.60694, 
    47.62155, 47.63592, 47.65005, 47.66395, 47.67761, 47.69104, 47.70422, 
    47.71717, 47.72988, 47.74235, 47.75458, 47.76657, 47.77832, 47.78983, 
    47.80111, 47.81214, 47.82293, 47.83349, 47.8438, 47.85387, 47.8637, 
    47.87329, 47.88264, 47.89175, 47.90062, 47.90924, 47.91763, 47.92577, 
    47.93367, 47.94133, 47.94874, 47.95591, 47.96284, 47.96953, 47.97597, 
    47.98217, 47.98813, 47.99385, 47.99932, 48.00455, 48.00953, 48.01427, 
    48.01877, 48.02303, 48.02703, 48.0308, 48.03432, 48.0376, 48.04064, 
    48.04343, 48.04597, 48.04827, 48.05033, 48.05215, 48.05371, 48.05504, 
    48.05612, 48.05696, 48.05755, 48.0579, 48.058, 48.05786, 48.05747, 
    48.05684, 48.05597, 48.05485, 48.05349, 48.05188, 48.05003, 48.04793, 
    48.04559, 48.043, 48.04017, 48.0371, 48.03378, 48.03022, 48.02642, 
    48.02237, 48.01808, 48.01354, 48.00876, 48.00374, 47.99847, 47.99296, 
    47.98721, 47.98121, 47.97497, 47.96849, 47.96176, 47.95479, 47.94758, 
    47.94013, 47.93243, 47.9245, 47.91632, 47.90789, 47.89923, 47.89033, 
    47.88118, 47.8718, 47.86217, 47.85229, 47.84219, 47.83183, 47.82124, 
    47.81041, 47.79934, 47.78803, 47.77648, 47.76469, 47.75266, 47.74039, 
    47.72788, 47.71514, 47.70215, 47.68893, 47.67547, 47.66177, 47.64783, 
    47.63366, 47.61925, 47.60461, 47.58972, 47.5746, 47.55925, 47.54366, 
    47.52783, 47.51177, 47.49548, 47.47894, 47.46218, 47.44518, 47.42795, 
    47.41048, 47.39278, 47.37485, 47.35669, 47.33829, 47.31966, 47.3008, 
    47.28171, 47.26238, 47.24283, 47.22305, 47.20303, 47.18279, 47.16232, 
    47.14161, 47.12068, 47.09953, 47.07814, 47.05652, 47.03468, 47.01261, 
    46.99032, 46.9678, 46.94505, 46.92207, 46.89888, 46.87545, 46.85181, 
    46.82794, 46.80384, 46.77953, 46.75499, 46.73022, 46.70523, 46.68003, 
    46.6546, 46.62895, 46.60308, 46.577, 46.55069, 46.52416, 46.49741, 
    46.47045, 46.44326, 46.41586, 46.38824, 46.36041, 46.33236, 46.3041, 
    46.27561, 46.24692, 46.21801, 46.18888, 46.15954, 46.12999, 46.10022, 
    46.07024, 46.04005, 46.00965, 45.97904, 45.94822, 45.91719, 45.88595, 
    45.8545, 45.82284, 45.79097, 45.75889, 45.72661, 45.69412, 45.66142, 
    45.62852, 45.59542, 45.5621, 45.52859, 45.49487, 45.46094, 45.42682, 
    45.39248, 45.35795, 45.32322, 45.28828, 45.25315, 45.21781, 45.18228, 
    45.14655, 45.11061, 45.07448, 45.03815, 45.00163, 44.9649, 44.92799, 
    44.89087, 44.85356, 44.81606, 44.77836, 44.74047, 44.70238, 44.6641, 
    44.62564,
  40.38373, 40.43787, 40.49187, 40.54572, 40.59943, 40.65299, 40.70641, 
    40.75968, 40.8128, 40.86577, 40.9186, 40.97127, 41.0238, 41.07618, 
    41.1284, 41.18048, 41.2324, 41.28417, 41.33579, 41.38726, 41.43857, 
    41.48973, 41.54073, 41.59158, 41.64228, 41.69281, 41.74319, 41.79342, 
    41.84348, 41.89339, 41.94314, 41.99273, 42.04216, 42.09143, 42.14054, 
    42.18949, 42.23828, 42.2869, 42.33536, 42.38366, 42.43179, 42.47976, 
    42.52757, 42.57521, 42.62268, 42.66999, 42.71713, 42.7641, 42.81091, 
    42.85754, 42.90401, 42.95031, 42.99643, 43.04239, 43.08818, 43.13379, 
    43.17923, 43.2245, 43.2696, 43.31452, 43.35927, 43.40384, 43.44824, 
    43.49246, 43.5365, 43.58037, 43.62406, 43.66758, 43.71091, 43.75407, 
    43.79704, 43.83984, 43.88245, 43.92488, 43.96714, 44.00921, 44.05109, 
    44.0928, 44.13432, 44.17566, 44.21681, 44.25777, 44.29856, 44.33915, 
    44.37956, 44.41978, 44.45981, 44.49965, 44.53931, 44.57878, 44.61805, 
    44.65714, 44.69603, 44.73473, 44.77325, 44.81157, 44.84969, 44.88762, 
    44.92536, 44.96291, 45.00026, 45.03741, 45.07436, 45.11113, 45.14769, 
    45.18406, 45.22023, 45.2562, 45.29197, 45.32754, 45.36291, 45.39808, 
    45.43305, 45.46782, 45.50239, 45.53675, 45.57092, 45.60487, 45.63863, 
    45.67218, 45.70552, 45.73866, 45.7716, 45.80433, 45.83685, 45.86916, 
    45.90126, 45.93316, 45.96485, 45.99633, 46.0276, 46.05867, 46.08952, 
    46.12016, 46.15059, 46.1808, 46.2108, 46.2406, 46.27017, 46.29954, 
    46.32869, 46.35762, 46.38634, 46.41485, 46.44314, 46.47121, 46.49907, 
    46.52671, 46.55413, 46.58134, 46.60832, 46.63509, 46.66164, 46.68797, 
    46.71407, 46.73996, 46.76563, 46.79107, 46.8163, 46.8413, 46.86608, 
    46.89064, 46.91497, 46.93908, 46.96296, 46.98663, 47.01006, 47.03327, 
    47.05626, 47.07902, 47.10155, 47.12386, 47.14594, 47.16779, 47.18941, 
    47.21081, 47.23198, 47.25291, 47.27362, 47.29411, 47.31435, 47.33437, 
    47.35416, 47.37372, 47.39305, 47.41215, 47.43101, 47.44964, 47.46804, 
    47.48621, 47.50414, 47.52184, 47.53931, 47.55655, 47.57354, 47.59031, 
    47.60684, 47.62313, 47.63919, 47.65501, 47.6706, 47.68595, 47.70107, 
    47.71594, 47.73058, 47.74499, 47.75916, 47.77308, 47.78677, 47.80022, 
    47.81344, 47.82641, 47.83915, 47.85165, 47.86391, 47.87592, 47.8877, 
    47.89924, 47.91054, 47.9216, 47.93242, 47.94299, 47.95333, 47.96342, 
    47.97327, 47.98288, 47.99226, 48.00138, 48.01027, 48.01891, 48.02732, 
    48.03547, 48.04339, 48.05107, 48.0585, 48.06569, 48.07263, 48.07933, 
    48.08579, 48.09201, 48.09798, 48.1037, 48.10919, 48.11443, 48.11942, 
    48.12418, 48.12868, 48.13295, 48.13697, 48.14074, 48.14427, 48.14756, 
    48.1506, 48.1534, 48.15595, 48.15825, 48.16032, 48.16213, 48.16371, 
    48.16504, 48.16612, 48.16695, 48.16755, 48.1679, 48.168, 48.16786, 
    48.16747, 48.16684, 48.16596, 48.16484, 48.16348, 48.16186, 48.16001, 
    48.15791, 48.15556, 48.15297, 48.15014, 48.14705, 48.14373, 48.14016, 
    48.13635, 48.13229, 48.12799, 48.12344, 48.11865, 48.11362, 48.10834, 
    48.10281, 48.09705, 48.09104, 48.08479, 48.07829, 48.07155, 48.06456, 
    48.05734, 48.04987, 48.04216, 48.0342, 48.026, 48.01756, 48.00888, 
    47.99995, 47.99079, 47.98138, 47.97173, 47.96184, 47.95171, 47.94133, 
    47.93072, 47.91986, 47.90877, 47.89743, 47.88585, 47.87404, 47.86198, 
    47.84969, 47.83715, 47.82438, 47.81136, 47.79811, 47.78462, 47.7709, 
    47.75693, 47.74273, 47.72828, 47.71361, 47.69869, 47.68354, 47.66815, 
    47.65253, 47.63667, 47.62057, 47.60424, 47.58767, 47.57087, 47.55383, 
    47.53656, 47.51906, 47.50132, 47.48335, 47.46515, 47.44671, 47.42804, 
    47.40914, 47.39001, 47.37064, 47.35105, 47.33122, 47.31116, 47.29088, 
    47.27036, 47.24962, 47.22864, 47.20744, 47.186, 47.16434, 47.14246, 
    47.12034, 47.098, 47.07543, 47.05264, 47.02961, 47.00637, 46.98289, 
    46.9592, 46.93528, 46.91113, 46.88676, 46.86217, 46.83736, 46.81232, 
    46.78706, 46.76159, 46.73588, 46.70996, 46.68382, 46.65745, 46.63087, 
    46.60407, 46.57705, 46.54981, 46.52235, 46.49468, 46.46679, 46.43868, 
    46.41035, 46.38182, 46.35306, 46.32409, 46.29491, 46.26551, 46.2359, 
    46.20607, 46.17603, 46.14578, 46.11532, 46.08465, 46.05376, 46.02267, 
    45.99137, 45.95985, 45.92813, 45.8962, 45.86406, 45.83171, 45.79916, 
    45.7664, 45.73343, 45.70026, 45.66688, 45.6333, 45.59951, 45.56553, 
    45.53133, 45.49693, 45.46233, 45.42753, 45.39253, 45.35733, 45.32193, 
    45.28632, 45.25052, 45.21452, 45.17832, 45.14192, 45.10532, 45.06853, 
    45.03154, 44.99436, 44.95698, 44.91941, 44.88164, 44.84367, 44.80552, 
    44.76717, 44.72863,
  40.47939, 40.53362, 40.58769, 40.64163, 40.69542, 40.74906, 40.80256, 
    40.85591, 40.90911, 40.96217, 41.01507, 41.06783, 41.12044, 41.1729, 
    41.2252, 41.27736, 41.32936, 41.38122, 41.43292, 41.48447, 41.53586, 
    41.5871, 41.63819, 41.68912, 41.73989, 41.79051, 41.84097, 41.89128, 
    41.94143, 41.99141, 42.04124, 42.09092, 42.14043, 42.18978, 42.23897, 
    42.28799, 42.33686, 42.38557, 42.43411, 42.48249, 42.5307, 42.57875, 
    42.62664, 42.67435, 42.72191, 42.76929, 42.81652, 42.86357, 42.91045, 
    42.95717, 43.00372, 43.05009, 43.0963, 43.14233, 43.1882, 43.23389, 
    43.27941, 43.32476, 43.36993, 43.41493, 43.45975, 43.50441, 43.54888, 
    43.59318, 43.6373, 43.68125, 43.72502, 43.76861, 43.81202, 43.85525, 
    43.8983, 43.94117, 43.98387, 44.02637, 44.0687, 44.11085, 44.15281, 
    44.19459, 44.23619, 44.2776, 44.31883, 44.35987, 44.40072, 44.44139, 
    44.48187, 44.52217, 44.56227, 44.60219, 44.64192, 44.68146, 44.72081, 
    44.75997, 44.79893, 44.83771, 44.87629, 44.91468, 44.95288, 44.99089, 
    45.02869, 45.06631, 45.10373, 45.14095, 45.17798, 45.21481, 45.25145, 
    45.28788, 45.32412, 45.36016, 45.396, 45.43164, 45.46708, 45.50232, 
    45.53736, 45.57219, 45.60683, 45.64126, 45.67549, 45.70951, 45.74333, 
    45.77695, 45.81036, 45.84356, 45.87656, 45.90936, 45.94194, 45.97432, 
    46.00649, 46.03845, 46.0702, 46.10175, 46.13308, 46.1642, 46.19511, 
    46.22581, 46.25631, 46.28658, 46.31665, 46.3465, 46.37614, 46.40556, 
    46.43477, 46.46376, 46.49254, 46.52111, 46.54945, 46.57759, 46.6055, 
    46.6332, 46.66068, 46.68793, 46.71498, 46.7418, 46.7684, 46.79478, 
    46.82095, 46.84689, 46.87261, 46.89811, 46.92338, 46.94844, 46.97327, 
    46.99788, 47.02226, 47.04642, 47.07035, 47.09406, 47.11755, 47.14081, 
    47.16384, 47.18665, 47.20923, 47.23158, 47.25371, 47.27561, 47.29728, 
    47.31872, 47.33993, 47.36092, 47.38167, 47.40219, 47.42249, 47.44255, 
    47.46238, 47.48198, 47.50135, 47.52049, 47.53939, 47.55807, 47.57651, 
    47.59471, 47.61269, 47.63042, 47.64793, 47.6652, 47.68224, 47.69904, 
    47.7156, 47.73193, 47.74802, 47.76388, 47.7795, 47.79489, 47.81004, 
    47.82494, 47.83962, 47.85405, 47.86825, 47.88221, 47.89593, 47.90941, 
    47.92265, 47.93566, 47.94842, 47.96095, 47.97323, 47.98528, 47.99708, 
    48.00864, 48.01997, 48.03105, 48.04189, 48.05249, 48.06285, 48.07296, 
    48.08284, 48.09247, 48.10186, 48.11101, 48.11992, 48.12858, 48.137, 
    48.14518, 48.15311, 48.1608, 48.16825, 48.17546, 48.18242, 48.18913, 
    48.19561, 48.20184, 48.20782, 48.21356, 48.21906, 48.22431, 48.22932, 
    48.23408, 48.2386, 48.24287, 48.2469, 48.25068, 48.25422, 48.25751, 
    48.26056, 48.26336, 48.26592, 48.26823, 48.2703, 48.27212, 48.2737, 
    48.27503, 48.27611, 48.27695, 48.27755, 48.2779, 48.278, 48.27786, 
    48.27747, 48.27684, 48.27596, 48.27483, 48.27346, 48.27185, 48.26999, 
    48.26788, 48.26553, 48.26294, 48.26009, 48.25701, 48.25367, 48.2501, 
    48.24628, 48.24221, 48.2379, 48.23334, 48.22854, 48.2235, 48.2182, 
    48.21267, 48.20689, 48.20087, 48.1946, 48.18809, 48.18133, 48.17433, 
    48.16709, 48.1596, 48.15187, 48.1439, 48.13568, 48.12723, 48.11853, 
    48.10958, 48.1004, 48.09097, 48.0813, 48.07138, 48.06123, 48.05083, 
    48.04019, 48.02931, 48.01819, 48.00683, 47.99523, 47.98339, 47.9713, 
    47.95898, 47.94642, 47.93362, 47.92057, 47.9073, 47.89378, 47.88002, 
    47.86602, 47.85178, 47.83731, 47.8226, 47.80766, 47.79247, 47.77705, 
    47.76139, 47.74549, 47.72936, 47.713, 47.69639, 47.67955, 47.66248, 
    47.64518, 47.62763, 47.60986, 47.59185, 47.5736, 47.55513, 47.53642, 
    47.51748, 47.49831, 47.4789, 47.45926, 47.43939, 47.41929, 47.39896, 
    47.3784, 47.35761, 47.33659, 47.31535, 47.29387, 47.27216, 47.25023, 
    47.22807, 47.20567, 47.18306, 47.16021, 47.13715, 47.11385, 47.09033, 
    47.06658, 47.04261, 47.01842, 46.994, 46.96935, 46.94449, 46.9194, 
    46.89408, 46.86855, 46.8428, 46.81682, 46.79063, 46.76421, 46.73757, 
    46.71071, 46.68364, 46.65634, 46.62883, 46.6011, 46.57315, 46.54499, 
    46.5166, 46.48801, 46.45919, 46.43016, 46.40092, 46.37146, 46.34179, 
    46.3119, 46.28181, 46.2515, 46.22097, 46.19024, 46.15929, 46.12814, 
    46.09677, 46.06519, 46.03341, 46.00141, 45.96921, 45.9368, 45.90418, 
    45.87136, 45.83833, 45.80509, 45.77164, 45.738, 45.70414, 45.67009, 
    45.63583, 45.60136, 45.5667, 45.53183, 45.49676, 45.46149, 45.42601, 
    45.39034, 45.35447, 45.3184, 45.28213, 45.24566, 45.209, 45.17214, 
    45.13508, 45.09782, 45.06037, 45.02273, 44.98489, 44.94685, 44.90862, 
    44.8702, 44.83159,
  40.575, 40.62931, 40.68347, 40.73749, 40.79136, 40.84509, 40.89867, 
    40.9521, 41.00538, 41.05852, 41.11151, 41.16434, 41.21704, 41.26958, 
    41.32196, 41.3742, 41.42629, 41.47823, 41.53001, 41.58163, 41.63311, 
    41.68443, 41.7356, 41.78661, 41.83747, 41.88817, 41.93871, 41.9891, 
    42.03933, 42.08939, 42.13931, 42.18906, 42.23865, 42.28808, 42.33735, 
    42.38646, 42.43541, 42.4842, 42.53282, 42.58128, 42.62957, 42.6777, 
    42.72567, 42.77346, 42.8211, 42.86856, 42.91587, 42.963, 43.00996, 
    43.05676, 43.10338, 43.14984, 43.19613, 43.24224, 43.28818, 43.33395, 
    43.37955, 43.42498, 43.47023, 43.51531, 43.56021, 43.60494, 43.64949, 
    43.69387, 43.73807, 43.78209, 43.82594, 43.86961, 43.91309, 43.95641, 
    43.99953, 44.04248, 44.08525, 44.12783, 44.17024, 44.21246, 44.2545, 
    44.29636, 44.33803, 44.37952, 44.42082, 44.46193, 44.50286, 44.54361, 
    44.58416, 44.62453, 44.66471, 44.7047, 44.7445, 44.78412, 44.82354, 
    44.86277, 44.90181, 44.94066, 44.97931, 45.01778, 45.05605, 45.09412, 
    45.132, 45.16969, 45.20718, 45.24447, 45.28157, 45.31847, 45.35518, 
    45.39168, 45.42799, 45.4641, 45.50001, 45.53572, 45.57122, 45.60653, 
    45.64164, 45.67654, 45.71124, 45.74574, 45.78004, 45.81413, 45.84801, 
    45.8817, 45.91517, 45.94844, 45.98151, 46.01437, 46.04702, 46.07946, 
    46.11169, 46.14372, 46.17553, 46.20714, 46.23854, 46.26972, 46.30069, 
    46.33146, 46.36201, 46.39235, 46.42247, 46.45238, 46.48208, 46.51157, 
    46.54083, 46.56989, 46.59872, 46.62735, 46.65575, 46.68394, 46.71191, 
    46.73967, 46.7672, 46.79452, 46.82161, 46.84849, 46.87515, 46.90159, 
    46.9278, 46.9538, 46.97957, 47.00512, 47.03045, 47.05556, 47.08044, 
    47.1051, 47.12954, 47.15375, 47.17773, 47.20149, 47.22503, 47.24834, 
    47.27142, 47.29427, 47.3169, 47.3393, 47.36148, 47.38342, 47.40514, 
    47.42662, 47.44788, 47.46891, 47.48971, 47.51028, 47.53061, 47.55072, 
    47.57059, 47.59024, 47.60965, 47.62883, 47.64777, 47.66648, 47.68496, 
    47.70321, 47.72122, 47.739, 47.75654, 47.77385, 47.79092, 47.80776, 
    47.82436, 47.84072, 47.85685, 47.87275, 47.8884, 47.90382, 47.919, 
    47.93394, 47.94865, 47.96311, 47.97734, 47.99133, 48.00508, 48.01859, 
    48.03186, 48.0449, 48.05769, 48.07024, 48.08255, 48.09462, 48.10645, 
    48.11805, 48.12939, 48.1405, 48.15136, 48.16199, 48.17237, 48.18251, 
    48.19241, 48.20206, 48.21147, 48.22064, 48.22956, 48.23825, 48.24669, 
    48.25488, 48.26284, 48.27054, 48.27801, 48.28523, 48.2922, 48.29893, 
    48.30542, 48.31166, 48.31767, 48.32342, 48.32893, 48.33419, 48.33921, 
    48.34398, 48.34851, 48.35279, 48.35683, 48.36062, 48.36417, 48.36747, 
    48.37052, 48.37333, 48.37589, 48.37821, 48.38028, 48.38211, 48.38369, 
    48.38502, 48.38611, 48.38695, 48.38755, 48.3879, 48.388, 48.38786, 
    48.38747, 48.38683, 48.38595, 48.38483, 48.38345, 48.38184, 48.37997, 
    48.37786, 48.3755, 48.3729, 48.37005, 48.36696, 48.36362, 48.36003, 
    48.3562, 48.35213, 48.34781, 48.34324, 48.33843, 48.33337, 48.32807, 
    48.32252, 48.31673, 48.3107, 48.30441, 48.29789, 48.29111, 48.2841, 
    48.27684, 48.26934, 48.26159, 48.2536, 48.24537, 48.23689, 48.22817, 
    48.2192, 48.21, 48.20055, 48.19086, 48.18092, 48.17074, 48.16032, 
    48.14966, 48.13876, 48.12761, 48.11623, 48.1046, 48.09273, 48.08062, 
    48.06827, 48.05568, 48.04285, 48.02978, 48.01647, 48.00292, 47.98914, 
    47.97511, 47.96084, 47.94633, 47.93159, 47.91661, 47.90139, 47.88594, 
    47.87025, 47.85432, 47.83815, 47.82175, 47.80511, 47.78823, 47.77113, 
    47.75378, 47.7362, 47.71839, 47.70034, 47.68206, 47.66354, 47.64479, 
    47.62581, 47.60659, 47.58715, 47.56747, 47.54755, 47.52741, 47.50704, 
    47.48643, 47.4656, 47.44453, 47.42324, 47.40172, 47.37997, 47.35799, 
    47.33578, 47.31334, 47.29067, 47.26778, 47.24466, 47.22132, 47.19775, 
    47.17395, 47.14993, 47.12569, 47.10122, 47.07652, 47.0516, 47.02646, 
    47.0011, 46.97551, 46.9497, 46.92367, 46.89742, 46.87095, 46.84426, 
    46.81734, 46.79021, 46.76286, 46.73529, 46.7075, 46.6795, 46.65128, 
    46.62283, 46.59418, 46.56531, 46.53622, 46.50692, 46.4774, 46.44767, 
    46.41772, 46.38756, 46.35719, 46.32661, 46.29581, 46.2648, 46.23358, 
    46.20215, 46.17051, 46.13866, 46.10661, 46.07434, 46.04187, 46.00918, 
    45.97629, 45.9432, 45.90989, 45.87638, 45.84267, 45.80875, 45.77463, 
    45.7403, 45.70577, 45.67104, 45.6361, 45.60096, 45.56562, 45.53008, 
    45.49434, 45.4584, 45.42226, 45.38592, 45.34938, 45.31265, 45.27572, 
    45.23859, 45.20126, 45.16374, 45.12602, 45.08811, 45.05001, 45.01171, 
    44.97321, 44.93452,
  40.67057, 40.72496, 40.77921, 40.83331, 40.88726, 40.94107, 40.99473, 
    41.04824, 41.10161, 41.15483, 41.2079, 41.26082, 41.31359, 41.36621, 
    41.41868, 41.471, 41.52317, 41.57519, 41.62705, 41.67876, 41.73032, 
    41.78172, 41.83297, 41.88407, 41.93501, 41.98579, 42.03641, 42.08688, 
    42.13719, 42.18734, 42.23733, 42.28716, 42.33684, 42.38635, 42.4357, 
    42.48489, 42.53392, 42.58279, 42.63149, 42.68003, 42.7284, 42.77662, 
    42.82466, 42.87254, 42.92025, 42.9678, 43.01518, 43.06239, 43.10944, 
    43.15631, 43.20301, 43.24955, 43.29591, 43.34211, 43.38813, 43.43398, 
    43.47966, 43.52517, 43.5705, 43.61565, 43.66063, 43.70544, 43.75007, 
    43.79453, 43.83881, 43.88291, 43.92683, 43.97057, 44.01414, 44.05753, 
    44.10073, 44.14376, 44.1866, 44.22927, 44.27175, 44.31404, 44.35616, 
    44.39809, 44.43984, 44.4814, 44.52278, 44.56397, 44.60497, 44.64579, 
    44.68642, 44.72686, 44.76712, 44.80719, 44.84706, 44.88675, 44.92624, 
    44.96555, 45.00466, 45.04358, 45.08231, 45.12085, 45.15919, 45.19733, 
    45.23529, 45.27304, 45.3106, 45.34797, 45.38514, 45.42211, 45.45889, 
    45.49546, 45.53184, 45.56802, 45.60399, 45.63977, 45.67535, 45.71072, 
    45.7459, 45.78087, 45.81564, 45.8502, 45.88457, 45.91873, 45.95268, 
    45.98643, 46.01997, 46.05331, 46.08644, 46.11936, 46.15207, 46.18458, 
    46.21688, 46.24897, 46.28085, 46.31252, 46.34398, 46.37522, 46.40626, 
    46.43708, 46.4677, 46.4981, 46.52828, 46.55825, 46.58801, 46.61755, 
    46.64688, 46.676, 46.7049, 46.73357, 46.76204, 46.79028, 46.81831, 
    46.84612, 46.87371, 46.90109, 46.92824, 46.95517, 46.98189, 47.00838, 
    47.03465, 47.0607, 47.08652, 47.11213, 47.13751, 47.16267, 47.18761, 
    47.21231, 47.2368, 47.26106, 47.2851, 47.30891, 47.3325, 47.35585, 
    47.37899, 47.40189, 47.42456, 47.44701, 47.46923, 47.49123, 47.51299, 
    47.53452, 47.55582, 47.5769, 47.59774, 47.61835, 47.63873, 47.65888, 
    47.6788, 47.69848, 47.71794, 47.73716, 47.75614, 47.77489, 47.79342, 
    47.8117, 47.82975, 47.84756, 47.86515, 47.88249, 47.8996, 47.91647, 
    47.93311, 47.94951, 47.96568, 47.98161, 47.99729, 48.01274, 48.02796, 
    48.04293, 48.05767, 48.07217, 48.08643, 48.10045, 48.11423, 48.12777, 
    48.14107, 48.15413, 48.16695, 48.17953, 48.19187, 48.20397, 48.21583, 
    48.22744, 48.23882, 48.24995, 48.26084, 48.27148, 48.28189, 48.29205, 
    48.30197, 48.31165, 48.32108, 48.33027, 48.33921, 48.34791, 48.35637, 
    48.36459, 48.37255, 48.38028, 48.38776, 48.395, 48.40199, 48.40874, 
    48.41524, 48.42149, 48.42751, 48.43327, 48.43879, 48.44407, 48.4491, 
    48.45388, 48.45842, 48.46271, 48.46676, 48.47056, 48.47411, 48.47742, 
    48.48048, 48.4833, 48.48587, 48.48819, 48.49026, 48.4921, 48.49368, 
    48.49501, 48.49611, 48.49695, 48.49754, 48.49789, 48.498, 48.49786, 
    48.49747, 48.49683, 48.49595, 48.49482, 48.49344, 48.49182, 48.48995, 
    48.48784, 48.48548, 48.48287, 48.48001, 48.47691, 48.47356, 48.46997, 
    48.46613, 48.46205, 48.45772, 48.45314, 48.44832, 48.44325, 48.43793, 
    48.43238, 48.42657, 48.42052, 48.41423, 48.40768, 48.4009, 48.39387, 
    48.38659, 48.37907, 48.37131, 48.3633, 48.35505, 48.34655, 48.33781, 
    48.32883, 48.3196, 48.31013, 48.30042, 48.29046, 48.28026, 48.26981, 
    48.25913, 48.2482, 48.23703, 48.22562, 48.21397, 48.20207, 48.18994, 
    48.17756, 48.16494, 48.15208, 48.13898, 48.12564, 48.11207, 48.09825, 
    48.08419, 48.06989, 48.05536, 48.04058, 48.02557, 48.01031, 47.99483, 
    47.9791, 47.96313, 47.94693, 47.9305, 47.91382, 47.89691, 47.87976, 
    47.86238, 47.84476, 47.82691, 47.80882, 47.7905, 47.77195, 47.75315, 
    47.73413, 47.71487, 47.69538, 47.67566, 47.65571, 47.63552, 47.61511, 
    47.59446, 47.57358, 47.55247, 47.53113, 47.50956, 47.48776, 47.46573, 
    47.44348, 47.42099, 47.39828, 47.37534, 47.35217, 47.32878, 47.30516, 
    47.28131, 47.25724, 47.23294, 47.20842, 47.18368, 47.15871, 47.13351, 
    47.10809, 47.08245, 47.05659, 47.03051, 47.0042, 46.97768, 46.95093, 
    46.92396, 46.89677, 46.86937, 46.84174, 46.81389, 46.78583, 46.75755, 
    46.72905, 46.70034, 46.67141, 46.64226, 46.6129, 46.58332, 46.55353, 
    46.52352, 46.4933, 46.46287, 46.43222, 46.40136, 46.37029, 46.33901, 
    46.30752, 46.27582, 46.2439, 46.21178, 46.17945, 46.14691, 46.11416, 
    46.08121, 46.04805, 46.01468, 45.9811, 45.94732, 45.91334, 45.87915, 
    45.84475, 45.81015, 45.77535, 45.74035, 45.70514, 45.66973, 45.63412, 
    45.59832, 45.56231, 45.5261, 45.48969, 45.45308, 45.41628, 45.37927, 
    45.34207, 45.30468, 45.26708, 45.22929, 45.19131, 45.15313, 45.11476, 
    45.07619, 45.03744,
  40.7661, 40.82057, 40.8749, 40.92908, 40.98311, 41.037, 41.09075, 41.14434, 
    41.19779, 41.25109, 41.30424, 41.35725, 41.4101, 41.46281, 41.51536, 
    41.56776, 41.62001, 41.67211, 41.72406, 41.77585, 41.82749, 41.87897, 
    41.93031, 41.98148, 42.0325, 42.08336, 42.13407, 42.18462, 42.23501, 
    42.28524, 42.33532, 42.38523, 42.43498, 42.48458, 42.53401, 42.58328, 
    42.63239, 42.68134, 42.73012, 42.77874, 42.8272, 42.87549, 42.92361, 
    42.97158, 43.01937, 43.067, 43.11446, 43.16175, 43.20887, 43.25583, 
    43.30261, 43.34923, 43.39567, 43.44194, 43.48805, 43.53398, 43.57973, 
    43.62532, 43.67073, 43.71596, 43.76102, 43.80591, 43.85062, 43.89515, 
    43.93951, 43.98369, 44.02769, 44.07151, 44.11515, 44.15862, 44.2019, 
    44.245, 44.28793, 44.33067, 44.37322, 44.4156, 44.45779, 44.49979, 
    44.54162, 44.58326, 44.62471, 44.66597, 44.70705, 44.74795, 44.78865, 
    44.82917, 44.8695, 44.90964, 44.94959, 44.98935, 45.02892, 45.0683, 
    45.10748, 45.14648, 45.18528, 45.22388, 45.2623, 45.30052, 45.33854, 
    45.37637, 45.41401, 45.45144, 45.48868, 45.52573, 45.56257, 45.59922, 
    45.63566, 45.67191, 45.70796, 45.7438, 45.77945, 45.8149, 45.85014, 
    45.88518, 45.92001, 45.95465, 45.98908, 46.0233, 46.05732, 46.09114, 
    46.12474, 46.15815, 46.19134, 46.22433, 46.25711, 46.28968, 46.32204, 
    46.3542, 46.38614, 46.41787, 46.44939, 46.48071, 46.5118, 46.54269, 
    46.57336, 46.60382, 46.63408, 46.66411, 46.69392, 46.72353, 46.75292, 
    46.78209, 46.81105, 46.83979, 46.86831, 46.89661, 46.9247, 46.95256, 
    46.98021, 47.00764, 47.03485, 47.06184, 47.08861, 47.11516, 47.14148, 
    47.16758, 47.19347, 47.21912, 47.24456, 47.26977, 47.29476, 47.31952, 
    47.34406, 47.36837, 47.39246, 47.41632, 47.43995, 47.46336, 47.48654, 
    47.50949, 47.53222, 47.55471, 47.57698, 47.59902, 47.62083, 47.64241, 
    47.66376, 47.68488, 47.70576, 47.72642, 47.74684, 47.76704, 47.78699, 
    47.80672, 47.82622, 47.84548, 47.86451, 47.8833, 47.90186, 47.92018, 
    47.93827, 47.95613, 47.97375, 47.99113, 48.00828, 48.02518, 48.04186, 
    48.0583, 48.0745, 48.09046, 48.10618, 48.12167, 48.13691, 48.15192, 
    48.16669, 48.18122, 48.19551, 48.20956, 48.22338, 48.23695, 48.25028, 
    48.26337, 48.27621, 48.28882, 48.30119, 48.31331, 48.3252, 48.33684, 
    48.34824, 48.35939, 48.3703, 48.38098, 48.3914, 48.40159, 48.41153, 
    48.42123, 48.43068, 48.43989, 48.44886, 48.45758, 48.46605, 48.47429, 
    48.48227, 48.49002, 48.49751, 48.50476, 48.51177, 48.51854, 48.52505, 
    48.53132, 48.53735, 48.54313, 48.54866, 48.55395, 48.55899, 48.56378, 
    48.56833, 48.57263, 48.57669, 48.5805, 48.58406, 48.58737, 48.59044, 
    48.59327, 48.59584, 48.59817, 48.60025, 48.60208, 48.60367, 48.60501, 
    48.6061, 48.60695, 48.60754, 48.60789, 48.608, 48.60786, 48.60747, 
    48.60683, 48.60595, 48.60481, 48.60343, 48.60181, 48.59993, 48.59781, 
    48.59545, 48.59283, 48.58997, 48.58686, 48.58351, 48.57991, 48.57606, 
    48.57197, 48.56763, 48.56304, 48.5582, 48.55313, 48.5478, 48.54223, 
    48.53641, 48.53035, 48.52404, 48.51748, 48.51068, 48.50364, 48.49635, 
    48.48881, 48.48103, 48.473, 48.46473, 48.45621, 48.44745, 48.43845, 
    48.4292, 48.41971, 48.40997, 48.39999, 48.38977, 48.3793, 48.3686, 
    48.35764, 48.34645, 48.33501, 48.32333, 48.31141, 48.29925, 48.28685, 
    48.2742, 48.26131, 48.24818, 48.23482, 48.22121, 48.20736, 48.19327, 
    48.17894, 48.16437, 48.14956, 48.13452, 48.11923, 48.10371, 48.08795, 
    48.07195, 48.05571, 48.03924, 48.02253, 48.00558, 47.9884, 47.97097, 
    47.95332, 47.93543, 47.9173, 47.89894, 47.88034, 47.86151, 47.84245, 
    47.82315, 47.80362, 47.78385, 47.76385, 47.74363, 47.72317, 47.70247, 
    47.68155, 47.6604, 47.63901, 47.61739, 47.59555, 47.57347, 47.55117, 
    47.52864, 47.50588, 47.48289, 47.45967, 47.43623, 47.41256, 47.38866, 
    47.36454, 47.34019, 47.31562, 47.29082, 47.2658, 47.24055, 47.21508, 
    47.18939, 47.16347, 47.13733, 47.11097, 47.08439, 47.05759, 47.03056, 
    47.00332, 46.97586, 46.94817, 46.92027, 46.89215, 46.86381, 46.83525, 
    46.80648, 46.77749, 46.74828, 46.71886, 46.68922, 46.65937, 46.6293, 
    46.59902, 46.56853, 46.53782, 46.5069, 46.47577, 46.44442, 46.41287, 
    46.3811, 46.34912, 46.31694, 46.28454, 46.25194, 46.21913, 46.1861, 
    46.15288, 46.11944, 46.0858, 46.05196, 46.0179, 45.98365, 45.94918, 
    45.91452, 45.87965, 45.84458, 45.8093, 45.77383, 45.73815, 45.70227, 
    45.66619, 45.62991, 45.59343, 45.55676, 45.51988, 45.4828, 45.44553, 
    45.40807, 45.3704, 45.33254, 45.29449, 45.25624, 45.21779, 45.17915, 
    45.14032,
  40.86158, 40.91613, 40.97054, 41.02481, 41.07893, 41.1329, 41.18672, 
    41.2404, 41.29393, 41.34732, 41.40055, 41.45364, 41.50657, 41.55936, 
    41.612, 41.66448, 41.71681, 41.76899, 41.82102, 41.87289, 41.92462, 
    41.97618, 42.0276, 42.07885, 42.12996, 42.1809, 42.23169, 42.28232, 
    42.33279, 42.38311, 42.43326, 42.48326, 42.53309, 42.58277, 42.63228, 
    42.68163, 42.73082, 42.77985, 42.82872, 42.87742, 42.92596, 42.97433, 
    43.02253, 43.07058, 43.11845, 43.16616, 43.2137, 43.26107, 43.30827, 
    43.35531, 43.40217, 43.44887, 43.49539, 43.54174, 43.58793, 43.63394, 
    43.67977, 43.72544, 43.77092, 43.81624, 43.86138, 43.90634, 43.95113, 
    43.99574, 44.04018, 44.08443, 44.12851, 44.17241, 44.21613, 44.25967, 
    44.30304, 44.34622, 44.38921, 44.43203, 44.47467, 44.51712, 44.55938, 
    44.60147, 44.64337, 44.68508, 44.72661, 44.76795, 44.80911, 44.85007, 
    44.89086, 44.93145, 44.97185, 45.01207, 45.05209, 45.09193, 45.13157, 
    45.17102, 45.21028, 45.24935, 45.28822, 45.3269, 45.36539, 45.40368, 
    45.44178, 45.47968, 45.51738, 45.55489, 45.5922, 45.62931, 45.66623, 
    45.70295, 45.73946, 45.77578, 45.8119, 45.84781, 45.88353, 45.91904, 
    45.95435, 45.98946, 46.02437, 46.05907, 46.09357, 46.12786, 46.16195, 
    46.19583, 46.2295, 46.26297, 46.29623, 46.32928, 46.36213, 46.39476, 
    46.42719, 46.45941, 46.49142, 46.52321, 46.5548, 46.58617, 46.61733, 
    46.64828, 46.67902, 46.70954, 46.73985, 46.76994, 46.79982, 46.82949, 
    46.85894, 46.88817, 46.91718, 46.94598, 46.97456, 47.00292, 47.03107, 
    47.05899, 47.0867, 47.11419, 47.14145, 47.1685, 47.19532, 47.22192, 
    47.2483, 47.27446, 47.3004, 47.32611, 47.35159, 47.37686, 47.4019, 
    47.42671, 47.4513, 47.47567, 47.49981, 47.52372, 47.5474, 47.57086, 
    47.59409, 47.61709, 47.63986, 47.6624, 47.68472, 47.70681, 47.72866, 
    47.75029, 47.77168, 47.79284, 47.81378, 47.83448, 47.85495, 47.87518, 
    47.89518, 47.91496, 47.93449, 47.95379, 47.97286, 47.9917, 48.0103, 
    48.02866, 48.04679, 48.06468, 48.08234, 48.09976, 48.11695, 48.13389, 
    48.1506, 48.16708, 48.18331, 48.19931, 48.21507, 48.23058, 48.24586, 
    48.26091, 48.27571, 48.29027, 48.30459, 48.31868, 48.33252, 48.34612, 
    48.35948, 48.3726, 48.38548, 48.39811, 48.4105, 48.42265, 48.43456, 
    48.44623, 48.45765, 48.46883, 48.47977, 48.49047, 48.50092, 48.51112, 
    48.52109, 48.53081, 48.54028, 48.54951, 48.5585, 48.56724, 48.57573, 
    48.58398, 48.59199, 48.59975, 48.60727, 48.61453, 48.62156, 48.62833, 
    48.63486, 48.64115, 48.64719, 48.65298, 48.65853, 48.66383, 48.66888, 
    48.67368, 48.67824, 48.68255, 48.68661, 48.69043, 48.694, 48.69733, 
    48.7004, 48.70323, 48.70581, 48.70815, 48.71023, 48.71207, 48.71366, 
    48.715, 48.71609, 48.71694, 48.71754, 48.7179, 48.718, 48.71786, 
    48.71746, 48.71683, 48.71594, 48.71481, 48.71342, 48.71179, 48.70992, 
    48.70779, 48.70542, 48.7028, 48.69993, 48.69682, 48.69345, 48.68985, 
    48.68599, 48.68189, 48.67754, 48.67294, 48.66809, 48.663, 48.65767, 
    48.65208, 48.64625, 48.64017, 48.63385, 48.62728, 48.62046, 48.6134, 
    48.60609, 48.59854, 48.59074, 48.5827, 48.57441, 48.56587, 48.55709, 
    48.54807, 48.5388, 48.52929, 48.51953, 48.50953, 48.49928, 48.48879, 
    48.47806, 48.46708, 48.45586, 48.4444, 48.4327, 48.42075, 48.40856, 
    48.39613, 48.38345, 48.37054, 48.35738, 48.34398, 48.33035, 48.31646, 
    48.30235, 48.28798, 48.27338, 48.25854, 48.24347, 48.22815, 48.21259, 
    48.19679, 48.18076, 48.16449, 48.14798, 48.13123, 48.11424, 48.09702, 
    48.07956, 48.06187, 48.04394, 48.02577, 48.00737, 47.98873, 47.96986, 
    47.95076, 47.93142, 47.91184, 47.89204, 47.87199, 47.85172, 47.83122, 
    47.81048, 47.78951, 47.76831, 47.74688, 47.72522, 47.70333, 47.68121, 
    47.65886, 47.63627, 47.61346, 47.59043, 47.56716, 47.54367, 47.51995, 
    47.496, 47.47183, 47.44743, 47.4228, 47.39795, 47.37288, 47.34758, 
    47.32206, 47.29631, 47.27034, 47.24414, 47.21773, 47.19109, 47.16423, 
    47.13715, 47.10985, 47.08233, 47.05459, 47.02663, 46.99845, 46.97005, 
    46.94144, 46.91261, 46.88356, 46.85429, 46.82481, 46.79511, 46.7652, 
    46.73507, 46.70473, 46.67417, 46.6434, 46.61242, 46.58122, 46.54982, 
    46.5182, 46.48637, 46.45433, 46.42208, 46.38961, 46.35695, 46.32407, 
    46.29098, 46.25769, 46.22419, 46.19048, 46.15657, 46.12245, 46.08812, 
    46.05359, 46.01886, 45.98392, 45.94878, 45.91344, 45.87789, 45.84215, 
    45.8062, 45.77005, 45.7337, 45.69715, 45.6604, 45.62346, 45.58631, 
    45.54897, 45.51143, 45.47369, 45.43576, 45.39764, 45.35931, 45.32079, 
    45.28209, 45.24318,
  40.95702, 41.01165, 41.06614, 41.12049, 41.17469, 41.22874, 41.28265, 
    41.33641, 41.39003, 41.44349, 41.49681, 41.54998, 41.603, 41.65587, 
    41.70858, 41.76115, 41.81357, 41.86583, 41.91794, 41.9699, 42.0217, 
    42.07335, 42.12484, 42.17618, 42.22737, 42.27839, 42.32927, 42.37998, 
    42.43053, 42.48093, 42.53117, 42.58124, 42.63116, 42.68092, 42.73051, 
    42.77995, 42.82922, 42.87833, 42.92727, 42.97606, 43.02467, 43.07313, 
    43.12141, 43.16954, 43.21749, 43.26528, 43.3129, 43.36036, 43.40764, 
    43.45475, 43.5017, 43.54847, 43.59508, 43.64151, 43.68777, 43.73386, 
    43.77978, 43.82552, 43.87109, 43.91648, 43.9617, 44.00674, 44.05161, 
    44.0963, 44.14082, 44.18515, 44.22931, 44.27328, 44.31708, 44.3607, 
    44.40414, 44.4474, 44.49047, 44.53337, 44.57608, 44.61861, 44.66095, 
    44.70311, 44.74509, 44.78688, 44.82848, 44.8699, 44.91113, 44.95218, 
    44.99303, 45.0337, 45.07418, 45.11447, 45.15456, 45.19447, 45.23419, 
    45.27372, 45.31305, 45.35219, 45.39114, 45.42989, 45.46845, 45.50681, 
    45.54498, 45.58295, 45.62073, 45.65831, 45.69569, 45.73288, 45.76987, 
    45.80665, 45.84324, 45.87963, 45.91581, 45.9518, 45.98759, 46.02317, 
    46.05855, 46.09372, 46.1287, 46.16347, 46.19803, 46.23239, 46.26654, 
    46.3005, 46.33424, 46.36777, 46.4011, 46.43422, 46.46712, 46.49983, 
    46.53232, 46.5646, 46.59667, 46.62853, 46.66018, 46.69162, 46.72284, 
    46.75386, 46.78465, 46.81524, 46.84561, 46.87576, 46.9057, 46.93543, 
    46.96494, 46.99423, 47.0233, 47.05216, 47.0808, 47.10922, 47.13742, 
    47.16541, 47.19317, 47.22071, 47.24804, 47.27514, 47.30201, 47.32867, 
    47.35511, 47.38132, 47.40731, 47.43307, 47.45862, 47.48394, 47.50903, 
    47.53389, 47.55854, 47.58295, 47.60714, 47.6311, 47.65483, 47.67834, 
    47.70162, 47.72467, 47.74749, 47.77008, 47.79245, 47.81458, 47.83648, 
    47.85815, 47.8796, 47.90081, 47.92178, 47.94253, 47.96304, 47.98332, 
    48.00336, 48.02318, 48.04276, 48.0621, 48.08121, 48.10009, 48.11873, 
    48.13713, 48.1553, 48.17323, 48.19093, 48.20839, 48.22561, 48.24259, 
    48.25934, 48.27585, 48.29212, 48.30815, 48.32394, 48.3395, 48.35481, 
    48.36989, 48.38472, 48.39931, 48.41367, 48.42778, 48.44165, 48.45529, 
    48.46868, 48.48182, 48.49473, 48.50739, 48.51981, 48.53199, 48.54393, 
    48.55562, 48.56707, 48.57828, 48.58924, 48.59996, 48.61043, 48.62066, 
    48.63065, 48.64039, 48.64988, 48.65913, 48.66814, 48.6769, 48.68541, 
    48.69368, 48.70171, 48.70948, 48.71701, 48.7243, 48.73134, 48.73813, 
    48.74468, 48.75098, 48.75703, 48.76283, 48.76839, 48.7737, 48.77877, 
    48.78358, 48.78815, 48.79247, 48.79655, 48.80037, 48.80395, 48.80728, 
    48.81036, 48.8132, 48.81578, 48.81812, 48.82021, 48.82206, 48.82365, 
    48.82499, 48.82609, 48.82694, 48.82754, 48.8279, 48.828, 48.82785, 
    48.82747, 48.82682, 48.82594, 48.8248, 48.82341, 48.82178, 48.8199, 
    48.81777, 48.81539, 48.81277, 48.80989, 48.80677, 48.8034, 48.79978, 
    48.79592, 48.79181, 48.78745, 48.78284, 48.77798, 48.77288, 48.76753, 
    48.76193, 48.75609, 48.75, 48.74366, 48.73708, 48.73024, 48.72316, 
    48.71584, 48.70827, 48.70045, 48.69239, 48.68408, 48.67553, 48.66673, 
    48.65769, 48.6484, 48.63886, 48.62908, 48.61906, 48.60879, 48.59828, 
    48.58752, 48.57652, 48.56528, 48.55379, 48.54206, 48.53008, 48.51786, 
    48.50541, 48.4927, 48.47976, 48.46658, 48.45315, 48.43948, 48.42557, 
    48.41142, 48.39702, 48.38239, 48.36752, 48.35241, 48.33705, 48.32146, 
    48.30563, 48.28956, 48.27325, 48.25671, 48.23992, 48.2229, 48.20564, 
    48.18814, 48.17041, 48.15244, 48.13424, 48.1158, 48.09712, 48.07821, 
    48.05906, 48.03968, 48.02006, 48.00021, 47.98013, 47.95981, 47.93926, 
    47.91848, 47.89746, 47.87622, 47.85474, 47.83303, 47.8111, 47.78893, 
    47.76653, 47.7439, 47.72104, 47.69796, 47.67464, 47.6511, 47.62733, 
    47.60333, 47.57911, 47.55465, 47.52998, 47.50507, 47.47995, 47.45459, 
    47.42902, 47.40321, 47.37719, 47.35094, 47.32447, 47.29778, 47.27086, 
    47.24373, 47.21637, 47.18879, 47.161, 47.13298, 47.10474, 47.07629, 
    47.04761, 47.01872, 46.98961, 46.96029, 46.93074, 46.90098, 46.87101, 
    46.84082, 46.81041, 46.7798, 46.74896, 46.71792, 46.68666, 46.65519, 
    46.62351, 46.59161, 46.55951, 46.52719, 46.49467, 46.46193, 46.42899, 
    46.39584, 46.36248, 46.32891, 46.29514, 46.26116, 46.22697, 46.19258, 
    46.15798, 46.12318, 46.08817, 46.05296, 46.01755, 45.98194, 45.94612, 
    45.9101, 45.87389, 45.83747, 45.80085, 45.76403, 45.72701, 45.68979, 
    45.65238, 45.61477, 45.57696, 45.53896, 45.50076, 45.46236, 45.42377, 
    45.38499, 45.34601,
  41.05241, 41.10713, 41.1617, 41.21613, 41.27041, 41.32455, 41.37854, 
    41.43238, 41.48608, 41.53963, 41.59303, 41.64628, 41.69938, 41.75233, 
    41.80513, 41.85778, 41.91028, 41.96262, 42.01482, 42.06686, 42.11874, 
    42.17048, 42.22205, 42.27347, 42.32474, 42.37585, 42.4268, 42.4776, 
    42.52823, 42.57871, 42.62903, 42.67919, 42.72919, 42.77903, 42.8287, 
    42.87822, 42.92757, 42.97676, 43.02579, 43.07466, 43.12336, 43.17189, 
    43.22026, 43.26846, 43.3165, 43.36437, 43.41207, 43.4596, 43.50697, 
    43.55416, 43.60119, 43.64804, 43.69473, 43.74124, 43.78758, 43.83375, 
    43.87975, 43.92557, 43.97121, 44.01669, 44.06199, 44.10711, 44.15205, 
    44.19682, 44.24142, 44.28583, 44.33007, 44.37412, 44.418, 44.4617, 
    44.50521, 44.54855, 44.5917, 44.63467, 44.67746, 44.72007, 44.76249, 
    44.80473, 44.84678, 44.88865, 44.93032, 44.97182, 45.01313, 45.05424, 
    45.09518, 45.13592, 45.17647, 45.21684, 45.25701, 45.29699, 45.33678, 
    45.37638, 45.41579, 45.45501, 45.49403, 45.53285, 45.57148, 45.60992, 
    45.64816, 45.68621, 45.72406, 45.76171, 45.79916, 45.83642, 45.87348, 
    45.91034, 45.94699, 45.98345, 46.01971, 46.05576, 46.09162, 46.12727, 
    46.16272, 46.19796, 46.23301, 46.26785, 46.30248, 46.33691, 46.37112, 
    46.40514, 46.43895, 46.47255, 46.50594, 46.53913, 46.57211, 46.60487, 
    46.63743, 46.66977, 46.70191, 46.73383, 46.76555, 46.79705, 46.82833, 
    46.85941, 46.89027, 46.92092, 46.95135, 46.98157, 47.01157, 47.04136, 
    47.07092, 47.10027, 47.12941, 47.15833, 47.18702, 47.2155, 47.24376, 
    47.2718, 47.29963, 47.32722, 47.3546, 47.38176, 47.4087, 47.43541, 
    47.4619, 47.48817, 47.51421, 47.54003, 47.56563, 47.591, 47.61614, 
    47.64106, 47.66576, 47.69022, 47.71446, 47.73848, 47.76226, 47.78582, 
    47.80915, 47.83224, 47.85512, 47.87776, 47.90017, 47.92235, 47.9443, 
    47.96601, 47.9875, 48.00876, 48.02978, 48.05057, 48.07113, 48.09145, 
    48.11154, 48.13139, 48.15102, 48.1704, 48.18956, 48.20847, 48.22715, 
    48.24559, 48.26381, 48.28178, 48.29951, 48.31701, 48.33427, 48.35129, 
    48.36807, 48.38462, 48.40092, 48.41699, 48.43282, 48.44841, 48.46375, 
    48.47886, 48.49373, 48.50836, 48.52274, 48.53689, 48.55079, 48.56445, 
    48.57787, 48.59105, 48.60398, 48.61667, 48.62912, 48.64133, 48.65329, 
    48.66501, 48.67648, 48.68771, 48.6987, 48.70944, 48.71994, 48.73019, 
    48.7402, 48.74997, 48.75948, 48.76875, 48.77778, 48.78656, 48.79509, 
    48.80338, 48.81142, 48.81922, 48.82677, 48.83407, 48.84112, 48.84793, 
    48.85449, 48.8608, 48.86687, 48.87269, 48.87826, 48.88358, 48.88866, 
    48.89348, 48.89806, 48.90239, 48.90648, 48.91031, 48.91389, 48.91723, 
    48.92032, 48.92316, 48.92575, 48.9281, 48.93019, 48.93204, 48.93364, 
    48.93499, 48.93609, 48.93694, 48.93754, 48.93789, 48.938, 48.93785, 
    48.93746, 48.93682, 48.93593, 48.93479, 48.9334, 48.93177, 48.92988, 
    48.92775, 48.92536, 48.92273, 48.91985, 48.91672, 48.91335, 48.90972, 
    48.90585, 48.90172, 48.89735, 48.89273, 48.88787, 48.88276, 48.87739, 
    48.87178, 48.86592, 48.85982, 48.85347, 48.84687, 48.84002, 48.83293, 
    48.82559, 48.818, 48.81017, 48.80209, 48.79376, 48.78519, 48.77637, 
    48.7673, 48.75799, 48.74844, 48.73864, 48.72859, 48.7183, 48.70776, 
    48.69698, 48.68596, 48.67469, 48.66317, 48.65141, 48.63941, 48.62717, 
    48.61468, 48.60195, 48.58898, 48.57576, 48.56231, 48.54861, 48.53466, 
    48.52048, 48.50606, 48.49139, 48.47649, 48.46134, 48.44596, 48.43033, 
    48.41446, 48.39836, 48.38202, 48.36543, 48.34861, 48.33155, 48.31425, 
    48.29672, 48.27895, 48.26094, 48.24269, 48.22421, 48.20549, 48.18654, 
    48.16735, 48.14793, 48.12827, 48.10838, 48.08825, 48.06789, 48.04729, 
    48.02647, 48.00541, 47.98412, 47.9626, 47.94084, 47.91885, 47.89664, 
    47.87419, 47.85151, 47.82861, 47.80547, 47.78211, 47.75851, 47.7347, 
    47.71064, 47.68637, 47.66187, 47.63714, 47.61218, 47.587, 47.5616, 
    47.53596, 47.51011, 47.48403, 47.45773, 47.4312, 47.40445, 47.37748, 
    47.35029, 47.32288, 47.29524, 47.26738, 47.23931, 47.21101, 47.1825, 
    47.15377, 47.12481, 47.09565, 47.06626, 47.03666, 47.00684, 46.9768, 
    46.94655, 46.91608, 46.8854, 46.85451, 46.8234, 46.79208, 46.76054, 
    46.7288, 46.69684, 46.66467, 46.63229, 46.5997, 46.5669, 46.53389, 
    46.50068, 46.46725, 46.43362, 46.39977, 46.36573, 46.33147, 46.29701, 
    46.26235, 46.22748, 46.1924, 46.15712, 46.12164, 46.08596, 46.05008, 
    46.01398, 45.9777, 45.94121, 45.90452, 45.86763, 45.83054, 45.79325, 
    45.75577, 45.71808, 45.6802, 45.64213, 45.60386, 45.56539, 45.52672, 
    45.48787, 45.44881,
  41.14775, 41.20256, 41.25721, 41.31172, 41.36609, 41.42031, 41.47438, 
    41.52831, 41.58209, 41.63572, 41.6892, 41.74253, 41.79572, 41.84875, 
    41.90164, 41.95437, 42.00695, 42.05938, 42.11165, 42.16378, 42.21574, 
    42.26756, 42.31922, 42.37072, 42.42207, 42.47326, 42.5243, 42.57517, 
    42.62589, 42.67645, 42.72685, 42.7771, 42.82718, 42.8771, 42.92686, 
    42.97646, 43.02589, 43.07516, 43.12427, 43.17322, 43.222, 43.27061, 
    43.31906, 43.36735, 43.41547, 43.46341, 43.5112, 43.55881, 43.60626, 
    43.65353, 43.70064, 43.74757, 43.79434, 43.84093, 43.88736, 43.93361, 
    43.97968, 44.02558, 44.07131, 44.11686, 44.16224, 44.20744, 44.25247, 
    44.29731, 44.34198, 44.38648, 44.43079, 44.47493, 44.51888, 44.56266, 
    44.60625, 44.64967, 44.6929, 44.73595, 44.77881, 44.8215, 44.86399, 
    44.90631, 44.94844, 44.99038, 45.03214, 45.07371, 45.11509, 45.15628, 
    45.19729, 45.23811, 45.27874, 45.31918, 45.35943, 45.39948, 45.43935, 
    45.47902, 45.51851, 45.55779, 45.59689, 45.63579, 45.67449, 45.71301, 
    45.75132, 45.78944, 45.82736, 45.86508, 45.90261, 45.93993, 45.97706, 
    46.01399, 46.05072, 46.08725, 46.12358, 46.1597, 46.19563, 46.23135, 
    46.26687, 46.30218, 46.33729, 46.3722, 46.4069, 46.44139, 46.47569, 
    46.50977, 46.54364, 46.57731, 46.61077, 46.64402, 46.67706, 46.7099, 
    46.74252, 46.77493, 46.80713, 46.83912, 46.8709, 46.90246, 46.93381, 
    46.96495, 46.99587, 47.02658, 47.05708, 47.08735, 47.11742, 47.14726, 
    47.17689, 47.2063, 47.2355, 47.26447, 47.29323, 47.32177, 47.35009, 
    47.37819, 47.40607, 47.43372, 47.46116, 47.48837, 47.51537, 47.54214, 
    47.56868, 47.59501, 47.6211, 47.64698, 47.67263, 47.69805, 47.72325, 
    47.74822, 47.77297, 47.79749, 47.82178, 47.84584, 47.86968, 47.89328, 
    47.91666, 47.93981, 47.96273, 47.98542, 48.00788, 48.03011, 48.0521, 
    48.07387, 48.0954, 48.1167, 48.13777, 48.1586, 48.1792, 48.19957, 
    48.2197, 48.2396, 48.25927, 48.2787, 48.29789, 48.31685, 48.33557, 
    48.35405, 48.3723, 48.39031, 48.40808, 48.42562, 48.44292, 48.45998, 
    48.4768, 48.49338, 48.50972, 48.52583, 48.54169, 48.55731, 48.57269, 
    48.58783, 48.60273, 48.61739, 48.63181, 48.64598, 48.65992, 48.67361, 
    48.68706, 48.70027, 48.71323, 48.72595, 48.73843, 48.75066, 48.76265, 
    48.77439, 48.7859, 48.79715, 48.80816, 48.81893, 48.82945, 48.83973, 
    48.84975, 48.85954, 48.86908, 48.87837, 48.88742, 48.89622, 48.90477, 
    48.91307, 48.92113, 48.92895, 48.93651, 48.94383, 48.9509, 48.95773, 
    48.9643, 48.97063, 48.97671, 48.98254, 48.98812, 48.99346, 48.99854, 
    49.00338, 49.00797, 49.01231, 49.0164, 49.02025, 49.02384, 49.02719, 
    49.03028, 49.03313, 49.03573, 49.03808, 49.04018, 49.04203, 49.04363, 
    49.04498, 49.04608, 49.04694, 49.04754, 49.04789, 49.048, 49.04786, 
    49.04746, 49.04682, 49.04593, 49.04478, 49.04339, 49.04175, 49.03986, 
    49.03772, 49.03534, 49.0327, 49.02981, 49.02667, 49.02329, 49.01965, 
    49.01577, 49.01164, 49.00726, 49.00263, 48.99775, 48.99263, 48.98726, 
    48.98163, 48.97576, 48.96964, 48.96328, 48.95666, 48.9498, 48.94269, 
    48.93533, 48.92773, 48.91988, 48.91178, 48.90343, 48.89484, 48.886, 
    48.87692, 48.86758, 48.85801, 48.84819, 48.83812, 48.8278, 48.81724, 
    48.80643, 48.79539, 48.78409, 48.77255, 48.76077, 48.74874, 48.73647, 
    48.72395, 48.7112, 48.69819, 48.68495, 48.67146, 48.65773, 48.64376, 
    48.62955, 48.61509, 48.60039, 48.58545, 48.57027, 48.55486, 48.53919, 
    48.52329, 48.50715, 48.49077, 48.47415, 48.45729, 48.4402, 48.42286, 
    48.40529, 48.38748, 48.36943, 48.35115, 48.33262, 48.31387, 48.29487, 
    48.27564, 48.25617, 48.23647, 48.21654, 48.19637, 48.17596, 48.15532, 
    48.13445, 48.11335, 48.09201, 48.07044, 48.04864, 48.0266, 48.00434, 
    47.98185, 47.95912, 47.93616, 47.91298, 47.88956, 47.86592, 47.84205, 
    47.81795, 47.79362, 47.76907, 47.74429, 47.71928, 47.69404, 47.66858, 
    47.6429, 47.61699, 47.59085, 47.5645, 47.53792, 47.51111, 47.48409, 
    47.45684, 47.42936, 47.40167, 47.37376, 47.34562, 47.31727, 47.2887, 
    47.25991, 47.2309, 47.20167, 47.17222, 47.14256, 47.11267, 47.08258, 
    47.05227, 47.02174, 46.99099, 46.96004, 46.92886, 46.89748, 46.86588, 
    46.83407, 46.80205, 46.76982, 46.73737, 46.70472, 46.67185, 46.63877, 
    46.60549, 46.572, 46.5383, 46.50439, 46.47028, 46.43595, 46.40142, 
    46.36669, 46.33175, 46.29661, 46.26126, 46.22571, 46.18996, 46.154, 
    46.11784, 46.08149, 46.04493, 46.00816, 45.9712, 45.93404, 45.89668, 
    45.85913, 45.82137, 45.78342, 45.74527, 45.70692, 45.66838, 45.62965, 
    45.59072, 45.55159,
  41.24305, 41.29794, 41.35268, 41.40727, 41.46172, 41.51602, 41.57018, 
    41.62419, 41.67805, 41.73177, 41.78533, 41.83875, 41.89201, 41.94513, 
    41.9981, 42.05091, 42.10358, 42.15609, 42.20845, 42.26065, 42.3127, 
    42.3646, 42.41634, 42.46793, 42.51936, 42.57063, 42.62175, 42.67271, 
    42.72351, 42.77415, 42.82463, 42.87496, 42.92512, 42.97512, 43.02497, 
    43.07465, 43.12416, 43.17352, 43.22271, 43.27174, 43.3206, 43.3693, 
    43.41783, 43.46619, 43.51439, 43.56242, 43.61029, 43.65799, 43.70551, 
    43.75287, 43.80006, 43.84707, 43.89392, 43.94059, 43.98709, 44.03342, 
    44.07958, 44.12556, 44.17137, 44.217, 44.26245, 44.30774, 44.35284, 
    44.39777, 44.44252, 44.48709, 44.53149, 44.5757, 44.61973, 44.66359, 
    44.70726, 44.75075, 44.79406, 44.83719, 44.88013, 44.92289, 44.96547, 
    45.00786, 45.05006, 45.09208, 45.13392, 45.17556, 45.21703, 45.2583, 
    45.29938, 45.34027, 45.38098, 45.42149, 45.46181, 45.50195, 45.54189, 
    45.58164, 45.62119, 45.66055, 45.69972, 45.7387, 45.77748, 45.81606, 
    45.85445, 45.89264, 45.93063, 45.96843, 46.00603, 46.04343, 46.08062, 
    46.11763, 46.15443, 46.19102, 46.22742, 46.26362, 46.29961, 46.33541, 
    46.37099, 46.40638, 46.44156, 46.47653, 46.5113, 46.54586, 46.58022, 
    46.61437, 46.64832, 46.68205, 46.71558, 46.74889, 46.782, 46.8149, 
    46.84759, 46.88006, 46.91233, 46.94438, 46.97622, 47.00785, 47.03926, 
    47.07047, 47.10145, 47.13223, 47.16278, 47.19312, 47.22325, 47.25315, 
    47.28284, 47.31232, 47.34157, 47.37061, 47.39943, 47.42802, 47.4564, 
    47.48456, 47.51249, 47.54021, 47.5677, 47.59497, 47.62202, 47.64885, 
    47.67545, 47.70183, 47.72798, 47.75391, 47.77961, 47.80509, 47.83034, 
    47.85537, 47.88017, 47.90474, 47.92908, 47.95319, 47.97708, 48.00074, 
    48.02417, 48.04736, 48.07033, 48.09307, 48.11558, 48.13785, 48.1599, 
    48.18171, 48.20329, 48.22464, 48.24575, 48.26663, 48.28727, 48.30769, 
    48.32786, 48.34781, 48.36751, 48.38698, 48.40622, 48.42522, 48.44398, 
    48.46251, 48.48079, 48.49884, 48.51665, 48.53423, 48.55156, 48.56866, 
    48.58552, 48.60214, 48.61852, 48.63465, 48.65055, 48.66621, 48.68163, 
    48.6968, 48.71173, 48.72643, 48.74088, 48.75508, 48.76905, 48.78277, 
    48.79625, 48.80948, 48.82248, 48.83522, 48.84773, 48.85999, 48.87201, 
    48.88378, 48.8953, 48.90659, 48.91762, 48.92841, 48.93895, 48.94925, 
    48.9593, 48.96911, 48.97867, 48.98799, 48.99705, 49.00587, 49.01445, 
    49.02277, 49.03085, 49.03868, 49.04626, 49.0536, 49.06068, 49.06752, 
    49.07411, 49.08045, 49.08654, 49.09239, 49.09798, 49.10333, 49.10843, 
    49.11328, 49.11788, 49.12223, 49.12633, 49.13018, 49.13379, 49.13714, 
    49.14024, 49.1431, 49.1457, 49.14806, 49.15016, 49.15201, 49.15362, 
    49.15497, 49.15608, 49.15693, 49.15754, 49.15789, 49.158, 49.15786, 
    49.15746, 49.15681, 49.15592, 49.15478, 49.15338, 49.15174, 49.14984, 
    49.1477, 49.14531, 49.14266, 49.13977, 49.13662, 49.13323, 49.12959, 
    49.1257, 49.12156, 49.11717, 49.11253, 49.10764, 49.1025, 49.09712, 
    49.09148, 49.0856, 49.07946, 49.07309, 49.06646, 49.05958, 49.05245, 
    49.04508, 49.03746, 49.02959, 49.02147, 49.01311, 49.00449, 48.99564, 
    48.98653, 48.97718, 48.96758, 48.95773, 48.94764, 48.9373, 48.92672, 
    48.91589, 48.90482, 48.8935, 48.88193, 48.87012, 48.85807, 48.84577, 
    48.83323, 48.82044, 48.80741, 48.79413, 48.78061, 48.76685, 48.75285, 
    48.73861, 48.72412, 48.70938, 48.69442, 48.6792, 48.66375, 48.64805, 
    48.63212, 48.61594, 48.59953, 48.58287, 48.56597, 48.54884, 48.53146, 
    48.51385, 48.496, 48.47792, 48.45959, 48.44103, 48.42223, 48.40319, 
    48.38392, 48.36441, 48.34467, 48.32469, 48.30447, 48.28402, 48.26334, 
    48.24242, 48.22128, 48.19989, 48.17828, 48.15643, 48.13435, 48.11203, 
    48.08949, 48.06672, 48.04371, 48.02048, 47.99701, 47.97332, 47.94939, 
    47.92524, 47.90086, 47.87626, 47.85143, 47.82636, 47.80107, 47.77556, 
    47.74982, 47.72386, 47.69767, 47.67126, 47.64462, 47.61776, 47.59068, 
    47.56337, 47.53584, 47.50809, 47.48012, 47.45193, 47.42352, 47.39488, 
    47.36603, 47.33696, 47.30767, 47.27816, 47.24844, 47.21849, 47.18834, 
    47.15796, 47.12737, 47.09657, 47.06554, 47.03431, 47.00286, 46.9712, 
    46.93933, 46.90724, 46.87494, 46.84243, 46.80971, 46.77678, 46.74364, 
    46.71029, 46.67673, 46.64296, 46.60899, 46.5748, 46.54041, 46.50581, 
    46.47101, 46.436, 46.40079, 46.36538, 46.32976, 46.29393, 46.25791, 
    46.22168, 46.18525, 46.14862, 46.11179, 46.07475, 46.03752, 46.00009, 
    45.96246, 45.92463, 45.88661, 45.84839, 45.80997, 45.77135, 45.73254, 
    45.69354, 45.65434,
  41.33831, 41.39327, 41.4481, 41.50277, 41.5573, 41.61169, 41.66593, 
    41.72002, 41.77397, 41.82777, 41.88142, 41.93491, 41.98827, 42.04147, 
    42.09451, 42.14741, 42.20016, 42.25275, 42.30519, 42.35748, 42.40961, 
    42.46159, 42.51342, 42.56509, 42.6166, 42.66796, 42.71916, 42.7702, 
    42.82109, 42.87181, 42.92238, 42.97278, 43.02303, 43.07312, 43.12304, 
    43.1728, 43.2224, 43.27184, 43.32111, 43.37022, 43.41916, 43.46794, 
    43.51656, 43.565, 43.61329, 43.6614, 43.70934, 43.75712, 43.80473, 
    43.85217, 43.89943, 43.94653, 43.99346, 44.04021, 44.08679, 44.1332, 
    44.17944, 44.2255, 44.27139, 44.3171, 44.36264, 44.408, 44.45319, 
    44.49819, 44.54302, 44.58767, 44.63214, 44.67644, 44.72055, 44.76448, 
    44.80824, 44.8518, 44.89519, 44.9384, 44.98142, 45.02425, 45.06691, 
    45.10938, 45.15166, 45.19376, 45.23567, 45.27739, 45.31893, 45.36028, 
    45.40144, 45.44241, 45.48318, 45.52378, 45.56417, 45.60438, 45.6444, 
    45.68422, 45.72385, 45.76329, 45.80253, 45.84158, 45.88043, 45.91909, 
    45.95755, 45.99581, 46.03388, 46.07175, 46.10942, 46.14689, 46.18416, 
    46.22123, 46.25811, 46.29478, 46.33125, 46.36751, 46.40358, 46.43944, 
    46.4751, 46.51055, 46.5458, 46.58084, 46.61568, 46.65031, 46.68474, 
    46.71896, 46.75297, 46.78677, 46.82036, 46.85374, 46.88692, 46.91988, 
    46.95264, 46.98518, 47.01751, 47.04963, 47.08153, 47.11322, 47.1447, 
    47.17597, 47.20702, 47.23785, 47.26847, 47.29887, 47.32906, 47.35903, 
    47.38878, 47.41832, 47.44763, 47.47673, 47.5056, 47.53426, 47.56269, 
    47.59091, 47.61891, 47.64668, 47.67423, 47.70156, 47.72866, 47.75554, 
    47.7822, 47.80864, 47.83484, 47.86083, 47.88659, 47.91212, 47.93742, 
    47.9625, 47.98735, 48.01197, 48.03637, 48.06054, 48.08447, 48.10818, 
    48.13166, 48.15491, 48.17793, 48.20071, 48.22327, 48.24559, 48.26768, 
    48.28954, 48.31117, 48.33256, 48.35372, 48.37465, 48.39534, 48.41579, 
    48.43601, 48.456, 48.47575, 48.49526, 48.51454, 48.53358, 48.55238, 
    48.57095, 48.58928, 48.60737, 48.62522, 48.64283, 48.66021, 48.67734, 
    48.69423, 48.71089, 48.7273, 48.74348, 48.75941, 48.7751, 48.79055, 
    48.80576, 48.82073, 48.83545, 48.84993, 48.86417, 48.87817, 48.89192, 
    48.90543, 48.9187, 48.93172, 48.9445, 48.95703, 48.96931, 48.98136, 
    48.99316, 49.00471, 49.01601, 49.02708, 49.03789, 49.04846, 49.05878, 
    49.06886, 49.07869, 49.08826, 49.0976, 49.10669, 49.11553, 49.12412, 
    49.13246, 49.14056, 49.14841, 49.15601, 49.16336, 49.17046, 49.17731, 
    49.18392, 49.19028, 49.19638, 49.20224, 49.20785, 49.21321, 49.21832, 
    49.22318, 49.22779, 49.23215, 49.23626, 49.24012, 49.24373, 49.24709, 
    49.2502, 49.25306, 49.25567, 49.25803, 49.26014, 49.262, 49.26361, 
    49.26497, 49.26608, 49.26693, 49.26754, 49.26789, 49.268, 49.26785, 
    49.26746, 49.26681, 49.26591, 49.26477, 49.26337, 49.26172, 49.25982, 
    49.25768, 49.25528, 49.25262, 49.24973, 49.24658, 49.24318, 49.23952, 
    49.23563, 49.23148, 49.22707, 49.22243, 49.21753, 49.21238, 49.20698, 
    49.20133, 49.19543, 49.18929, 49.18289, 49.17625, 49.16935, 49.16221, 
    49.15482, 49.14718, 49.13929, 49.13116, 49.12278, 49.11415, 49.10527, 
    49.09614, 49.08677, 49.07714, 49.06728, 49.05716, 49.0468, 49.0362, 
    49.02534, 49.01424, 49.0029, 48.99131, 48.97947, 48.96739, 48.95506, 
    48.94249, 48.92968, 48.91661, 48.90331, 48.88976, 48.87597, 48.86194, 
    48.84766, 48.83314, 48.81838, 48.80337, 48.78812, 48.77264, 48.7569, 
    48.74094, 48.72472, 48.70827, 48.69158, 48.67464, 48.65747, 48.64006, 
    48.62241, 48.60452, 48.5864, 48.56803, 48.54942, 48.53058, 48.51151, 
    48.49219, 48.47264, 48.45285, 48.43283, 48.41257, 48.39208, 48.37135, 
    48.35039, 48.32919, 48.30776, 48.2861, 48.2642, 48.24208, 48.21972, 
    48.19712, 48.1743, 48.15125, 48.12796, 48.10445, 48.0807, 48.05673, 
    48.03253, 48.00809, 47.98344, 47.95855, 47.93343, 47.90809, 47.88253, 
    47.85673, 47.83072, 47.80447, 47.778, 47.75131, 47.72439, 47.69725, 
    47.66989, 47.6423, 47.61449, 47.58646, 47.55821, 47.52974, 47.50105, 
    47.47214, 47.44301, 47.41366, 47.38409, 47.3543, 47.3243, 47.29408, 
    47.26364, 47.23299, 47.20212, 47.17104, 47.13974, 47.10823, 47.0765, 
    47.04456, 47.01241, 46.98005, 46.94747, 46.91468, 46.88169, 46.84848, 
    46.81506, 46.78144, 46.7476, 46.71356, 46.67931, 46.64485, 46.61018, 
    46.57531, 46.54024, 46.50496, 46.46947, 46.43378, 46.39788, 46.36179, 
    46.32549, 46.28899, 46.25229, 46.21538, 46.17828, 46.14098, 46.10347, 
    46.06577, 46.02787, 45.98977, 45.95148, 45.91299, 45.8743, 45.83541, 
    45.79634, 45.75706,
  41.43351, 41.48856, 41.54347, 41.59823, 41.65284, 41.70731, 41.76164, 
    41.81581, 41.86984, 41.92372, 41.97746, 42.03104, 42.08447, 42.13775, 
    42.19089, 42.24387, 42.2967, 42.34937, 42.4019, 42.45427, 42.50649, 
    42.55855, 42.61046, 42.66221, 42.71381, 42.76525, 42.81653, 42.86765, 
    42.91862, 42.96943, 43.02008, 43.07057, 43.1209, 43.17106, 43.22107, 
    43.27092, 43.32059, 43.37011, 43.41947, 43.46866, 43.51769, 43.56655, 
    43.61525, 43.66377, 43.71214, 43.76033, 43.80836, 43.85622, 43.9039, 
    43.95142, 43.99878, 44.04595, 44.09296, 44.13979, 44.18646, 44.23295, 
    44.27927, 44.32541, 44.37138, 44.41717, 44.46279, 44.50823, 44.55349, 
    44.59858, 44.64349, 44.68822, 44.73277, 44.77714, 44.82133, 44.86535, 
    44.90918, 44.95282, 44.99629, 45.03957, 45.08267, 45.12559, 45.16832, 
    45.21087, 45.25323, 45.2954, 45.33739, 45.37919, 45.4208, 45.46223, 
    45.50346, 45.54451, 45.58537, 45.62603, 45.6665, 45.70679, 45.74688, 
    45.78678, 45.82648, 45.86599, 45.90531, 45.94443, 45.98336, 46.02209, 
    46.06062, 46.09896, 46.1371, 46.17504, 46.21279, 46.25033, 46.28767, 
    46.32482, 46.36176, 46.3985, 46.43504, 46.47138, 46.50751, 46.54345, 
    46.57917, 46.6147, 46.65002, 46.68513, 46.72004, 46.75474, 46.78923, 
    46.82352, 46.8576, 46.89146, 46.92513, 46.95858, 46.99182, 47.02485, 
    47.05767, 47.09027, 47.12267, 47.15485, 47.18682, 47.21858, 47.25012, 
    47.28145, 47.31256, 47.34346, 47.37414, 47.40461, 47.43486, 47.46489, 
    47.4947, 47.5243, 47.55367, 47.58283, 47.61176, 47.64048, 47.66898, 
    47.69725, 47.7253, 47.75314, 47.78074, 47.80813, 47.83529, 47.86223, 
    47.88894, 47.91543, 47.9417, 47.96774, 47.99355, 48.01913, 48.04449, 
    48.06962, 48.09452, 48.1192, 48.14365, 48.16787, 48.19186, 48.21561, 
    48.23914, 48.26244, 48.28551, 48.30835, 48.33095, 48.35332, 48.37546, 
    48.39737, 48.41904, 48.44048, 48.46168, 48.48265, 48.50339, 48.52389, 
    48.54416, 48.56419, 48.58398, 48.60353, 48.62285, 48.64194, 48.66078, 
    48.67939, 48.69775, 48.71589, 48.73378, 48.75143, 48.76884, 48.78601, 
    48.80294, 48.81964, 48.83609, 48.85229, 48.86826, 48.88399, 48.89948, 
    48.91472, 48.92972, 48.94448, 48.95899, 48.97326, 48.98729, 49.00107, 
    49.01461, 49.02791, 49.04096, 49.05376, 49.06632, 49.07864, 49.09071, 
    49.10253, 49.11411, 49.12544, 49.13653, 49.14737, 49.15796, 49.1683, 
    49.1784, 49.18826, 49.19786, 49.20721, 49.21632, 49.22518, 49.23379, 
    49.24215, 49.25027, 49.25814, 49.26575, 49.27312, 49.28024, 49.28711, 
    49.29373, 49.3001, 49.30622, 49.31209, 49.31771, 49.32308, 49.32821, 
    49.33308, 49.3377, 49.34207, 49.34619, 49.35006, 49.35368, 49.35704, 
    49.36016, 49.36303, 49.36564, 49.36801, 49.37012, 49.37199, 49.3736, 
    49.37496, 49.37607, 49.37693, 49.37754, 49.3779, 49.378, 49.37785, 
    49.37746, 49.37681, 49.37591, 49.37476, 49.37336, 49.37171, 49.3698, 
    49.36765, 49.36525, 49.36259, 49.35968, 49.35653, 49.35312, 49.34946, 
    49.34555, 49.34139, 49.33698, 49.33232, 49.32741, 49.32225, 49.31684, 
    49.31118, 49.30527, 49.29911, 49.2927, 49.28604, 49.27913, 49.27197, 
    49.26456, 49.25691, 49.249, 49.24085, 49.23244, 49.2238, 49.2149, 
    49.20575, 49.19635, 49.18671, 49.17682, 49.16669, 49.1563, 49.14567, 
    49.13479, 49.12367, 49.1123, 49.10068, 49.08882, 49.07671, 49.06435, 
    49.05175, 49.03891, 49.02582, 49.01249, 48.99891, 48.98508, 48.97102, 
    48.95671, 48.94216, 48.92736, 48.91232, 48.89704, 48.88152, 48.86575, 
    48.84975, 48.8335, 48.81701, 48.80028, 48.78331, 48.7661, 48.74865, 
    48.73096, 48.71303, 48.69487, 48.67646, 48.65781, 48.63893, 48.61981, 
    48.60046, 48.58086, 48.56103, 48.54097, 48.52066, 48.50013, 48.47935, 
    48.45834, 48.4371, 48.41563, 48.39392, 48.37197, 48.3498, 48.32739, 
    48.30475, 48.28188, 48.25877, 48.23544, 48.21187, 48.18808, 48.16405, 
    48.1398, 48.11531, 48.0906, 48.06566, 48.04049, 48.0151, 47.98948, 
    47.96363, 47.93756, 47.91125, 47.88473, 47.85798, 47.83101, 47.80381, 
    47.77639, 47.74874, 47.72088, 47.69279, 47.66448, 47.63595, 47.6072, 
    47.57823, 47.54904, 47.51963, 47.49, 47.46015, 47.43009, 47.3998, 
    47.3693, 47.33859, 47.30766, 47.27651, 47.24515, 47.21357, 47.18178, 
    47.14978, 47.11756, 47.08513, 47.05249, 47.01964, 46.98657, 46.9533, 
    46.91982, 46.88612, 46.85222, 46.81811, 46.78379, 46.74926, 46.71453, 
    46.67959, 46.64444, 46.60909, 46.57354, 46.53778, 46.50181, 46.46564, 
    46.42928, 46.3927, 46.35593, 46.31895, 46.28178, 46.2444, 46.20683, 
    46.16906, 46.13108, 46.09291, 46.05454, 46.01598, 45.97721, 45.93826, 
    45.89911, 45.85976,
  41.52867, 41.58381, 41.63879, 41.69364, 41.74834, 41.80289, 41.8573, 
    41.91156, 41.96567, 42.01963, 42.07345, 42.12712, 42.18063, 42.234, 
    42.28722, 42.34028, 42.39319, 42.44595, 42.49856, 42.55101, 42.60331, 
    42.65546, 42.70745, 42.75929, 42.81097, 42.86249, 42.91386, 42.96507, 
    43.01611, 43.06701, 43.11774, 43.16831, 43.21872, 43.26897, 43.31906, 
    43.36899, 43.41875, 43.46835, 43.51779, 43.56706, 43.61617, 43.66512, 
    43.71389, 43.7625, 43.81095, 43.85923, 43.90733, 43.95527, 44.00304, 
    44.05064, 44.09808, 44.14534, 44.19242, 44.23934, 44.28609, 44.33266, 
    44.37906, 44.42528, 44.47132, 44.5172, 44.5629, 44.60842, 44.65376, 
    44.69893, 44.74392, 44.78873, 44.83336, 44.87781, 44.92208, 44.96618, 
    45.01008, 45.05381, 45.09735, 45.14072, 45.1839, 45.22689, 45.2697, 
    45.31232, 45.35476, 45.39701, 45.43908, 45.48096, 45.52265, 45.56415, 
    45.60546, 45.64658, 45.68752, 45.72826, 45.76881, 45.80917, 45.84933, 
    45.88931, 45.92908, 45.96867, 46.00806, 46.04726, 46.08626, 46.12506, 
    46.16367, 46.20208, 46.2403, 46.27831, 46.31613, 46.35374, 46.39116, 
    46.42838, 46.46539, 46.5022, 46.53881, 46.57523, 46.61143, 46.64743, 
    46.68323, 46.71883, 46.75421, 46.78939, 46.82437, 46.85914, 46.8937, 
    46.92806, 46.9622, 46.99614, 47.02987, 47.06339, 47.09669, 47.12979, 
    47.16268, 47.19535, 47.22781, 47.26006, 47.2921, 47.32392, 47.35552, 
    47.38692, 47.41809, 47.44905, 47.4798, 47.51033, 47.54063, 47.57073, 
    47.6006, 47.63026, 47.65969, 47.68891, 47.71791, 47.74669, 47.77524, 
    47.80357, 47.83168, 47.85957, 47.88724, 47.91468, 47.9419, 47.9689, 
    47.99567, 48.02221, 48.04853, 48.07463, 48.10049, 48.12613, 48.15155, 
    48.17673, 48.20169, 48.22642, 48.25092, 48.27519, 48.29923, 48.32304, 
    48.34661, 48.36996, 48.39308, 48.41597, 48.43862, 48.46104, 48.48323, 
    48.50518, 48.5269, 48.54839, 48.56964, 48.59065, 48.61143, 48.63198, 
    48.65229, 48.67236, 48.6922, 48.7118, 48.73116, 48.75028, 48.76917, 
    48.78782, 48.80623, 48.8244, 48.84233, 48.86002, 48.87747, 48.89468, 
    48.91165, 48.92838, 48.94487, 48.96111, 48.97712, 48.99287, 49.0084, 
    49.02367, 49.0387, 49.05349, 49.06804, 49.08234, 49.09641, 49.11022, 
    49.12379, 49.13711, 49.15019, 49.16303, 49.17562, 49.18796, 49.20006, 
    49.21191, 49.22351, 49.23487, 49.24598, 49.25684, 49.26746, 49.27783, 
    49.28795, 49.29782, 49.30745, 49.31683, 49.32595, 49.33483, 49.34346, 
    49.35184, 49.35998, 49.36786, 49.3755, 49.38288, 49.39001, 49.3969, 
    49.40353, 49.40992, 49.41605, 49.42194, 49.42757, 49.43296, 49.43809, 
    49.44297, 49.44761, 49.45198, 49.45612, 49.45999, 49.46362, 49.467, 
    49.47012, 49.47299, 49.47562, 49.47799, 49.48011, 49.48197, 49.48359, 
    49.48495, 49.48606, 49.48693, 49.48754, 49.48789, 49.488, 49.48785, 
    49.48746, 49.48681, 49.4859, 49.48475, 49.48335, 49.48169, 49.47979, 
    49.47763, 49.47522, 49.47256, 49.46964, 49.46648, 49.46306, 49.4594, 
    49.45548, 49.45131, 49.44689, 49.44222, 49.43729, 49.43212, 49.4267, 
    49.42102, 49.4151, 49.40893, 49.4025, 49.39583, 49.3889, 49.38173, 
    49.37431, 49.36663, 49.35871, 49.35054, 49.34211, 49.33344, 49.32452, 
    49.31536, 49.30594, 49.29628, 49.28637, 49.2762, 49.2658, 49.25514, 
    49.24424, 49.23309, 49.22169, 49.21005, 49.19816, 49.18602, 49.17364, 
    49.16101, 49.14814, 49.13502, 49.12166, 49.10805, 49.0942, 49.0801, 
    49.06576, 49.05117, 49.03634, 49.02127, 49.00595, 48.9904, 48.9746, 
    48.95856, 48.94227, 48.92575, 48.90898, 48.89197, 48.87473, 48.85723, 
    48.83951, 48.82154, 48.80333, 48.78489, 48.7662, 48.74728, 48.72811, 
    48.70871, 48.68908, 48.6692, 48.64909, 48.62875, 48.60816, 48.58735, 
    48.56629, 48.545, 48.52348, 48.50172, 48.47973, 48.45751, 48.43505, 
    48.41236, 48.38944, 48.36629, 48.3429, 48.31929, 48.29544, 48.27136, 
    48.24706, 48.22252, 48.19776, 48.17276, 48.14754, 48.12209, 48.09642, 
    48.07051, 48.04438, 48.01803, 47.99145, 47.96464, 47.93761, 47.91036, 
    47.88288, 47.85518, 47.82726, 47.79911, 47.77074, 47.74215, 47.71334, 
    47.68431, 47.65505, 47.62558, 47.59589, 47.56598, 47.53585, 47.50551, 
    47.47495, 47.44417, 47.41317, 47.38197, 47.35054, 47.3189, 47.28704, 
    47.25497, 47.22269, 47.1902, 47.15749, 47.12457, 47.09144, 47.0581, 
    47.02455, 46.99079, 46.95682, 46.92264, 46.88825, 46.85366, 46.81885, 
    46.78384, 46.74863, 46.71321, 46.67758, 46.64175, 46.60572, 46.56948, 
    46.53304, 46.4964, 46.45955, 46.4225, 46.38525, 46.34781, 46.31016, 
    46.27231, 46.23426, 46.19602, 46.15758, 46.11894, 46.0801, 46.04107, 
    46.00185, 45.96242,
  41.62378, 41.679, 41.73407, 41.789, 41.84378, 41.89842, 41.95291, 42.00726, 
    42.06145, 42.1155, 42.1694, 42.22315, 42.27675, 42.3302, 42.3835, 
    42.43665, 42.48964, 42.54248, 42.59518, 42.64772, 42.7001, 42.75233, 
    42.8044, 42.85632, 42.90808, 42.95969, 43.01114, 43.06243, 43.11356, 
    43.16454, 43.21535, 43.26601, 43.3165, 43.36684, 43.41701, 43.46702, 
    43.51686, 43.56655, 43.61607, 43.66542, 43.71462, 43.76364, 43.8125, 
    43.86119, 43.90972, 43.95808, 44.00627, 44.05429, 44.10215, 44.14983, 
    44.19734, 44.24468, 44.29185, 44.33885, 44.38568, 44.43233, 44.47881, 
    44.52511, 44.57124, 44.6172, 44.66298, 44.70858, 44.754, 44.79925, 
    44.84431, 44.88921, 44.93392, 44.97845, 45.0228, 45.06697, 45.11096, 
    45.15476, 45.19839, 45.24183, 45.28508, 45.32816, 45.37104, 45.41375, 
    45.45626, 45.49859, 45.54074, 45.58269, 45.62446, 45.66604, 45.70743, 
    45.74863, 45.78963, 45.83045, 45.87108, 45.91151, 45.95176, 45.99181, 
    46.03166, 46.07132, 46.11079, 46.15006, 46.18913, 46.22801, 46.2667, 
    46.30518, 46.34347, 46.38155, 46.41944, 46.45713, 46.49462, 46.53191, 
    46.569, 46.60588, 46.64257, 46.67905, 46.71532, 46.7514, 46.78726, 
    46.82293, 46.85839, 46.89364, 46.92868, 46.96352, 46.99815, 47.03258, 
    47.06679, 47.1008, 47.13459, 47.16817, 47.20155, 47.23471, 47.26767, 
    47.30041, 47.33294, 47.36525, 47.39735, 47.42923, 47.46091, 47.49236, 
    47.5236, 47.55463, 47.58543, 47.61602, 47.6464, 47.67655, 47.70649, 
    47.73621, 47.76571, 47.79498, 47.82404, 47.85287, 47.88149, 47.90988, 
    47.93805, 47.966, 47.99372, 48.02122, 48.0485, 48.07555, 48.10238, 
    48.12898, 48.15536, 48.18151, 48.20743, 48.23312, 48.25859, 48.28383, 
    48.30884, 48.33362, 48.35817, 48.3825, 48.40659, 48.43045, 48.45408, 
    48.47748, 48.50064, 48.52358, 48.54628, 48.56875, 48.59098, 48.61298, 
    48.63475, 48.65628, 48.67758, 48.69864, 48.71947, 48.74006, 48.76041, 
    48.78053, 48.80041, 48.82005, 48.83946, 48.85863, 48.87755, 48.89624, 
    48.91469, 48.9329, 48.95087, 48.9686, 48.98609, 49.00334, 49.02035, 
    49.03711, 49.05364, 49.06992, 49.08596, 49.10175, 49.11731, 49.13262, 
    49.14769, 49.16251, 49.17709, 49.19143, 49.20551, 49.21936, 49.23296, 
    49.24632, 49.25943, 49.27229, 49.2849, 49.29728, 49.3094, 49.32128, 
    49.33291, 49.34429, 49.35543, 49.36632, 49.37696, 49.38735, 49.39749, 
    49.40739, 49.41703, 49.42643, 49.43558, 49.44448, 49.45313, 49.46153, 
    49.46968, 49.47758, 49.48524, 49.49264, 49.49979, 49.50669, 49.51334, 
    49.51974, 49.52589, 49.53179, 49.53744, 49.54283, 49.54798, 49.55287, 
    49.55751, 49.5619, 49.56604, 49.56993, 49.57356, 49.57695, 49.58008, 
    49.58296, 49.58559, 49.58796, 49.59009, 49.59196, 49.59358, 49.59494, 
    49.59606, 49.59692, 49.59753, 49.59789, 49.598, 49.59785, 49.59745, 
    49.59681, 49.5959, 49.59475, 49.59334, 49.59168, 49.58977, 49.5876, 
    49.58519, 49.58252, 49.5796, 49.57643, 49.57301, 49.56933, 49.5654, 
    49.56123, 49.55679, 49.55211, 49.54718, 49.542, 49.53656, 49.53087, 
    49.52494, 49.51875, 49.51231, 49.50562, 49.49868, 49.49149, 49.48404, 
    49.47635, 49.46841, 49.46022, 49.45178, 49.44309, 49.43415, 49.42496, 
    49.41553, 49.40584, 49.3959, 49.38572, 49.37529, 49.36461, 49.35368, 
    49.34251, 49.33109, 49.31942, 49.3075, 49.29534, 49.28292, 49.27027, 
    49.25737, 49.24422, 49.23082, 49.21719, 49.2033, 49.18917, 49.1748, 
    49.16018, 49.14532, 49.13021, 49.11486, 49.09927, 49.08344, 49.06736, 
    49.05104, 49.03448, 49.01767, 49.00063, 48.98334, 48.96581, 48.94804, 
    48.93004, 48.91179, 48.8933, 48.87458, 48.85561, 48.83641, 48.81696, 
    48.79728, 48.77737, 48.75721, 48.73682, 48.71619, 48.69533, 48.67423, 
    48.65289, 48.63132, 48.60952, 48.58748, 48.56521, 48.54271, 48.51997, 
    48.49699, 48.47379, 48.45036, 48.42669, 48.40279, 48.37866, 48.35431, 
    48.32972, 48.3049, 48.27985, 48.25458, 48.22907, 48.20334, 48.17738, 
    48.1512, 48.12479, 48.09815, 48.07129, 48.0442, 48.01689, 47.98935, 
    47.96159, 47.93361, 47.90541, 47.87698, 47.84833, 47.81946, 47.79036, 
    47.76105, 47.73152, 47.70177, 47.6718, 47.64161, 47.6112, 47.58057, 
    47.54973, 47.51867, 47.4874, 47.45591, 47.42421, 47.39228, 47.36015, 
    47.3278, 47.29524, 47.26247, 47.22948, 47.19629, 47.16288, 47.12926, 
    47.09543, 47.06139, 47.02715, 46.99269, 46.95802, 46.92315, 46.88808, 
    46.85279, 46.8173, 46.7816, 46.7457, 46.7096, 46.67329, 46.63678, 
    46.60006, 46.56314, 46.52602, 46.4887, 46.45118, 46.41346, 46.37554, 
    46.33742, 46.29911, 46.26059, 46.22188, 46.18297, 46.14386, 46.10456, 
    46.06506,
  41.71885, 41.77415, 41.82931, 41.88432, 41.93919, 41.9939, 42.04848, 
    42.10291, 42.15718, 42.21132, 42.2653, 42.31913, 42.37282, 42.42635, 
    42.47974, 42.53297, 42.58605, 42.63897, 42.69175, 42.74437, 42.79684, 
    42.84915, 42.90131, 42.95331, 43.00516, 43.05685, 43.10838, 43.15976, 
    43.21097, 43.26203, 43.31293, 43.36367, 43.41424, 43.46466, 43.51492, 
    43.56501, 43.61494, 43.66471, 43.71431, 43.76375, 43.81302, 43.86213, 
    43.91107, 43.95985, 44.00846, 44.0569, 44.10517, 44.15327, 44.20121, 
    44.24897, 44.29657, 44.34399, 44.39124, 44.43832, 44.48523, 44.53196, 
    44.57852, 44.62491, 44.67112, 44.71716, 44.76301, 44.8087, 44.8542, 
    44.89953, 44.94468, 44.98965, 45.03444, 45.07905, 45.12348, 45.16773, 
    45.2118, 45.25568, 45.29939, 45.34291, 45.38624, 45.42939, 45.47236, 
    45.51514, 45.55774, 45.60014, 45.64236, 45.68439, 45.72624, 45.76789, 
    45.80936, 45.85064, 45.89172, 45.93262, 45.97332, 46.01383, 46.05415, 
    46.09428, 46.1342, 46.17394, 46.21349, 46.25283, 46.29198, 46.33093, 
    46.36969, 46.40825, 46.44661, 46.48477, 46.52273, 46.56049, 46.59806, 
    46.63542, 46.67258, 46.70953, 46.74629, 46.78284, 46.81919, 46.85533, 
    46.89127, 46.92701, 46.96254, 46.99786, 47.03297, 47.06788, 47.10258, 
    47.13707, 47.17136, 47.20543, 47.23929, 47.27295, 47.30639, 47.33962, 
    47.37263, 47.40544, 47.43803, 47.47042, 47.50258, 47.53453, 47.56627, 
    47.59779, 47.62909, 47.66018, 47.69105, 47.72171, 47.75214, 47.78236, 
    47.81236, 47.84214, 47.8717, 47.90104, 47.93015, 47.95905, 47.98772, 
    48.01617, 48.0444, 48.07241, 48.10019, 48.12775, 48.15509, 48.1822, 
    48.20908, 48.23574, 48.26217, 48.28837, 48.31435, 48.3401, 48.36562, 
    48.39091, 48.41598, 48.44081, 48.46542, 48.48979, 48.51394, 48.53785, 
    48.56153, 48.58498, 48.6082, 48.63118, 48.65393, 48.67645, 48.69873, 
    48.72078, 48.7426, 48.76418, 48.78552, 48.80663, 48.8275, 48.84813, 
    48.86853, 48.88869, 48.90862, 48.9283, 48.94775, 48.96696, 48.98593, 
    49.00466, 49.02315, 49.0414, 49.05941, 49.07718, 49.09471, 49.112, 
    49.12904, 49.14584, 49.1624, 49.17872, 49.1948, 49.21063, 49.22622, 
    49.24156, 49.25666, 49.27152, 49.28613, 49.3005, 49.31462, 49.3285, 
    49.34213, 49.35551, 49.36865, 49.38155, 49.39419, 49.40659, 49.41874, 
    49.43064, 49.4423, 49.45371, 49.46487, 49.47579, 49.48645, 49.49687, 
    49.50703, 49.51695, 49.52662, 49.53604, 49.54521, 49.55413, 49.5628, 
    49.57122, 49.57939, 49.58731, 49.59498, 49.6024, 49.60957, 49.61648, 
    49.62315, 49.62956, 49.63573, 49.64164, 49.6473, 49.65271, 49.65786, 
    49.66277, 49.66742, 49.67182, 49.67597, 49.67986, 49.68351, 49.6869, 
    49.69004, 49.69292, 49.69556, 49.69794, 49.70007, 49.70195, 49.70357, 
    49.70494, 49.70605, 49.70692, 49.70753, 49.70789, 49.708, 49.70785, 
    49.70745, 49.7068, 49.7059, 49.70474, 49.70333, 49.70166, 49.69975, 
    49.69758, 49.69516, 49.69249, 49.68956, 49.68638, 49.68295, 49.67926, 
    49.67533, 49.67114, 49.6667, 49.66201, 49.65706, 49.65187, 49.64642, 
    49.64072, 49.63477, 49.62856, 49.62211, 49.61541, 49.60845, 49.60124, 
    49.59378, 49.58607, 49.57812, 49.5699, 49.56145, 49.55274, 49.54378, 
    49.53457, 49.52511, 49.5154, 49.50544, 49.49524, 49.48478, 49.47408, 
    49.46312, 49.45192, 49.44048, 49.42878, 49.41684, 49.40464, 49.39221, 
    49.37952, 49.36659, 49.35341, 49.33999, 49.32632, 49.3124, 49.29824, 
    49.28384, 49.26919, 49.25429, 49.23915, 49.22377, 49.20814, 49.19227, 
    49.17616, 49.1598, 49.1432, 49.12636, 49.10928, 49.09195, 49.07438, 
    49.05658, 49.03853, 49.02024, 49.00171, 48.98294, 48.96394, 48.94469, 
    48.92521, 48.90548, 48.88552, 48.86532, 48.84489, 48.82421, 48.8033, 
    48.78216, 48.76078, 48.73916, 48.71731, 48.69522, 48.6729, 48.65034, 
    48.62756, 48.60454, 48.58128, 48.5578, 48.53408, 48.51013, 48.48595, 
    48.46154, 48.4369, 48.41203, 48.38693, 48.3616, 48.33604, 48.31026, 
    48.28424, 48.258, 48.23154, 48.20484, 48.17792, 48.15078, 48.12341, 
    48.09581, 48.068, 48.03996, 48.01169, 47.9832, 47.95449, 47.92556, 
    47.89641, 47.86703, 47.83744, 47.80763, 47.7776, 47.74734, 47.71687, 
    47.68618, 47.65528, 47.62416, 47.59282, 47.56126, 47.52949, 47.49751, 
    47.46531, 47.4329, 47.40027, 47.36743, 47.33437, 47.30111, 47.26764, 
    47.23395, 47.20005, 47.16595, 47.13163, 47.09711, 47.06237, 47.02743, 
    46.99228, 46.95693, 46.92137, 46.8856, 46.84963, 46.81345, 46.77707, 
    46.74049, 46.7037, 46.66671, 46.62952, 46.59213, 46.55453, 46.51674, 
    46.47875, 46.44056, 46.40216, 46.36357, 46.32478, 46.2858, 46.24662, 
    46.20724, 46.16767,
  41.81387, 41.86925, 41.92449, 41.97959, 42.03454, 42.08934, 42.144, 
    42.19851, 42.25288, 42.30709, 42.36116, 42.41507, 42.46884, 42.52246, 
    42.57593, 42.62924, 42.68241, 42.73542, 42.78828, 42.84098, 42.89354, 
    42.94593, 42.99817, 43.05026, 43.10219, 43.15396, 43.20558, 43.25704, 
    43.30834, 43.35948, 43.41046, 43.46128, 43.51194, 43.56244, 43.61278, 
    43.66296, 43.71297, 43.76282, 43.81251, 43.86203, 43.91138, 43.96058, 
    44.0096, 44.05846, 44.10715, 44.15567, 44.20403, 44.25222, 44.30023, 
    44.34808, 44.39576, 44.44326, 44.4906, 44.53776, 44.58475, 44.63156, 
    44.6782, 44.72467, 44.77096, 44.81708, 44.86302, 44.90878, 44.95436, 
    44.99977, 45.04501, 45.09005, 45.13493, 45.17962, 45.22413, 45.26846, 
    45.3126, 45.35657, 45.40035, 45.44395, 45.48737, 45.53059, 45.57364, 
    45.6165, 45.65917, 45.70166, 45.74396, 45.78607, 45.82799, 45.86972, 
    45.91127, 45.95262, 45.99379, 46.03476, 46.07553, 46.11612, 46.15652, 
    46.19672, 46.23672, 46.27654, 46.31615, 46.35558, 46.3948, 46.43383, 
    46.47266, 46.51129, 46.54972, 46.58796, 46.626, 46.66383, 46.70147, 
    46.7389, 46.77613, 46.81316, 46.84999, 46.88661, 46.92303, 46.95925, 
    46.99526, 47.03106, 47.06666, 47.10205, 47.13724, 47.17221, 47.20699, 
    47.24155, 47.2759, 47.31004, 47.34397, 47.37769, 47.4112, 47.4445, 
    47.47758, 47.51046, 47.54312, 47.57556, 47.6078, 47.63981, 47.67161, 
    47.7032, 47.73457, 47.76572, 47.79665, 47.82737, 47.85787, 47.88815, 
    47.91821, 47.94805, 47.97767, 48.00707, 48.03625, 48.0652, 48.09394, 
    48.12245, 48.15074, 48.17881, 48.20665, 48.23426, 48.26166, 48.28882, 
    48.31577, 48.34248, 48.36897, 48.39523, 48.42126, 48.44706, 48.47264, 
    48.49799, 48.52311, 48.54799, 48.57265, 48.59708, 48.62127, 48.64524, 
    48.66897, 48.69247, 48.71574, 48.73877, 48.76157, 48.78414, 48.80647, 
    48.82857, 48.85043, 48.87206, 48.89344, 48.9146, 48.93552, 48.9562, 
    48.97664, 48.99685, 49.01682, 49.03654, 49.05603, 49.07529, 49.0943, 
    49.11307, 49.1316, 49.14989, 49.16794, 49.18575, 49.20332, 49.22064, 
    49.23773, 49.25457, 49.27116, 49.28752, 49.30363, 49.3195, 49.33512, 
    49.3505, 49.36564, 49.38053, 49.39517, 49.40957, 49.42373, 49.43763, 
    49.45129, 49.46471, 49.47788, 49.4908, 49.50348, 49.5159, 49.52808, 
    49.54001, 49.5517, 49.56313, 49.57432, 49.58525, 49.59594, 49.60638, 
    49.61657, 49.62651, 49.6362, 49.64565, 49.65484, 49.66378, 49.67247, 
    49.68091, 49.68909, 49.69703, 49.70472, 49.71215, 49.71934, 49.72627, 
    49.73295, 49.73938, 49.74556, 49.75148, 49.75716, 49.76258, 49.76775, 
    49.77266, 49.77732, 49.78173, 49.78589, 49.7898, 49.79345, 49.79685, 
    49.8, 49.80289, 49.80553, 49.80792, 49.81005, 49.81193, 49.81356, 
    49.81493, 49.81605, 49.81692, 49.81753, 49.81789, 49.818, 49.81785, 
    49.81745, 49.8168, 49.81589, 49.81473, 49.81332, 49.81165, 49.80973, 
    49.80756, 49.80513, 49.80245, 49.79951, 49.79633, 49.79289, 49.7892, 
    49.78525, 49.78106, 49.7766, 49.7719, 49.76694, 49.76174, 49.75628, 
    49.75056, 49.7446, 49.73838, 49.73191, 49.72519, 49.71822, 49.71099, 
    49.70352, 49.69579, 49.68782, 49.67959, 49.67111, 49.66238, 49.6534, 
    49.64417, 49.63469, 49.62496, 49.61498, 49.60475, 49.59427, 49.58354, 
    49.57256, 49.56134, 49.54987, 49.53814, 49.52617, 49.51395, 49.50149, 
    49.48877, 49.47581, 49.4626, 49.44915, 49.43545, 49.4215, 49.40731, 
    49.39287, 49.37819, 49.36326, 49.34809, 49.33267, 49.31701, 49.3011, 
    49.28495, 49.26855, 49.25192, 49.23504, 49.21792, 49.20055, 49.18295, 
    49.1651, 49.14701, 49.12868, 49.11012, 49.0913, 49.07226, 49.05297, 
    49.03344, 49.01367, 48.99367, 48.97342, 48.95294, 48.93222, 48.91127, 
    48.89008, 48.86865, 48.84698, 48.82508, 48.80295, 48.78058, 48.75798, 
    48.73514, 48.71207, 48.68877, 48.66523, 48.64146, 48.61746, 48.59323, 
    48.56876, 48.54407, 48.51915, 48.49399, 48.46861, 48.443, 48.41716, 
    48.39109, 48.36479, 48.33827, 48.31152, 48.28454, 48.25734, 48.22991, 
    48.20226, 48.17438, 48.14628, 48.11796, 48.08941, 48.06064, 48.03165, 
    48.00243, 47.973, 47.94334, 47.91347, 47.88337, 47.85306, 47.82253, 
    47.79177, 47.7608, 47.72962, 47.69822, 47.6666, 47.63476, 47.60271, 
    47.57045, 47.53796, 47.50527, 47.47237, 47.43925, 47.40591, 47.37237, 
    47.33862, 47.30465, 47.27048, 47.23609, 47.2015, 47.1667, 47.13169, 
    47.09647, 47.06104, 47.02541, 46.98957, 46.95353, 46.91729, 46.88083, 
    46.84418, 46.80732, 46.77026, 46.73299, 46.69553, 46.65786, 46.61999, 
    46.58192, 46.54366, 46.50519, 46.46653, 46.42767, 46.38861, 46.34935, 
    46.3099, 46.27025,
  41.90884, 41.96431, 42.01963, 42.07481, 42.12984, 42.18473, 42.23948, 
    42.29407, 42.34852, 42.40282, 42.45697, 42.51097, 42.56482, 42.61852, 
    42.67207, 42.72548, 42.77872, 42.83182, 42.88476, 42.93755, 42.99018, 
    43.04267, 43.09499, 43.14716, 43.19918, 43.25103, 43.30273, 43.35427, 
    43.40566, 43.45688, 43.50795, 43.55885, 43.6096, 43.66018, 43.71061, 
    43.76086, 43.81096, 43.86089, 43.91066, 43.96027, 44.00971, 44.05898, 
    44.10809, 44.15703, 44.20581, 44.25441, 44.30285, 44.35112, 44.39922, 
    44.44715, 44.49491, 44.5425, 44.58991, 44.63715, 44.68422, 44.73112, 
    44.77784, 44.82439, 44.87077, 44.91696, 44.96298, 45.00883, 45.0545, 
    45.09998, 45.14529, 45.19043, 45.23538, 45.28015, 45.32474, 45.36915, 
    45.41338, 45.45742, 45.50129, 45.54496, 45.58846, 45.63176, 45.67489, 
    45.71783, 45.76058, 45.80314, 45.84552, 45.88771, 45.92971, 45.97152, 
    46.01314, 46.05457, 46.09581, 46.13686, 46.17772, 46.21838, 46.25885, 
    46.29913, 46.33921, 46.3791, 46.41879, 46.45829, 46.49759, 46.53669, 
    46.5756, 46.6143, 46.65281, 46.69112, 46.72923, 46.76714, 46.80485, 
    46.84236, 46.87966, 46.91676, 46.95366, 46.99036, 47.02685, 47.06314, 
    47.09922, 47.13509, 47.17076, 47.20623, 47.24148, 47.27653, 47.31137, 
    47.346, 47.38042, 47.41463, 47.44863, 47.48242, 47.516, 47.54936, 
    47.58251, 47.61545, 47.64818, 47.68069, 47.71299, 47.74507, 47.77694, 
    47.80859, 47.84002, 47.87123, 47.90224, 47.93301, 47.96358, 47.99392, 
    48.02404, 48.05395, 48.08363, 48.11309, 48.14233, 48.17135, 48.20014, 
    48.22871, 48.25706, 48.28519, 48.31309, 48.34076, 48.36821, 48.39544, 
    48.42244, 48.44921, 48.47575, 48.50207, 48.52815, 48.55401, 48.57964, 
    48.60505, 48.63022, 48.65516, 48.67987, 48.70435, 48.7286, 48.75261, 
    48.7764, 48.79995, 48.82327, 48.84635, 48.8692, 48.89182, 48.9142, 
    48.93634, 48.95825, 48.97993, 49.00137, 49.02256, 49.04353, 49.06425, 
    49.08474, 49.105, 49.12501, 49.14478, 49.16431, 49.18361, 49.20266, 
    49.22147, 49.24004, 49.25838, 49.27647, 49.29432, 49.31192, 49.32928, 
    49.34641, 49.36329, 49.37992, 49.39631, 49.41246, 49.42836, 49.44402, 
    49.45943, 49.47461, 49.48953, 49.50421, 49.51864, 49.53283, 49.54676, 
    49.56046, 49.5739, 49.5871, 49.60005, 49.61275, 49.62521, 49.63742, 
    49.64938, 49.66109, 49.67255, 49.68376, 49.69472, 49.70543, 49.7159, 
    49.72611, 49.73607, 49.74579, 49.75525, 49.76446, 49.77342, 49.78213, 
    49.79059, 49.7988, 49.80676, 49.81446, 49.82191, 49.82911, 49.83606, 
    49.84276, 49.8492, 49.85539, 49.86133, 49.86702, 49.87245, 49.87763, 
    49.88256, 49.88723, 49.89165, 49.89582, 49.89973, 49.90339, 49.9068, 
    49.90995, 49.91286, 49.9155, 49.91789, 49.92003, 49.92192, 49.92355, 
    49.92492, 49.92605, 49.92692, 49.92753, 49.92789, 49.928, 49.92785, 
    49.92745, 49.9268, 49.92589, 49.92472, 49.92331, 49.92163, 49.91971, 
    49.91753, 49.9151, 49.91241, 49.90947, 49.90628, 49.90283, 49.89913, 
    49.89518, 49.89097, 49.88651, 49.88179, 49.87683, 49.87161, 49.86613, 
    49.86041, 49.85443, 49.8482, 49.84171, 49.83498, 49.82799, 49.82075, 
    49.81326, 49.80551, 49.79752, 49.78927, 49.78077, 49.77202, 49.76302, 
    49.75377, 49.74427, 49.73452, 49.72451, 49.71426, 49.70375, 49.693, 
    49.682, 49.67075, 49.65925, 49.6475, 49.6355, 49.62326, 49.61076, 
    49.59802, 49.58503, 49.57179, 49.55831, 49.54457, 49.5306, 49.51637, 
    49.5019, 49.48718, 49.47222, 49.45702, 49.44156, 49.42587, 49.40992, 
    49.39373, 49.3773, 49.36063, 49.34372, 49.32656, 49.30915, 49.29151, 
    49.27362, 49.25549, 49.23713, 49.21851, 49.19966, 49.18057, 49.16124, 
    49.14167, 49.12186, 49.10181, 49.08152, 49.06099, 49.04023, 49.01923, 
    48.99799, 48.97651, 48.9548, 48.93285, 48.91067, 48.88825, 48.8656, 
    48.84271, 48.81959, 48.79624, 48.77265, 48.74883, 48.72478, 48.70049, 
    48.67598, 48.65123, 48.62625, 48.60104, 48.57561, 48.54994, 48.52404, 
    48.49792, 48.47157, 48.44498, 48.41818, 48.39114, 48.36388, 48.3364, 
    48.30869, 48.28075, 48.25259, 48.22421, 48.1956, 48.16677, 48.13772, 
    48.10844, 48.07895, 48.04923, 48.01929, 47.98914, 47.95876, 47.92816, 
    47.89735, 47.86631, 47.83506, 47.80359, 47.77191, 47.74001, 47.70789, 
    47.67556, 47.64302, 47.61026, 47.57728, 47.5441, 47.5107, 47.47709, 
    47.44326, 47.40923, 47.37499, 47.34053, 47.30587, 47.271, 47.23592, 
    47.20063, 47.16513, 47.12943, 47.09352, 47.05741, 47.02109, 46.98457, 
    46.94784, 46.91091, 46.87377, 46.83644, 46.7989, 46.76116, 46.72322, 
    46.68507, 46.64674, 46.6082, 46.56946, 46.53052, 46.49139, 46.45205, 
    46.41253, 46.3728,
  42.00376, 42.05931, 42.11472, 42.16998, 42.2251, 42.28008, 42.3349, 
    42.38958, 42.44411, 42.4985, 42.55273, 42.60682, 42.66076, 42.71454, 
    42.76817, 42.82166, 42.87499, 42.92817, 42.9812, 43.03407, 43.08679, 
    43.13935, 43.19176, 43.24402, 43.29612, 43.34806, 43.39985, 43.45147, 
    43.50294, 43.55424, 43.6054, 43.65638, 43.70721, 43.75788, 43.80838, 
    43.85873, 43.90891, 43.95893, 44.00878, 44.05847, 44.10799, 44.15735, 
    44.20654, 44.25556, 44.30442, 44.35311, 44.40163, 44.44998, 44.49817, 
    44.54618, 44.59402, 44.64169, 44.68919, 44.73651, 44.78366, 44.83064, 
    44.87745, 44.92408, 44.97053, 45.01681, 45.06292, 45.10884, 45.15459, 
    45.20016, 45.24555, 45.29076, 45.33579, 45.38065, 45.42532, 45.46981, 
    45.51411, 45.55824, 45.60218, 45.64594, 45.68951, 45.7329, 45.7761, 
    45.81912, 45.86195, 45.90459, 45.94705, 45.98932, 46.0314, 46.07329, 
    46.11499, 46.15649, 46.19781, 46.23894, 46.27987, 46.32061, 46.36116, 
    46.40151, 46.44167, 46.48164, 46.5214, 46.56097, 46.60035, 46.63953, 
    46.67851, 46.71729, 46.75587, 46.79426, 46.83244, 46.87042, 46.90821, 
    46.94579, 46.98317, 47.02034, 47.05731, 47.09408, 47.13064, 47.167, 
    47.20316, 47.2391, 47.27484, 47.31038, 47.3457, 47.38082, 47.41573, 
    47.45043, 47.48492, 47.5192, 47.55326, 47.58712, 47.62077, 47.6542, 
    47.68742, 47.72043, 47.75322, 47.7858, 47.81816, 47.85031, 47.88224, 
    47.91396, 47.94545, 47.97673, 48.0078, 48.03864, 48.06927, 48.09967, 
    48.12986, 48.15982, 48.18957, 48.21909, 48.24839, 48.27747, 48.30633, 
    48.33496, 48.36337, 48.39155, 48.41951, 48.44725, 48.47475, 48.50204, 
    48.52909, 48.55592, 48.58252, 48.60889, 48.63504, 48.66095, 48.68664, 
    48.71209, 48.73732, 48.76231, 48.78708, 48.81161, 48.83591, 48.85998, 
    48.88382, 48.90742, 48.93079, 48.95392, 48.97682, 48.99949, 49.02192, 
    49.04411, 49.06607, 49.08779, 49.10927, 49.13052, 49.15153, 49.1723, 
    49.19284, 49.21313, 49.23319, 49.25301, 49.27258, 49.29192, 49.31101, 
    49.32987, 49.34848, 49.36686, 49.38499, 49.40287, 49.42052, 49.43792, 
    49.45508, 49.472, 49.48867, 49.5051, 49.52128, 49.53722, 49.55292, 
    49.56837, 49.58357, 49.59853, 49.61324, 49.6277, 49.64192, 49.65589, 
    49.66961, 49.68309, 49.69632, 49.7093, 49.72203, 49.73452, 49.74675, 
    49.75874, 49.77047, 49.78196, 49.7932, 49.80418, 49.81492, 49.82541, 
    49.83565, 49.84563, 49.85537, 49.86485, 49.87408, 49.88307, 49.8918, 
    49.90028, 49.9085, 49.91648, 49.9242, 49.93167, 49.93888, 49.94585, 
    49.95256, 49.95902, 49.96523, 49.97118, 49.97688, 49.98232, 49.98751, 
    49.99245, 49.99714, 50.00157, 50.00574, 50.00967, 50.01334, 50.01675, 
    50.01991, 50.02282, 50.02547, 50.02787, 50.03001, 50.0319, 50.03354, 
    50.03492, 50.03604, 50.03691, 50.03753, 50.03789, 50.038, 50.03785, 
    50.03745, 50.03679, 50.03588, 50.03472, 50.03329, 50.03162, 50.02969, 
    50.02751, 50.02507, 50.02238, 50.01943, 50.01623, 50.01278, 50.00906, 
    50.0051, 50.00089, 49.99641, 49.99169, 49.98671, 49.98148, 49.97599, 
    49.97025, 49.96426, 49.95802, 49.95152, 49.94476, 49.93776, 49.9305, 
    49.92299, 49.91523, 49.90722, 49.89895, 49.89043, 49.88166, 49.87264, 
    49.86337, 49.85384, 49.84407, 49.83405, 49.82377, 49.81324, 49.80246, 
    49.79144, 49.78016, 49.76863, 49.75686, 49.74483, 49.73256, 49.72003, 
    49.70726, 49.69424, 49.68098, 49.66746, 49.6537, 49.63969, 49.62543, 
    49.61093, 49.59618, 49.58118, 49.56594, 49.55045, 49.53472, 49.51874, 
    49.50252, 49.48605, 49.46934, 49.45238, 49.43518, 49.41774, 49.40006, 
    49.38213, 49.36396, 49.34555, 49.3269, 49.30801, 49.28888, 49.2695, 
    49.24989, 49.23003, 49.20994, 49.18961, 49.16903, 49.14822, 49.12717, 
    49.10589, 49.08437, 49.06261, 49.04062, 49.01838, 48.99591, 48.97321, 
    48.95028, 48.9271, 48.9037, 48.88006, 48.85619, 48.83208, 48.80775, 
    48.78318, 48.75838, 48.73335, 48.70808, 48.68259, 48.65687, 48.63092, 
    48.60474, 48.57833, 48.55169, 48.52483, 48.49773, 48.47042, 48.44287, 
    48.4151, 48.38711, 48.35889, 48.33044, 48.30178, 48.27289, 48.24377, 
    48.21444, 48.18488, 48.1551, 48.1251, 48.09488, 48.06444, 48.03378, 
    48.0029, 47.9718, 47.94049, 47.90895, 47.8772, 47.84524, 47.81306, 
    47.78066, 47.74805, 47.71522, 47.68218, 47.64893, 47.61546, 47.58178, 
    47.54789, 47.51379, 47.47947, 47.44495, 47.41022, 47.37528, 47.34013, 
    47.30477, 47.2692, 47.23343, 47.19745, 47.16126, 47.12487, 47.08828, 
    47.05148, 47.01447, 46.97726, 46.93985, 46.90224, 46.86443, 46.82642, 
    46.7882, 46.74978, 46.71117, 46.67236, 46.63335, 46.59414, 46.55473, 
    46.51513, 46.47533,
  42.09863, 42.15427, 42.20976, 42.26511, 42.32031, 42.37537, 42.43028, 
    42.48504, 42.53966, 42.59413, 42.64845, 42.70262, 42.75664, 42.81051, 
    42.86423, 42.9178, 42.97121, 43.02448, 43.07759, 43.13055, 43.18335, 
    43.236, 43.28849, 43.34084, 43.39302, 43.44504, 43.49691, 43.54862, 
    43.60017, 43.65157, 43.7028, 43.75387, 43.80478, 43.85553, 43.90612, 
    43.95655, 44.00681, 44.05692, 44.10685, 44.15662, 44.20623, 44.25567, 
    44.30495, 44.35405, 44.40299, 44.45177, 44.50037, 44.54881, 44.59707, 
    44.64516, 44.69309, 44.74084, 44.78842, 44.83583, 44.88306, 44.93013, 
    44.97701, 45.02372, 45.07026, 45.11662, 45.16281, 45.20882, 45.25464, 
    45.3003, 45.34577, 45.39106, 45.43618, 45.48111, 45.52586, 45.57043, 
    45.61482, 45.65902, 45.70304, 45.74688, 45.79053, 45.834, 45.87729, 
    45.92038, 45.96329, 46.00602, 46.04855, 46.0909, 46.13305, 46.17502, 
    46.2168, 46.25838, 46.29978, 46.34098, 46.38199, 46.42281, 46.46344, 
    46.50386, 46.5441, 46.58414, 46.62399, 46.66363, 46.70308, 46.74234, 
    46.78139, 46.82025, 46.85891, 46.89737, 46.93562, 46.97368, 47.01154, 
    47.04919, 47.08664, 47.12389, 47.16093, 47.19777, 47.23441, 47.27084, 
    47.30706, 47.34308, 47.37889, 47.4145, 47.4499, 47.48508, 47.52006, 
    47.55483, 47.58939, 47.62374, 47.65788, 47.6918, 47.72552, 47.75902, 
    47.7923, 47.82538, 47.85824, 47.89088, 47.92332, 47.95553, 47.98753, 
    48.01931, 48.05087, 48.08222, 48.11334, 48.14425, 48.17494, 48.20541, 
    48.23566, 48.26569, 48.29549, 48.32508, 48.35444, 48.38358, 48.4125, 
    48.44119, 48.46966, 48.4979, 48.52592, 48.55371, 48.58128, 48.60862, 
    48.63573, 48.66262, 48.68927, 48.71571, 48.74191, 48.76788, 48.79362, 
    48.81913, 48.84441, 48.86946, 48.89428, 48.91886, 48.94321, 48.96733, 
    48.99122, 49.01487, 49.0383, 49.06148, 49.08443, 49.10714, 49.12962, 
    49.15187, 49.17387, 49.19564, 49.21717, 49.23847, 49.25953, 49.28034, 
    49.30092, 49.32126, 49.34136, 49.36122, 49.38084, 49.40022, 49.41936, 
    49.43826, 49.45691, 49.47533, 49.4935, 49.51143, 49.52911, 49.54655, 
    49.56375, 49.58071, 49.59742, 49.61388, 49.6301, 49.64608, 49.66181, 
    49.67729, 49.69253, 49.70752, 49.72226, 49.73676, 49.75101, 49.76501, 
    49.77877, 49.79227, 49.80553, 49.81854, 49.8313, 49.84381, 49.85608, 
    49.86809, 49.87986, 49.89137, 49.90263, 49.91365, 49.92441, 49.93492, 
    49.94518, 49.95519, 49.96495, 49.97445, 49.98371, 49.99271, 50.00146, 
    50.00996, 50.0182, 50.0262, 50.03394, 50.04142, 50.04866, 50.05563, 
    50.06236, 50.06884, 50.07505, 50.08102, 50.08673, 50.09219, 50.0974, 
    50.10235, 50.10704, 50.11148, 50.11567, 50.1196, 50.12328, 50.12671, 
    50.12987, 50.13279, 50.13544, 50.13785, 50.14, 50.14189, 50.14353, 
    50.14491, 50.14604, 50.14691, 50.14753, 50.14789, 50.148, 50.14785, 
    50.14745, 50.14679, 50.14588, 50.14471, 50.14328, 50.14161, 50.13967, 
    50.13748, 50.13504, 50.13234, 50.12939, 50.12618, 50.12271, 50.119, 
    50.11502, 50.1108, 50.10632, 50.10158, 50.09659, 50.09135, 50.08585, 
    50.08009, 50.07409, 50.06783, 50.06131, 50.05455, 50.04753, 50.04025, 
    50.03273, 50.02495, 50.01691, 50.00863, 50.00009, 49.9913, 49.98226, 
    49.97297, 49.96342, 49.95362, 49.94357, 49.93327, 49.92272, 49.91192, 
    49.90087, 49.88956, 49.87801, 49.86621, 49.85416, 49.84185, 49.8293, 
    49.8165, 49.80345, 49.79015, 49.77661, 49.76281, 49.74877, 49.73449, 
    49.71995, 49.70516, 49.69013, 49.67486, 49.65934, 49.64357, 49.62755, 
    49.61129, 49.59479, 49.57804, 49.56105, 49.54381, 49.52633, 49.50861, 
    49.49064, 49.47243, 49.45398, 49.43528, 49.41635, 49.39717, 49.37775, 
    49.3581, 49.3382, 49.31806, 49.29768, 49.27707, 49.25621, 49.23512, 
    49.21378, 49.19221, 49.17041, 49.14836, 49.12608, 49.10357, 49.08081, 
    49.05783, 49.03461, 49.01115, 48.98746, 48.96354, 48.93938, 48.91499, 
    48.89037, 48.86551, 48.84042, 48.81511, 48.78956, 48.76378, 48.73778, 
    48.71154, 48.68507, 48.65838, 48.63146, 48.60431, 48.57693, 48.54933, 
    48.5215, 48.49345, 48.46517, 48.43666, 48.40794, 48.37899, 48.34981, 
    48.32041, 48.29079, 48.26095, 48.23089, 48.2006, 48.1701, 48.13938, 
    48.10843, 48.07727, 48.04589, 48.01429, 47.98248, 47.95045, 47.9182, 
    47.88573, 47.85306, 47.82016, 47.78706, 47.75373, 47.7202, 47.68645, 
    47.65249, 47.61832, 47.58394, 47.54935, 47.51455, 47.47953, 47.44431, 
    47.40888, 47.37325, 47.3374, 47.30135, 47.26509, 47.22863, 47.19196, 
    47.15509, 47.11801, 47.08073, 47.04325, 47.00556, 46.96767, 46.92958, 
    46.8913, 46.85281, 46.81412, 46.77523, 46.73614, 46.69686, 46.65738, 
    46.61769, 46.57782,
  42.19345, 42.24918, 42.30475, 42.36018, 42.41547, 42.47062, 42.52561, 
    42.58046, 42.63516, 42.68971, 42.74412, 42.79837, 42.85248, 42.90643, 
    42.96024, 43.01389, 43.06739, 43.12074, 43.17393, 43.22698, 43.27987, 
    43.3326, 43.38518, 43.4376, 43.48987, 43.54198, 43.59393, 43.64573, 
    43.69736, 43.74884, 43.80016, 43.85131, 43.90231, 43.95314, 44.00382, 
    44.05433, 44.10468, 44.15486, 44.20488, 44.25474, 44.30443, 44.35395, 
    44.40331, 44.4525, 44.50153, 44.55038, 44.59907, 44.64759, 44.69593, 
    44.74411, 44.79212, 44.83995, 44.88762, 44.93511, 44.98243, 45.02957, 
    45.07654, 45.12334, 45.16995, 45.2164, 45.26266, 45.30875, 45.35466, 
    45.4004, 45.44595, 45.49133, 45.53652, 45.58154, 45.62637, 45.67102, 
    45.71548, 45.75977, 45.80387, 45.84779, 45.89153, 45.93507, 45.97844, 
    46.02161, 46.0646, 46.1074, 46.15002, 46.19244, 46.23468, 46.27672, 
    46.31858, 46.36024, 46.40171, 46.443, 46.48409, 46.52498, 46.56568, 
    46.60619, 46.6465, 46.68662, 46.72654, 46.76626, 46.80579, 46.84512, 
    46.88425, 46.92318, 46.96191, 47.00045, 47.03878, 47.07691, 47.11484, 
    47.15257, 47.19009, 47.22741, 47.26453, 47.30145, 47.33815, 47.37466, 
    47.41095, 47.44704, 47.48293, 47.5186, 47.55407, 47.58932, 47.62437, 
    47.65921, 47.69384, 47.72826, 47.76247, 47.79646, 47.83025, 47.86382, 
    47.89717, 47.93031, 47.96324, 47.99595, 48.02845, 48.06073, 48.09279, 
    48.12464, 48.15627, 48.18768, 48.21887, 48.24984, 48.28059, 48.31113, 
    48.34144, 48.37153, 48.4014, 48.43105, 48.46047, 48.48967, 48.51865, 
    48.5474, 48.57593, 48.60424, 48.63231, 48.66016, 48.68779, 48.71519, 
    48.74236, 48.7693, 48.79602, 48.8225, 48.84876, 48.87479, 48.90059, 
    48.92615, 48.95148, 48.97659, 49.00146, 49.0261, 49.0505, 49.07468, 
    49.09862, 49.12232, 49.14579, 49.16903, 49.19203, 49.21479, 49.23732, 
    49.25961, 49.28167, 49.30349, 49.32507, 49.34641, 49.36751, 49.38837, 
    49.409, 49.42938, 49.44953, 49.46943, 49.4891, 49.50852, 49.5277, 
    49.54664, 49.56534, 49.58379, 49.60201, 49.61997, 49.6377, 49.65518, 
    49.67242, 49.68941, 49.70615, 49.72266, 49.73891, 49.75492, 49.77069, 
    49.78621, 49.80148, 49.81651, 49.83128, 49.84581, 49.8601, 49.87413, 
    49.88792, 49.90145, 49.91475, 49.92778, 49.94057, 49.95311, 49.9654, 
    49.97745, 49.98924, 50.00078, 50.01207, 50.02311, 50.03389, 50.04443, 
    50.05471, 50.06474, 50.07452, 50.08405, 50.09333, 50.10235, 50.11112, 
    50.11964, 50.1279, 50.13591, 50.14367, 50.15117, 50.15842, 50.16542, 
    50.17216, 50.17865, 50.18489, 50.19087, 50.19659, 50.20206, 50.20728, 
    50.21224, 50.21695, 50.2214, 50.2256, 50.22954, 50.23322, 50.23665, 
    50.23983, 50.24275, 50.24541, 50.24782, 50.24998, 50.25187, 50.25352, 
    50.2549, 50.25603, 50.25691, 50.25753, 50.25789, 50.258, 50.25785, 
    50.25745, 50.25679, 50.25587, 50.2547, 50.25327, 50.25159, 50.24965, 
    50.24746, 50.24501, 50.24231, 50.23935, 50.23613, 50.23266, 50.22893, 
    50.22495, 50.22071, 50.21622, 50.21147, 50.20647, 50.20121, 50.1957, 
    50.18994, 50.18392, 50.17764, 50.17111, 50.16433, 50.1573, 50.15001, 
    50.14246, 50.13466, 50.12661, 50.11831, 50.10975, 50.10094, 50.09188, 
    50.08256, 50.07299, 50.06317, 50.0531, 50.04278, 50.0322, 50.02137, 
    50.0103, 49.99897, 49.98739, 49.97556, 49.96348, 49.95115, 49.93857, 
    49.92574, 49.91266, 49.89933, 49.88575, 49.87193, 49.85786, 49.84353, 
    49.82896, 49.81415, 49.79908, 49.78377, 49.76822, 49.75241, 49.73636, 
    49.72006, 49.70352, 49.68674, 49.6697, 49.65243, 49.63491, 49.61715, 
    49.59914, 49.58089, 49.5624, 49.54366, 49.52468, 49.50546, 49.486, 
    49.4663, 49.44636, 49.42617, 49.40575, 49.38509, 49.36419, 49.34304, 
    49.32167, 49.30005, 49.27819, 49.2561, 49.23377, 49.21121, 49.1884, 
    49.16537, 49.14209, 49.11859, 49.09484, 49.07087, 49.04666, 49.02222, 
    48.99754, 48.97263, 48.94749, 48.92212, 48.89652, 48.87069, 48.84462, 
    48.81833, 48.79181, 48.76506, 48.73808, 48.71087, 48.68344, 48.65577, 
    48.62789, 48.59977, 48.57143, 48.54287, 48.51408, 48.48507, 48.45583, 
    48.42637, 48.39669, 48.36679, 48.33666, 48.30631, 48.27575, 48.24496, 
    48.21395, 48.18272, 48.15128, 48.11962, 48.08773, 48.05564, 48.02332, 
    47.99079, 47.95805, 47.92508, 47.89191, 47.85852, 47.82492, 47.7911, 
    47.75707, 47.72283, 47.68838, 47.65372, 47.61885, 47.58376, 47.54847, 
    47.51297, 47.47726, 47.44135, 47.40522, 47.3689, 47.33236, 47.29562, 
    47.25867, 47.22152, 47.18417, 47.14661, 47.10885, 47.07089, 47.03273, 
    46.99437, 46.9558, 46.91704, 46.87807, 46.83891, 46.79955, 46.75999, 
    46.72024, 46.68028,
  42.28823, 42.34403, 42.3997, 42.45521, 42.51059, 42.56581, 42.62089, 
    42.67583, 42.73061, 42.78525, 42.83974, 42.89408, 42.94827, 43.00231, 
    43.0562, 43.10994, 43.16352, 43.21696, 43.27024, 43.32336, 43.37634, 
    43.42915, 43.48182, 43.53432, 43.58668, 43.63887, 43.69091, 43.74279, 
    43.79451, 43.84607, 43.89747, 43.94872, 43.99979, 44.05071, 44.10147, 
    44.15207, 44.2025, 44.25277, 44.30287, 44.35281, 44.40258, 44.45219, 
    44.50164, 44.55091, 44.60002, 44.64896, 44.69773, 44.74633, 44.79476, 
    44.84302, 44.89111, 44.93903, 44.98678, 45.03435, 45.08175, 45.12898, 
    45.17603, 45.22291, 45.26961, 45.31613, 45.36248, 45.40865, 45.45465, 
    45.50046, 45.5461, 45.59155, 45.63683, 45.68192, 45.72684, 45.77157, 
    45.81612, 45.86049, 45.90467, 45.94867, 45.99248, 46.03611, 46.07955, 
    46.12281, 46.16587, 46.20876, 46.25145, 46.29395, 46.33627, 46.37839, 
    46.42033, 46.46207, 46.50362, 46.54498, 46.58614, 46.62712, 46.6679, 
    46.70848, 46.74887, 46.78906, 46.82906, 46.86886, 46.90847, 46.94787, 
    46.98708, 47.02608, 47.06489, 47.1035, 47.14191, 47.18011, 47.21812, 
    47.25592, 47.29352, 47.33091, 47.3681, 47.40509, 47.44187, 47.47845, 
    47.51482, 47.55098, 47.58693, 47.62268, 47.65822, 47.69355, 47.72866, 
    47.76358, 47.79827, 47.83276, 47.86704, 47.9011, 47.93495, 47.96859, 
    48.00201, 48.03522, 48.06822, 48.101, 48.13356, 48.16591, 48.19804, 
    48.22995, 48.26165, 48.29312, 48.32438, 48.35542, 48.38623, 48.41683, 
    48.4472, 48.47736, 48.50729, 48.537, 48.56649, 48.59575, 48.62479, 
    48.6536, 48.68219, 48.71055, 48.73869, 48.7666, 48.79429, 48.82174, 
    48.84897, 48.87597, 48.90274, 48.92929, 48.9556, 48.98169, 49.00754, 
    49.03316, 49.05855, 49.08371, 49.10863, 49.13332, 49.15778, 49.18201, 
    49.206, 49.22976, 49.25328, 49.27657, 49.29961, 49.32243, 49.34501, 
    49.36735, 49.38945, 49.41132, 49.43295, 49.45433, 49.47548, 49.4964, 
    49.51707, 49.53749, 49.55769, 49.57763, 49.59734, 49.61681, 49.63603, 
    49.65501, 49.67375, 49.69225, 49.7105, 49.72851, 49.74628, 49.7638, 
    49.78107, 49.7981, 49.81489, 49.83143, 49.84772, 49.86377, 49.87957, 
    49.89513, 49.91043, 49.92549, 49.9403, 49.95486, 49.96918, 49.98325, 
    49.99707, 50.01063, 50.02395, 50.03702, 50.04984, 50.06241, 50.07473, 
    50.0868, 50.09861, 50.11018, 50.1215, 50.13256, 50.14337, 50.15393, 
    50.16424, 50.17429, 50.1841, 50.19365, 50.20295, 50.21199, 50.22078, 
    50.22932, 50.2376, 50.24563, 50.2534, 50.26093, 50.26819, 50.27521, 
    50.28196, 50.28847, 50.29472, 50.30071, 50.30645, 50.31193, 50.31716, 
    50.32214, 50.32685, 50.33131, 50.33552, 50.33947, 50.34317, 50.3466, 
    50.34979, 50.35271, 50.35538, 50.3578, 50.35996, 50.36186, 50.36351, 
    50.36489, 50.36603, 50.36691, 50.36753, 50.36789, 50.368, 50.36785, 
    50.36745, 50.36678, 50.36587, 50.36469, 50.36326, 50.36158, 50.35963, 
    50.35743, 50.35498, 50.35227, 50.3493, 50.34608, 50.3426, 50.33886, 
    50.33487, 50.33062, 50.32612, 50.32137, 50.31635, 50.31108, 50.30556, 
    50.29978, 50.29374, 50.28746, 50.28091, 50.27411, 50.26706, 50.25975, 
    50.25219, 50.24437, 50.23631, 50.22798, 50.21941, 50.21058, 50.20149, 
    50.19215, 50.18256, 50.17272, 50.16262, 50.15228, 50.14168, 50.13083, 
    50.11972, 50.10837, 50.09676, 50.0849, 50.0728, 50.06044, 50.04783, 
    50.03497, 50.02186, 50.0085, 49.9949, 49.98104, 49.96693, 49.95258, 
    49.93798, 49.92313, 49.90803, 49.89268, 49.87709, 49.86125, 49.84516, 
    49.82883, 49.81225, 49.79543, 49.77835, 49.76104, 49.74348, 49.72568, 
    49.70763, 49.68934, 49.67081, 49.65203, 49.63301, 49.61375, 49.59424, 
    49.57449, 49.55451, 49.53428, 49.51381, 49.4931, 49.47215, 49.45097, 
    49.42954, 49.40788, 49.38597, 49.36383, 49.34145, 49.31884, 49.29599, 
    49.2729, 49.24957, 49.22601, 49.20222, 49.17819, 49.15393, 49.12943, 
    49.1047, 49.07974, 49.05455, 49.02912, 49.00346, 48.97757, 48.95145, 
    48.92511, 48.89853, 48.87172, 48.84468, 48.81742, 48.78992, 48.7622, 
    48.73426, 48.70608, 48.67768, 48.64906, 48.62021, 48.59113, 48.56184, 
    48.53231, 48.50257, 48.4726, 48.44241, 48.412, 48.38137, 48.35052, 
    48.31945, 48.28815, 48.25665, 48.22492, 48.19297, 48.1608, 48.12843, 
    48.09583, 48.06301, 48.02999, 47.99674, 47.96328, 47.92961, 47.89573, 
    47.86163, 47.82732, 47.7928, 47.75807, 47.72313, 47.68797, 47.65261, 
    47.61704, 47.58126, 47.54527, 47.50908, 47.47268, 47.43607, 47.39925, 
    47.36223, 47.32501, 47.28758, 47.24995, 47.21212, 47.17408, 47.13585, 
    47.09741, 47.05877, 47.01993, 46.98089, 46.94165, 46.90221, 46.86258, 
    46.82275, 46.78272,
  42.38295, 42.43884, 42.49459, 42.55019, 42.60565, 42.66096, 42.71613, 
    42.77114, 42.82602, 42.88074, 42.93531, 42.98974, 43.04401, 43.09814, 
    43.15211, 43.20593, 43.25961, 43.31313, 43.36649, 43.4197, 43.47276, 
    43.52567, 43.57841, 43.631, 43.68344, 43.73572, 43.78784, 43.83981, 
    43.89161, 43.94326, 43.99474, 44.04607, 44.09724, 44.14824, 44.19908, 
    44.24976, 44.30028, 44.35063, 44.40082, 44.45084, 44.5007, 44.55039, 
    44.59992, 44.64928, 44.69847, 44.74749, 44.79635, 44.84503, 44.89355, 
    44.94189, 44.99006, 45.03807, 45.0859, 45.13355, 45.18103, 45.22834, 
    45.27548, 45.32244, 45.36922, 45.41583, 45.46226, 45.50851, 45.55459, 
    45.60049, 45.64621, 45.69174, 45.7371, 45.78228, 45.82727, 45.87209, 
    45.91672, 45.96116, 46.00543, 46.04951, 46.0934, 46.13711, 46.18063, 
    46.22397, 46.26712, 46.31008, 46.35285, 46.39543, 46.43782, 46.48003, 
    46.52204, 46.56386, 46.60549, 46.64693, 46.68818, 46.72923, 46.77008, 
    46.81075, 46.85121, 46.89148, 46.93156, 46.97143, 47.01111, 47.05059, 
    47.08987, 47.12896, 47.16784, 47.20652, 47.24501, 47.28329, 47.32137, 
    47.35924, 47.39692, 47.43438, 47.47165, 47.50871, 47.54556, 47.58221, 
    47.61865, 47.65488, 47.69091, 47.72673, 47.76234, 47.79774, 47.83293, 
    47.86791, 47.90268, 47.93724, 47.97158, 48.00572, 48.03964, 48.07335, 
    48.10684, 48.14011, 48.17318, 48.20602, 48.23866, 48.27107, 48.30326, 
    48.33524, 48.367, 48.39854, 48.42987, 48.46097, 48.49185, 48.52251, 
    48.55295, 48.58317, 48.61316, 48.64293, 48.67248, 48.70181, 48.73091, 
    48.75978, 48.78843, 48.81686, 48.84505, 48.87302, 48.90077, 48.92828, 
    48.95557, 48.98263, 49.00946, 49.03606, 49.06243, 49.08857, 49.11448, 
    49.14015, 49.1656, 49.19081, 49.21579, 49.24054, 49.26505, 49.28933, 
    49.31337, 49.33718, 49.36076, 49.38409, 49.40719, 49.43006, 49.45269, 
    49.47507, 49.49723, 49.51914, 49.54082, 49.56225, 49.58345, 49.60441, 
    49.62513, 49.6456, 49.66584, 49.68583, 49.70558, 49.72509, 49.74436, 
    49.76338, 49.78216, 49.8007, 49.81899, 49.83704, 49.85485, 49.87241, 
    49.88972, 49.90679, 49.92362, 49.94019, 49.95652, 49.97261, 49.98845, 
    50.00404, 50.01937, 50.03447, 50.04932, 50.06391, 50.07826, 50.09236, 
    50.10621, 50.11981, 50.13316, 50.14626, 50.1591, 50.1717, 50.18405, 
    50.19614, 50.20799, 50.21959, 50.23093, 50.24201, 50.25285, 50.26344, 
    50.27377, 50.28384, 50.29367, 50.30324, 50.31256, 50.32162, 50.33044, 
    50.33899, 50.34729, 50.35534, 50.36314, 50.37068, 50.37796, 50.38499, 
    50.39176, 50.39828, 50.40454, 50.41055, 50.41631, 50.4218, 50.42704, 
    50.43203, 50.43676, 50.44123, 50.44545, 50.44941, 50.45311, 50.45655, 
    50.45974, 50.46268, 50.46535, 50.46778, 50.46994, 50.47185, 50.4735, 
    50.47489, 50.47602, 50.4769, 50.47753, 50.47789, 50.478, 50.47785, 
    50.47744, 50.47678, 50.47586, 50.47469, 50.47325, 50.47156, 50.46962, 
    50.46741, 50.46495, 50.46223, 50.45926, 50.45603, 50.45254, 50.4488, 
    50.44479, 50.44054, 50.43602, 50.43126, 50.42623, 50.42095, 50.41541, 
    50.40962, 50.40357, 50.39727, 50.39071, 50.3839, 50.37682, 50.3695, 
    50.36192, 50.35409, 50.346, 50.33766, 50.32906, 50.32021, 50.3111, 
    50.30175, 50.29213, 50.28227, 50.27215, 50.26178, 50.25115, 50.24028, 
    50.22915, 50.21777, 50.20613, 50.19425, 50.18211, 50.16973, 50.15709, 
    50.1442, 50.13106, 50.11767, 50.10403, 50.09015, 50.07601, 50.06162, 
    50.04698, 50.0321, 50.01696, 50.00158, 49.98596, 49.97008, 49.95396, 
    49.93759, 49.92097, 49.90411, 49.887, 49.86965, 49.85205, 49.83421, 
    49.81612, 49.79778, 49.77921, 49.76039, 49.74133, 49.72202, 49.70247, 
    49.68268, 49.66265, 49.64238, 49.62186, 49.60111, 49.58011, 49.55888, 
    49.5374, 49.51569, 49.49374, 49.47155, 49.44912, 49.42646, 49.40355, 
    49.38042, 49.35704, 49.33343, 49.30959, 49.2855, 49.26119, 49.23664, 
    49.21185, 49.18684, 49.16159, 49.13611, 49.11039, 49.08445, 49.05827, 
    49.03187, 49.00523, 48.97837, 48.95127, 48.92395, 48.89639, 48.86861, 
    48.84061, 48.81237, 48.78392, 48.75523, 48.72632, 48.69718, 48.66782, 
    48.63824, 48.60843, 48.5784, 48.54815, 48.51767, 48.48698, 48.45606, 
    48.42493, 48.39357, 48.36199, 48.3302, 48.29819, 48.26596, 48.23351, 
    48.20084, 48.16796, 48.13486, 48.10155, 48.06803, 48.03429, 48.00033, 
    47.96617, 47.93179, 47.89719, 47.86239, 47.82738, 47.79216, 47.75672, 
    47.72108, 47.68523, 47.64917, 47.6129, 47.57643, 47.53975, 47.50286, 
    47.46577, 47.42847, 47.39097, 47.35326, 47.31536, 47.27724, 47.23893, 
    47.20042, 47.16171, 47.12279, 47.08368, 47.04436, 47.00485, 46.96514, 
    46.92523, 46.88512,
  42.47763, 42.5336, 42.58944, 42.64512, 42.70066, 42.75606, 42.81131, 
    42.86641, 42.92137, 42.97618, 43.03084, 43.08535, 43.13971, 43.19392, 
    43.24798, 43.30188, 43.35564, 43.40924, 43.4627, 43.516, 43.56914, 
    43.62212, 43.67496, 43.72763, 43.78016, 43.83252, 43.88473, 43.93678, 
    43.98867, 44.0404, 44.09197, 44.14338, 44.19463, 44.24572, 44.29665, 
    44.34741, 44.39801, 44.44845, 44.49872, 44.54883, 44.59877, 44.64855, 
    44.69816, 44.7476, 44.79688, 44.84599, 44.89492, 44.94369, 44.99229, 
    45.04072, 45.08898, 45.13706, 45.18497, 45.23272, 45.28028, 45.32767, 
    45.37489, 45.42193, 45.4688, 45.51549, 45.562, 45.60834, 45.6545, 
    45.70048, 45.74628, 45.7919, 45.83734, 45.8826, 45.92767, 45.97256, 
    46.01728, 46.06181, 46.10615, 46.15031, 46.19429, 46.23808, 46.28168, 
    46.32509, 46.36832, 46.41136, 46.45422, 46.49688, 46.53935, 46.58163, 
    46.62373, 46.66563, 46.70734, 46.74885, 46.79017, 46.8313, 46.87223, 
    46.91298, 46.95352, 46.99387, 47.03402, 47.07397, 47.11373, 47.15329, 
    47.19265, 47.2318, 47.27076, 47.30952, 47.34808, 47.38644, 47.42459, 
    47.46254, 47.50029, 47.53783, 47.57517, 47.6123, 47.64923, 47.68595, 
    47.72246, 47.75877, 47.79487, 47.83076, 47.86644, 47.90191, 47.93718, 
    47.97223, 48.00706, 48.04169, 48.07611, 48.11031, 48.1443, 48.17808, 
    48.21164, 48.24498, 48.27811, 48.31103, 48.34373, 48.37621, 48.40847, 
    48.44051, 48.47234, 48.50395, 48.53534, 48.5665, 48.59745, 48.62817, 
    48.65868, 48.68896, 48.71902, 48.74885, 48.77846, 48.80785, 48.83701, 
    48.86595, 48.89466, 48.92314, 48.9514, 48.97943, 49.00723, 49.03481, 
    49.06215, 49.08927, 49.11616, 49.14281, 49.16924, 49.19544, 49.22141, 
    49.24714, 49.27264, 49.2979, 49.32294, 49.34774, 49.3723, 49.39664, 
    49.42073, 49.44459, 49.46822, 49.49161, 49.51476, 49.53767, 49.56035, 
    49.58279, 49.605, 49.62696, 49.64868, 49.67016, 49.69141, 49.71241, 
    49.73317, 49.7537, 49.77398, 49.79401, 49.81381, 49.83336, 49.85268, 
    49.87174, 49.89056, 49.90915, 49.92748, 49.94557, 49.96341, 49.98101, 
    49.99837, 50.01548, 50.03234, 50.04895, 50.06532, 50.08144, 50.09731, 
    50.11294, 50.12831, 50.14344, 50.15832, 50.17295, 50.18733, 50.20147, 
    50.21535, 50.22898, 50.24236, 50.25549, 50.26836, 50.28099, 50.29337, 
    50.30549, 50.31736, 50.32898, 50.34035, 50.35146, 50.36233, 50.37294, 
    50.38329, 50.39339, 50.40324, 50.41283, 50.42218, 50.43126, 50.44009, 
    50.44867, 50.45699, 50.46506, 50.47287, 50.48043, 50.48773, 50.49477, 
    50.50156, 50.50809, 50.51437, 50.5204, 50.52616, 50.53167, 50.53692, 
    50.54192, 50.54666, 50.55114, 50.55537, 50.55934, 50.56305, 50.56651, 
    50.5697, 50.57264, 50.57533, 50.57775, 50.57992, 50.58183, 50.58348, 
    50.58488, 50.58602, 50.5869, 50.58752, 50.58789, 50.588, 50.58785, 
    50.58744, 50.58678, 50.58586, 50.58468, 50.58324, 50.58155, 50.57959, 
    50.57738, 50.57492, 50.57219, 50.56921, 50.56598, 50.56248, 50.55873, 
    50.55472, 50.55045, 50.54593, 50.54115, 50.53611, 50.53082, 50.52526, 
    50.51946, 50.5134, 50.50708, 50.5005, 50.49368, 50.48659, 50.47925, 
    50.47165, 50.4638, 50.45569, 50.44733, 50.43871, 50.42984, 50.42072, 
    50.41133, 50.4017, 50.39181, 50.38167, 50.37127, 50.36063, 50.34972, 
    50.33857, 50.32716, 50.3155, 50.30359, 50.29143, 50.27901, 50.26634, 
    50.25343, 50.24026, 50.22684, 50.21317, 50.19925, 50.18507, 50.17065, 
    50.15599, 50.14107, 50.1259, 50.11049, 50.09482, 50.07891, 50.06275, 
    50.04634, 50.02969, 50.01279, 49.99564, 49.97825, 49.96061, 49.94273, 
    49.92459, 49.90622, 49.8876, 49.86874, 49.84964, 49.83029, 49.8107, 
    49.79086, 49.77078, 49.75047, 49.7299, 49.70911, 49.68806, 49.66678, 
    49.64526, 49.6235, 49.6015, 49.57926, 49.55678, 49.53407, 49.51111, 
    49.48792, 49.4645, 49.44083, 49.41693, 49.3928, 49.36843, 49.34383, 
    49.31899, 49.29392, 49.26862, 49.24308, 49.21731, 49.19131, 49.16508, 
    49.13861, 49.11192, 49.085, 49.05784, 49.03046, 49.00285, 48.97501, 
    48.94695, 48.91865, 48.89013, 48.86139, 48.83241, 48.80322, 48.77379, 
    48.74414, 48.71428, 48.68418, 48.65387, 48.62333, 48.59257, 48.56159, 
    48.53038, 48.49896, 48.46732, 48.43546, 48.40338, 48.37108, 48.33857, 
    48.30584, 48.27289, 48.23972, 48.20634, 48.17275, 48.13894, 48.10492, 
    48.07068, 48.03623, 48.00157, 47.96669, 47.93161, 47.89632, 47.86081, 
    47.8251, 47.78917, 47.75304, 47.7167, 47.68015, 47.6434, 47.60644, 
    47.56927, 47.5319, 47.49433, 47.45655, 47.41857, 47.38038, 47.342, 
    47.30341, 47.26461, 47.22562, 47.18643, 47.14704, 47.10745, 47.06767, 
    47.02768, 46.9875,
  42.57225, 42.62831, 42.68423, 42.74, 42.79563, 42.85111, 42.90645, 
    42.96164, 43.01668, 43.07157, 43.12631, 43.18091, 43.23536, 43.28965, 
    43.3438, 43.39779, 43.45163, 43.50532, 43.55886, 43.61224, 43.66547, 
    43.71854, 43.77146, 43.82422, 43.87683, 43.92928, 43.98157, 44.0337, 
    44.08568, 44.13749, 44.18915, 44.24065, 44.29198, 44.34315, 44.39417, 
    44.44501, 44.4957, 44.54622, 44.59658, 44.64677, 44.6968, 44.74666, 
    44.79636, 44.84589, 44.89524, 44.94444, 44.99346, 45.04231, 45.091, 
    45.13951, 45.18785, 45.23602, 45.28401, 45.33184, 45.37949, 45.42696, 
    45.47426, 45.52139, 45.56834, 45.61511, 45.66171, 45.70813, 45.75437, 
    45.80043, 45.84631, 45.89201, 45.93753, 45.98288, 46.02803, 46.07301, 
    46.1178, 46.16241, 46.20684, 46.25108, 46.29514, 46.339, 46.38269, 
    46.42619, 46.46949, 46.51262, 46.55555, 46.59829, 46.64084, 46.6832, 
    46.72538, 46.76736, 46.80914, 46.85074, 46.89214, 46.93335, 46.97436, 
    47.01518, 47.0558, 47.09623, 47.13645, 47.17648, 47.21632, 47.25595, 
    47.29539, 47.33462, 47.37366, 47.41249, 47.45113, 47.48956, 47.52778, 
    47.56581, 47.60363, 47.64125, 47.67866, 47.71587, 47.75287, 47.78966, 
    47.82625, 47.86263, 47.8988, 47.93476, 47.97052, 48.00606, 48.04139, 
    48.07652, 48.11143, 48.14613, 48.18061, 48.21488, 48.24894, 48.28279, 
    48.31642, 48.34983, 48.38303, 48.41601, 48.44878, 48.48133, 48.51366, 
    48.54577, 48.57766, 48.60933, 48.64079, 48.67202, 48.70303, 48.73382, 
    48.76439, 48.79473, 48.82485, 48.85475, 48.88442, 48.91387, 48.9431, 
    48.9721, 49.00087, 49.02941, 49.05773, 49.08582, 49.11369, 49.14132, 
    49.16872, 49.1959, 49.22284, 49.24956, 49.27604, 49.3023, 49.32832, 
    49.3541, 49.37966, 49.40498, 49.43007, 49.45493, 49.47955, 49.50393, 
    49.52808, 49.55199, 49.57567, 49.59911, 49.62231, 49.64528, 49.66801, 
    49.6905, 49.71275, 49.73476, 49.75653, 49.77806, 49.79935, 49.82041, 
    49.84122, 49.86178, 49.88211, 49.90219, 49.92203, 49.94163, 49.96098, 
    49.98009, 49.99896, 50.01758, 50.03596, 50.05409, 50.07198, 50.08961, 
    50.10701, 50.12415, 50.14106, 50.15771, 50.17411, 50.19027, 50.20618, 
    50.22184, 50.23725, 50.25241, 50.26733, 50.28199, 50.2964, 50.31057, 
    50.32448, 50.33814, 50.35155, 50.36471, 50.37762, 50.39028, 50.40268, 
    50.41483, 50.42673, 50.43838, 50.44977, 50.46091, 50.4718, 50.48243, 
    50.49281, 50.50294, 50.51281, 50.52243, 50.53179, 50.54089, 50.54975, 
    50.55834, 50.56668, 50.57477, 50.5826, 50.59018, 50.59749, 50.60455, 
    50.61136, 50.61791, 50.6242, 50.63024, 50.63602, 50.64154, 50.6468, 
    50.65181, 50.65656, 50.66106, 50.66529, 50.66927, 50.67299, 50.67645, 
    50.67966, 50.68261, 50.6853, 50.68773, 50.6899, 50.69182, 50.69347, 
    50.69487, 50.69601, 50.6969, 50.69753, 50.69789, 50.698, 50.69785, 
    50.69744, 50.69678, 50.69585, 50.69467, 50.69323, 50.69153, 50.68958, 
    50.68736, 50.68489, 50.68216, 50.67917, 50.67592, 50.67242, 50.66866, 
    50.66464, 50.66036, 50.65583, 50.65104, 50.64599, 50.64068, 50.63512, 
    50.6293, 50.62322, 50.61689, 50.6103, 50.60345, 50.59635, 50.58899, 
    50.58138, 50.57351, 50.56538, 50.557, 50.54836, 50.53947, 50.53032, 
    50.52092, 50.51126, 50.50135, 50.49119, 50.48077, 50.4701, 50.45917, 
    50.44799, 50.43655, 50.42487, 50.41293, 50.40074, 50.38829, 50.3756, 
    50.36265, 50.34945, 50.336, 50.3223, 50.30834, 50.29414, 50.27969, 
    50.26498, 50.25003, 50.23483, 50.21938, 50.20368, 50.18773, 50.17154, 
    50.15509, 50.1384, 50.12146, 50.10427, 50.08684, 50.06916, 50.05124, 
    50.03307, 50.01465, 49.99599, 49.97709, 49.95794, 49.93855, 49.91891, 
    49.89903, 49.87891, 49.85855, 49.83794, 49.81709, 49.79601, 49.77467, 
    49.75311, 49.7313, 49.70925, 49.68696, 49.66443, 49.64167, 49.61866, 
    49.59542, 49.57194, 49.54823, 49.52428, 49.50009, 49.47567, 49.45101, 
    49.42612, 49.40099, 49.37563, 49.35004, 49.32421, 49.29816, 49.27187, 
    49.24535, 49.2186, 49.19162, 49.1644, 49.13696, 49.10929, 49.08139, 
    49.05326, 49.02491, 48.99633, 48.96752, 48.93849, 48.90923, 48.87975, 
    48.85004, 48.8201, 48.78994, 48.75956, 48.72896, 48.69814, 48.66709, 
    48.63583, 48.60434, 48.57263, 48.5407, 48.50856, 48.47619, 48.44361, 
    48.41081, 48.37779, 48.34456, 48.31111, 48.27745, 48.24357, 48.20948, 
    48.17517, 48.14065, 48.10592, 48.07097, 48.03582, 48.00045, 47.96487, 
    47.92909, 47.89309, 47.85689, 47.82048, 47.78386, 47.74703, 47.71, 
    47.67276, 47.63531, 47.59766, 47.55981, 47.52175, 47.48349, 47.44503, 
    47.40636, 47.3675, 47.32843, 47.28916, 47.24969, 47.21003, 47.17017, 
    47.1301, 47.08984,
  42.66682, 42.72297, 42.77897, 42.83483, 42.89054, 42.94611, 43.00153, 
    43.05681, 43.11193, 43.16691, 43.22174, 43.27642, 43.33096, 43.38533, 
    43.43956, 43.49364, 43.54757, 43.60135, 43.65497, 43.70844, 43.76175, 
    43.81491, 43.86791, 43.92076, 43.97345, 44.02599, 44.07837, 44.13058, 
    44.18264, 44.23455, 44.28629, 44.33787, 44.38929, 44.44055, 44.49165, 
    44.54258, 44.59335, 44.64396, 44.6944, 44.74467, 44.79479, 44.84473, 
    44.89451, 44.94413, 44.99357, 45.04285, 45.09195, 45.14089, 45.18966, 
    45.23825, 45.28668, 45.33493, 45.38301, 45.43092, 45.47865, 45.52621, 
    45.5736, 45.6208, 45.66784, 45.71469, 45.76138, 45.80788, 45.8542, 
    45.90034, 45.94631, 45.99209, 46.0377, 46.08312, 46.12836, 46.17342, 
    46.21829, 46.26299, 46.30749, 46.35181, 46.39595, 46.4399, 46.48367, 
    46.52724, 46.57063, 46.61383, 46.65685, 46.69967, 46.7423, 46.78474, 
    46.827, 46.86905, 46.91092, 46.95259, 46.99408, 47.03536, 47.07645, 
    47.11735, 47.15805, 47.19855, 47.23886, 47.27896, 47.31887, 47.35859, 
    47.3981, 47.43741, 47.47652, 47.51543, 47.55414, 47.59265, 47.63095, 
    47.66905, 47.70695, 47.74464, 47.78213, 47.81941, 47.85648, 47.89335, 
    47.93001, 47.96646, 48.00271, 48.03874, 48.07457, 48.11018, 48.14559, 
    48.18078, 48.21576, 48.25053, 48.28509, 48.31943, 48.35356, 48.38747, 
    48.42117, 48.45465, 48.48792, 48.52097, 48.55381, 48.58642, 48.61882, 
    48.651, 48.68296, 48.7147, 48.74622, 48.77751, 48.80859, 48.83944, 
    48.87008, 48.90049, 48.93067, 48.96063, 48.99037, 49.01988, 49.04917, 
    49.07822, 49.10706, 49.13567, 49.16404, 49.1922, 49.22012, 49.24781, 
    49.27528, 49.30251, 49.32951, 49.35629, 49.38283, 49.40914, 49.43521, 
    49.46106, 49.48667, 49.51205, 49.53719, 49.5621, 49.58678, 49.61121, 
    49.63542, 49.65939, 49.68311, 49.70661, 49.72986, 49.75288, 49.77566, 
    49.79819, 49.8205, 49.84256, 49.86438, 49.88596, 49.9073, 49.92839, 
    49.94925, 49.96986, 49.99023, 50.01036, 50.03025, 50.04989, 50.06929, 
    50.08844, 50.10735, 50.12601, 50.14443, 50.1626, 50.18053, 50.19821, 
    50.21564, 50.23283, 50.24976, 50.26646, 50.2829, 50.29909, 50.31504, 
    50.33073, 50.34618, 50.36138, 50.37633, 50.39102, 50.40547, 50.41967, 
    50.43361, 50.4473, 50.46075, 50.47393, 50.48687, 50.49956, 50.51199, 
    50.52417, 50.5361, 50.54777, 50.55919, 50.57036, 50.58127, 50.59193, 
    50.60233, 50.61248, 50.62238, 50.63202, 50.6414, 50.65053, 50.6594, 
    50.66801, 50.67638, 50.68448, 50.69233, 50.69992, 50.70726, 50.71434, 
    50.72116, 50.72772, 50.73403, 50.74008, 50.74587, 50.75141, 50.75668, 
    50.7617, 50.76646, 50.77097, 50.77522, 50.7792, 50.78293, 50.7864, 
    50.78962, 50.79257, 50.79527, 50.7977, 50.79988, 50.8018, 50.80346, 
    50.80487, 50.80601, 50.8069, 50.80752, 50.80789, 50.808, 50.80785, 
    50.80744, 50.80677, 50.80585, 50.80466, 50.80322, 50.80152, 50.79956, 
    50.79734, 50.79486, 50.79212, 50.78912, 50.78587, 50.78236, 50.77859, 
    50.77456, 50.77028, 50.76573, 50.76093, 50.75587, 50.75055, 50.74497, 
    50.73914, 50.73305, 50.7267, 50.72009, 50.71323, 50.70611, 50.69874, 
    50.6911, 50.68322, 50.67507, 50.66667, 50.65801, 50.6491, 50.63993, 
    50.63051, 50.62083, 50.61089, 50.6007, 50.59026, 50.57956, 50.56861, 
    50.5574, 50.54594, 50.53423, 50.52226, 50.51004, 50.49757, 50.48484, 
    50.47187, 50.45864, 50.44516, 50.43142, 50.41744, 50.4032, 50.38871, 
    50.37398, 50.35899, 50.34375, 50.32827, 50.31253, 50.29655, 50.28032, 
    50.26383, 50.2471, 50.23013, 50.2129, 50.19543, 50.17771, 50.15974, 
    50.14153, 50.12307, 50.10437, 50.08543, 50.06623, 50.0468, 50.02712, 
    50.00719, 49.98703, 49.96662, 49.94596, 49.92507, 49.90393, 49.88256, 
    49.86094, 49.83908, 49.81698, 49.79465, 49.77207, 49.74925, 49.7262, 
    49.70291, 49.67937, 49.65561, 49.6316, 49.60736, 49.58289, 49.55818, 
    49.53323, 49.50805, 49.48264, 49.45699, 49.43111, 49.40499, 49.37865, 
    49.35207, 49.32526, 49.29822, 49.27095, 49.24345, 49.21572, 49.18776, 
    49.15957, 49.13116, 49.10251, 49.07364, 49.04455, 49.01523, 48.98568, 
    48.95591, 48.92591, 48.89569, 48.86525, 48.83458, 48.80369, 48.77258, 
    48.74125, 48.70969, 48.67792, 48.64592, 48.61371, 48.58128, 48.54863, 
    48.51576, 48.48268, 48.44938, 48.41586, 48.38212, 48.34818, 48.31401, 
    48.27964, 48.24504, 48.21024, 48.17523, 48.14, 48.10456, 48.06892, 
    48.03305, 47.99699, 47.96071, 47.92422, 47.88753, 47.85063, 47.81352, 
    47.77621, 47.73869, 47.70097, 47.66304, 47.6249, 47.58657, 47.54803, 
    47.50929, 47.47035, 47.43121, 47.39186, 47.35232, 47.31258, 47.27263, 
    47.23249, 47.19216,
  42.76134, 42.81758, 42.87367, 42.92961, 42.98541, 43.04106, 43.09657, 
    43.15193, 43.20714, 43.26221, 43.31712, 43.37189, 43.42651, 43.48097, 
    43.53529, 43.58945, 43.64346, 43.69732, 43.75103, 43.80458, 43.85799, 
    43.91123, 43.96432, 44.01725, 44.07003, 44.12265, 44.17511, 44.22742, 
    44.27956, 44.33155, 44.38338, 44.43505, 44.48655, 44.5379, 44.58908, 
    44.64009, 44.69095, 44.74165, 44.79217, 44.84253, 44.89273, 44.94276, 
    44.99263, 45.04232, 45.09185, 45.14121, 45.1904, 45.23943, 45.28828, 
    45.33696, 45.38547, 45.4338, 45.48197, 45.52996, 45.57778, 45.62542, 
    45.67289, 45.72018, 45.7673, 45.81424, 45.861, 45.90759, 45.95399, 
    46.00022, 46.04626, 46.09213, 46.13782, 46.18332, 46.22865, 46.27379, 
    46.31874, 46.36352, 46.40811, 46.45251, 46.49673, 46.54076, 46.58461, 
    46.62827, 46.67174, 46.71502, 46.75811, 46.80101, 46.84373, 46.88625, 
    46.92858, 46.97072, 47.01266, 47.05442, 47.09598, 47.13734, 47.17851, 
    47.21949, 47.26027, 47.30085, 47.34123, 47.38142, 47.4214, 47.46119, 
    47.50078, 47.54017, 47.57936, 47.61834, 47.65713, 47.69571, 47.73409, 
    47.77227, 47.81024, 47.848, 47.88557, 47.92292, 47.96007, 47.99701, 
    48.03374, 48.07027, 48.10659, 48.1427, 48.17859, 48.21428, 48.24976, 
    48.28502, 48.32008, 48.35492, 48.38954, 48.42395, 48.45815, 48.49214, 
    48.52591, 48.55946, 48.5928, 48.62592, 48.65882, 48.6915, 48.72396, 
    48.75621, 48.78823, 48.82004, 48.85163, 48.88299, 48.91413, 48.94505, 
    48.97575, 49.00622, 49.03647, 49.06649, 49.09629, 49.12587, 49.15522, 
    49.18434, 49.21323, 49.24191, 49.27034, 49.29855, 49.32654, 49.35429, 
    49.38181, 49.40911, 49.43617, 49.463, 49.4896, 49.51597, 49.5421, 49.568, 
    49.59367, 49.6191, 49.6443, 49.66927, 49.69399, 49.71849, 49.74274, 
    49.76676, 49.79054, 49.81409, 49.83739, 49.86046, 49.88329, 49.90588, 
    49.92823, 49.95034, 49.97221, 49.99384, 50.01522, 50.03637, 50.05727, 
    50.07793, 50.09835, 50.11852, 50.13845, 50.15814, 50.17758, 50.19678, 
    50.21573, 50.23443, 50.2529, 50.27111, 50.28907, 50.30679, 50.32427, 
    50.34149, 50.35847, 50.3752, 50.39168, 50.40791, 50.42389, 50.43962, 
    50.4551, 50.47034, 50.48532, 50.50005, 50.51453, 50.52876, 50.54274, 
    50.55646, 50.56993, 50.58316, 50.59612, 50.60884, 50.6213, 50.63351, 
    50.64546, 50.65717, 50.66861, 50.6798, 50.69074, 50.70142, 50.71185, 
    50.72202, 50.73194, 50.7416, 50.75101, 50.76015, 50.76905, 50.77769, 
    50.78607, 50.79419, 50.80206, 50.80967, 50.81702, 50.82412, 50.83095, 
    50.83753, 50.84385, 50.84992, 50.85572, 50.86127, 50.86656, 50.87159, 
    50.87637, 50.88088, 50.88514, 50.88913, 50.89287, 50.89635, 50.89957, 
    50.90253, 50.90524, 50.90768, 50.90986, 50.91179, 50.91345, 50.91486, 
    50.916, 50.91689, 50.91752, 50.91789, 50.918, 50.91785, 50.91744, 
    50.91677, 50.91584, 50.91465, 50.91321, 50.9115, 50.90953, 50.90731, 
    50.90483, 50.90208, 50.89908, 50.89582, 50.8923, 50.88852, 50.88448, 
    50.88018, 50.87563, 50.87082, 50.86574, 50.86041, 50.85482, 50.84898, 
    50.84287, 50.83651, 50.82989, 50.82301, 50.81587, 50.80848, 50.80083, 
    50.79292, 50.78476, 50.77634, 50.76766, 50.75873, 50.74953, 50.74009, 
    50.73039, 50.72043, 50.71022, 50.69975, 50.68903, 50.67805, 50.66682, 
    50.65533, 50.64359, 50.6316, 50.61935, 50.60685, 50.59409, 50.58108, 
    50.56782, 50.55431, 50.54054, 50.52653, 50.51226, 50.49774, 50.48297, 
    50.46795, 50.45267, 50.43715, 50.42138, 50.40536, 50.38909, 50.37257, 
    50.3558, 50.33878, 50.32152, 50.30401, 50.28625, 50.26824, 50.24999, 
    50.23149, 50.21275, 50.19376, 50.17452, 50.15504, 50.13531, 50.11535, 
    50.09513, 50.07468, 50.05398, 50.03304, 50.01186, 49.99043, 49.96877, 
    49.94686, 49.92471, 49.90232, 49.8797, 49.85683, 49.83372, 49.81038, 
    49.7868, 49.76298, 49.73892, 49.71463, 49.6901, 49.66533, 49.64033, 
    49.6151, 49.58963, 49.56392, 49.53798, 49.51181, 49.48541, 49.45877, 
    49.4319, 49.4048, 49.37748, 49.34991, 49.32213, 49.29411, 49.26586, 
    49.23738, 49.20868, 49.17975, 49.15059, 49.12121, 49.09159, 49.06176, 
    49.0317, 49.00142, 48.97091, 48.94017, 48.90922, 48.87804, 48.84665, 
    48.81503, 48.78318, 48.75113, 48.71885, 48.68634, 48.65363, 48.62069, 
    48.58754, 48.55416, 48.52058, 48.48678, 48.45276, 48.41853, 48.38408, 
    48.34942, 48.31454, 48.27946, 48.24416, 48.20865, 48.17293, 48.137, 
    48.10086, 48.06451, 48.02795, 47.99118, 47.95421, 47.91703, 47.87964, 
    47.84204, 47.80424, 47.76624, 47.72803, 47.68962, 47.65101, 47.61219, 
    47.57317, 47.53395, 47.49453, 47.45491, 47.41509, 47.37507, 47.33485, 
    47.29444,
  42.85582, 42.91214, 42.96831, 43.02434, 43.08022, 43.13596, 43.19156, 
    43.247, 43.3023, 43.35745, 43.41245, 43.4673, 43.52201, 43.57656, 
    43.63096, 43.68521, 43.73931, 43.79325, 43.84705, 43.90069, 43.95417, 
    44.0075, 44.06068, 44.1137, 44.16656, 44.21927, 44.27182, 44.32421, 
    44.37644, 44.42851, 44.48042, 44.53218, 44.58377, 44.6352, 44.68647, 
    44.73757, 44.78851, 44.83929, 44.8899, 44.94035, 44.99063, 45.04075, 
    45.09069, 45.14048, 45.19009, 45.23954, 45.28881, 45.33792, 45.38686, 
    45.43562, 45.48421, 45.53263, 45.58088, 45.62896, 45.67686, 45.72459, 
    45.77214, 45.81952, 45.86672, 45.91374, 45.96059, 46.00726, 46.05375, 
    46.10006, 46.14619, 46.19213, 46.23791, 46.28349, 46.3289, 46.37412, 
    46.41916, 46.46402, 46.50869, 46.55317, 46.59747, 46.64159, 46.68552, 
    46.72926, 46.77281, 46.81617, 46.85934, 46.90233, 46.94512, 46.98772, 
    47.03013, 47.07235, 47.11438, 47.15621, 47.19785, 47.23929, 47.28054, 
    47.32159, 47.36245, 47.40311, 47.44357, 47.48384, 47.5239, 47.56377, 
    47.60343, 47.6429, 47.68216, 47.72123, 47.76009, 47.79875, 47.8372, 
    47.87545, 47.9135, 47.95134, 47.98898, 48.02641, 48.06363, 48.10065, 
    48.13745, 48.17405, 48.21045, 48.24662, 48.2826, 48.31836, 48.3539, 
    48.38924, 48.42437, 48.45927, 48.49397, 48.52846, 48.56273, 48.59678, 
    48.63062, 48.66424, 48.69765, 48.73083, 48.76381, 48.79655, 48.82909, 
    48.8614, 48.89349, 48.92537, 48.95702, 48.98845, 49.01965, 49.05064, 
    49.0814, 49.11194, 49.14225, 49.17234, 49.20221, 49.23184, 49.26125, 
    49.29044, 49.3194, 49.34813, 49.37663, 49.4049, 49.43294, 49.46075, 
    49.48834, 49.51569, 49.54281, 49.5697, 49.59636, 49.62278, 49.64897, 
    49.67493, 49.70065, 49.72614, 49.7514, 49.77642, 49.8012, 49.82574, 
    49.85006, 49.87413, 49.89796, 49.92156, 49.94492, 49.96804, 49.99092, 
    50.01356, 50.03596, 50.05812, 50.08003, 50.10171, 50.12315, 50.14434, 
    50.16529, 50.18599, 50.20646, 50.22668, 50.24665, 50.26638, 50.28587, 
    50.30511, 50.3241, 50.34285, 50.36135, 50.3796, 50.39761, 50.41537, 
    50.43289, 50.45015, 50.46717, 50.48394, 50.50045, 50.51672, 50.53274, 
    50.54851, 50.56403, 50.57929, 50.59431, 50.60907, 50.62359, 50.63785, 
    50.65186, 50.66562, 50.67912, 50.69237, 50.70537, 50.71811, 50.73061, 
    50.74284, 50.75483, 50.76655, 50.77803, 50.78924, 50.80021, 50.81091, 
    50.82137, 50.83156, 50.8415, 50.85118, 50.86061, 50.86979, 50.8787, 
    50.88736, 50.89576, 50.9039, 50.91179, 50.91941, 50.92678, 50.93389, 
    50.94075, 50.94734, 50.95368, 50.95976, 50.96558, 50.97114, 50.97644, 
    50.98148, 50.98627, 50.9908, 50.99506, 50.99907, 51.00282, 51.0063, 
    51.00953, 51.0125, 51.01521, 51.01765, 51.01984, 51.02177, 51.02344, 
    51.02485, 51.026, 51.02689, 51.02752, 51.02789, 51.028, 51.02785, 
    51.02744, 51.02677, 51.02584, 51.02465, 51.0232, 51.02148, 51.01952, 
    51.01728, 51.01479, 51.01205, 51.00904, 51.00577, 51.00224, 50.99845, 
    50.9944, 50.9901, 50.98553, 50.98071, 50.97562, 50.97028, 50.96468, 
    50.95881, 50.95269, 50.94632, 50.93968, 50.93279, 50.92563, 50.91822, 
    50.91055, 50.90263, 50.89444, 50.88601, 50.87731, 50.86835, 50.85914, 
    50.84967, 50.83995, 50.82997, 50.81973, 50.80924, 50.79849, 50.78749, 
    50.77623, 50.76471, 50.75294, 50.74092, 50.72865, 50.71611, 50.70333, 
    50.69029, 50.677, 50.66346, 50.64966, 50.63561, 50.62131, 50.60675, 
    50.59195, 50.5769, 50.56159, 50.54603, 50.53022, 50.51416, 50.49786, 
    50.4813, 50.46449, 50.44744, 50.43013, 50.41258, 50.39478, 50.37674, 
    50.35844, 50.3399, 50.32111, 50.30208, 50.2828, 50.26328, 50.24351, 
    50.22349, 50.20324, 50.18274, 50.16199, 50.141, 50.11977, 50.0983, 
    50.07658, 50.05463, 50.03243, 50.00999, 49.98731, 49.9644, 49.94124, 
    49.91784, 49.89421, 49.87033, 49.84623, 49.82188, 49.79729, 49.77248, 
    49.74742, 49.72213, 49.6966, 49.67084, 49.64484, 49.61862, 49.59216, 
    49.56546, 49.53854, 49.51138, 49.48399, 49.45637, 49.42852, 49.40044, 
    49.37213, 49.34359, 49.31483, 49.28584, 49.25661, 49.22717, 49.19749, 
    49.16759, 49.13747, 49.10712, 49.07655, 49.04575, 49.01473, 48.98349, 
    48.95203, 48.92034, 48.88843, 48.8563, 48.82396, 48.79139, 48.7586, 
    48.7256, 48.69238, 48.65894, 48.62528, 48.59141, 48.55732, 48.52302, 
    48.4885, 48.45377, 48.41882, 48.38366, 48.34829, 48.31271, 48.27692, 
    48.24092, 48.2047, 48.16828, 48.13165, 48.0948, 48.05775, 48.0205, 
    47.98304, 47.94537, 47.90749, 47.86942, 47.83113, 47.79264, 47.75396, 
    47.71506, 47.67596, 47.63667, 47.59717, 47.55747, 47.51758, 47.47748, 
    47.43718, 47.39669,
  42.95024, 43.00664, 43.0629, 43.11902, 43.17499, 43.23081, 43.28649, 
    43.34202, 43.39741, 43.45264, 43.50773, 43.56267, 43.61746, 43.6721, 
    43.72659, 43.78092, 43.83511, 43.88914, 43.94302, 43.99674, 44.05031, 
    44.10373, 44.15699, 44.2101, 44.26305, 44.31584, 44.36847, 44.42095, 
    44.47327, 44.52542, 44.57742, 44.62926, 44.68094, 44.73245, 44.78381, 
    44.835, 44.88602, 44.93689, 44.98759, 45.03812, 45.08849, 45.13869, 
    45.18872, 45.23859, 45.28829, 45.33782, 45.38718, 45.43637, 45.48539, 
    45.53424, 45.58292, 45.63143, 45.67976, 45.72792, 45.77591, 45.82372, 
    45.87135, 45.91882, 45.9661, 46.01321, 46.06013, 46.10689, 46.15346, 
    46.19986, 46.24607, 46.2921, 46.33796, 46.38363, 46.42911, 46.47442, 
    46.51954, 46.56448, 46.60923, 46.6538, 46.69818, 46.74238, 46.78638, 
    46.83021, 46.87384, 46.91729, 46.96054, 47.0036, 47.04648, 47.08916, 
    47.13165, 47.17395, 47.21606, 47.25797, 47.29969, 47.34121, 47.38254, 
    47.42367, 47.4646, 47.50534, 47.54588, 47.58622, 47.62637, 47.66631, 
    47.70605, 47.7456, 47.78494, 47.82408, 47.86302, 47.90175, 47.94028, 
    47.97861, 48.01674, 48.05465, 48.09236, 48.12987, 48.16716, 48.20425, 
    48.24113, 48.27781, 48.31427, 48.35053, 48.38657, 48.42241, 48.45802, 
    48.49343, 48.52863, 48.56361, 48.59838, 48.63293, 48.66727, 48.7014, 
    48.73531, 48.769, 48.80247, 48.83573, 48.86877, 48.90159, 48.93419, 
    48.96657, 48.99873, 49.03067, 49.06239, 49.09388, 49.12516, 49.15621, 
    49.18703, 49.21764, 49.24802, 49.27817, 49.30809, 49.3378, 49.36727, 
    49.39652, 49.42554, 49.45433, 49.48289, 49.51123, 49.53933, 49.5672, 
    49.59484, 49.62226, 49.64944, 49.67638, 49.7031, 49.72958, 49.75583, 
    49.78185, 49.80762, 49.83317, 49.85848, 49.88356, 49.90839, 49.93299, 
    49.95736, 49.98148, 50.00537, 50.02902, 50.05243, 50.0756, 50.09853, 
    50.12122, 50.14367, 50.16588, 50.18785, 50.20957, 50.23106, 50.2523, 
    50.27329, 50.29404, 50.31456, 50.33482, 50.35484, 50.37461, 50.39415, 
    50.41343, 50.43246, 50.45126, 50.4698, 50.4881, 50.50615, 50.52395, 
    50.5415, 50.5588, 50.57586, 50.59267, 50.60922, 50.62553, 50.64158, 
    50.65739, 50.67294, 50.68824, 50.7033, 50.71809, 50.73264, 50.74694, 
    50.76098, 50.77477, 50.7883, 50.80158, 50.81461, 50.82738, 50.8399, 
    50.85217, 50.86418, 50.87594, 50.88744, 50.89868, 50.90967, 50.9204, 
    50.93088, 50.9411, 50.95106, 50.96077, 50.97022, 50.97941, 50.98835, 
    50.99702, 51.00544, 51.01361, 51.02151, 51.02916, 51.03654, 51.04367, 
    51.05054, 51.05715, 51.0635, 51.0696, 51.07543, 51.08101, 51.08632, 
    51.09137, 51.09617, 51.1007, 51.10498, 51.109, 51.11275, 51.11625, 
    51.11948, 51.12246, 51.12518, 51.12763, 51.12983, 51.13176, 51.13343, 
    51.13485, 51.136, 51.13689, 51.13752, 51.13789, 51.138, 51.13785, 
    51.13744, 51.13676, 51.13583, 51.13464, 51.13318, 51.13147, 51.12949, 
    51.12726, 51.12476, 51.12201, 51.11899, 51.11572, 51.11218, 51.10838, 
    51.10432, 51.10001, 51.09543, 51.09059, 51.08549, 51.08014, 51.07452, 
    51.06865, 51.06252, 51.05612, 51.04947, 51.04256, 51.03539, 51.02796, 
    51.02028, 51.01233, 51.00413, 50.99567, 50.98695, 50.97797, 50.96874, 
    50.95925, 50.9495, 50.9395, 50.92924, 50.91872, 50.90795, 50.89692, 
    50.88564, 50.8741, 50.8623, 50.85025, 50.83794, 50.82538, 50.81257, 
    50.7995, 50.78618, 50.7726, 50.75877, 50.74469, 50.73036, 50.71577, 
    50.70093, 50.68584, 50.6705, 50.6549, 50.63906, 50.62296, 50.60662, 
    50.59002, 50.57318, 50.55608, 50.53874, 50.52115, 50.50331, 50.48522, 
    50.46688, 50.4483, 50.42947, 50.41039, 50.39107, 50.3715, 50.35169, 
    50.33163, 50.31133, 50.29078, 50.26999, 50.24895, 50.22767, 50.20615, 
    50.18439, 50.16238, 50.14014, 50.11765, 50.09492, 50.07195, 50.04874, 
    50.0253, 50.00161, 49.97768, 49.95352, 49.92912, 49.90448, 49.8796, 
    49.85449, 49.82915, 49.80356, 49.77775, 49.75169, 49.72541, 49.69889, 
    49.67214, 49.64515, 49.61794, 49.59049, 49.56281, 49.5349, 49.50676, 
    49.47839, 49.44979, 49.42096, 49.39191, 49.36263, 49.33311, 49.30338, 
    49.27341, 49.24323, 49.21281, 49.18217, 49.15131, 49.12022, 49.08892, 
    49.05738, 49.02563, 48.99366, 48.96146, 48.92905, 48.89641, 48.86356, 
    48.83049, 48.7972, 48.76369, 48.72996, 48.69602, 48.66186, 48.62748, 
    48.5929, 48.55809, 48.52308, 48.48785, 48.4524, 48.41675, 48.38088, 
    48.34481, 48.30852, 48.27202, 48.23532, 48.1984, 48.16128, 48.12395, 
    48.08641, 48.04867, 48.01072, 47.97256, 47.9342, 47.89564, 47.85687, 
    47.8179, 47.77873, 47.73936, 47.69978, 47.66001, 47.62003, 47.57986, 
    47.53948, 47.49891,
  43.04461, 43.1011, 43.15744, 43.21365, 43.2697, 43.32561, 43.38137, 
    43.43699, 43.49246, 43.54779, 43.60296, 43.65799, 43.71286, 43.76758, 
    43.82216, 43.87658, 43.93085, 43.98497, 44.03894, 44.09275, 44.1464, 
    44.19991, 44.25325, 44.30645, 44.35948, 44.41236, 44.46508, 44.51764, 
    44.57005, 44.62229, 44.67438, 44.7263, 44.77806, 44.82966, 44.8811, 
    44.93238, 44.98349, 45.03444, 45.08522, 45.13585, 45.1863, 45.23658, 
    45.28671, 45.33665, 45.38644, 45.43606, 45.4855, 45.53478, 45.58389, 
    45.63282, 45.68158, 45.73018, 45.77859, 45.82684, 45.87491, 45.9228, 
    45.97052, 46.01807, 46.06544, 46.11263, 46.15965, 46.20648, 46.25314, 
    46.29961, 46.34591, 46.39203, 46.43796, 46.48372, 46.52929, 46.57468, 
    46.61988, 46.6649, 46.70974, 46.75439, 46.79885, 46.84313, 46.88722, 
    46.93113, 46.97484, 47.01836, 47.0617, 47.10485, 47.1478, 47.19056, 
    47.23314, 47.27552, 47.3177, 47.35969, 47.40149, 47.44309, 47.4845, 
    47.52571, 47.56673, 47.60754, 47.64816, 47.68858, 47.72881, 47.76883, 
    47.80865, 47.84827, 47.88769, 47.92691, 47.96592, 48.00473, 48.04334, 
    48.08174, 48.11994, 48.15793, 48.19572, 48.2333, 48.27067, 48.30783, 
    48.34479, 48.38154, 48.41808, 48.45441, 48.49052, 48.52643, 48.56212, 
    48.5976, 48.63287, 48.66793, 48.70277, 48.73739, 48.7718, 48.806, 
    48.83997, 48.87374, 48.90728, 48.94061, 48.97371, 49.0066, 49.03927, 
    49.07172, 49.10395, 49.13596, 49.16774, 49.1993, 49.23064, 49.26176, 
    49.29265, 49.32332, 49.35376, 49.38398, 49.41397, 49.44373, 49.47327, 
    49.50258, 49.53166, 49.56052, 49.58914, 49.61753, 49.6457, 49.67363, 
    49.70134, 49.72881, 49.75605, 49.78305, 49.80983, 49.83637, 49.86267, 
    49.88875, 49.91459, 49.94019, 49.96555, 49.99068, 50.01557, 50.04023, 
    50.06464, 50.08883, 50.11277, 50.13647, 50.15993, 50.18315, 50.20613, 
    50.22887, 50.25138, 50.27364, 50.29565, 50.31742, 50.33895, 50.36024, 
    50.38129, 50.40209, 50.42265, 50.44296, 50.46302, 50.48284, 50.50241, 
    50.52174, 50.54082, 50.55966, 50.57824, 50.59658, 50.61467, 50.63251, 
    50.65011, 50.66745, 50.68455, 50.70139, 50.71798, 50.73433, 50.75042, 
    50.76626, 50.78185, 50.79719, 50.81227, 50.82711, 50.84169, 50.85602, 
    50.87009, 50.88391, 50.89748, 50.91079, 50.92385, 50.93666, 50.9492, 
    50.9615, 50.97354, 50.98532, 50.99685, 51.00812, 51.01913, 51.02989, 
    51.04039, 51.05064, 51.06062, 51.07035, 51.07982, 51.08904, 51.09799, 
    51.10669, 51.11513, 51.12331, 51.13123, 51.1389, 51.1463, 51.15345, 
    51.16033, 51.16696, 51.17333, 51.17944, 51.18528, 51.19087, 51.1962, 
    51.20126, 51.20607, 51.21062, 51.2149, 51.21893, 51.22269, 51.2262, 
    51.22944, 51.23242, 51.23515, 51.23761, 51.2398, 51.24174, 51.24342, 
    51.24484, 51.24599, 51.24689, 51.24752, 51.24789, 51.248, 51.24785, 
    51.24744, 51.24676, 51.24583, 51.24463, 51.24317, 51.24146, 51.23948, 
    51.23723, 51.23473, 51.23197, 51.22895, 51.22566, 51.22211, 51.21831, 
    51.21424, 51.20992, 51.20533, 51.20048, 51.19537, 51.19, 51.18438, 
    51.17849, 51.17234, 51.16593, 51.15926, 51.15234, 51.14515, 51.1377, 
    51.13, 51.12204, 51.11381, 51.10533, 51.09659, 51.0876, 51.07834, 
    51.06883, 51.05906, 51.04903, 51.03875, 51.02821, 51.01741, 51.00635, 
    50.99504, 50.98347, 50.97165, 50.95957, 50.94724, 50.93465, 50.9218, 
    50.9087, 50.89535, 50.88174, 50.86788, 50.85377, 50.8394, 50.82478, 
    50.80991, 50.79478, 50.7794, 50.76377, 50.74789, 50.73176, 50.71538, 
    50.69874, 50.68186, 50.66473, 50.64734, 50.62971, 50.61183, 50.5937, 
    50.57532, 50.55669, 50.53782, 50.5187, 50.49934, 50.47972, 50.45986, 
    50.43976, 50.41941, 50.39882, 50.37798, 50.35689, 50.33557, 50.314, 
    50.29218, 50.27013, 50.24783, 50.2253, 50.20251, 50.17949, 50.15623, 
    50.13273, 50.10899, 50.08501, 50.0608, 50.03634, 50.01165, 49.98672, 
    49.96156, 49.93615, 49.91051, 49.88464, 49.85853, 49.83219, 49.80561, 
    49.7788, 49.75175, 49.72448, 49.69697, 49.66923, 49.64126, 49.61306, 
    49.58463, 49.55597, 49.52708, 49.49796, 49.46861, 49.43904, 49.40924, 
    49.37921, 49.34896, 49.31848, 49.28778, 49.25685, 49.2257, 49.19432, 
    49.16273, 49.13091, 49.09887, 49.0666, 49.03412, 49.00142, 48.96849, 
    48.93535, 48.90199, 48.86841, 48.83461, 48.8006, 48.76637, 48.73193, 
    48.69727, 48.6624, 48.6273, 48.592, 48.55649, 48.52076, 48.48482, 
    48.44867, 48.41231, 48.37574, 48.33896, 48.30197, 48.26477, 48.22737, 
    48.18975, 48.15194, 48.11391, 48.07568, 48.03725, 47.9986, 47.95976, 
    47.92072, 47.88147, 47.84201, 47.80236, 47.76251, 47.72245, 47.6822, 
    47.64175, 47.6011,
  43.13892, 43.1955, 43.25193, 43.30822, 43.36436, 43.42036, 43.47621, 
    43.53191, 43.58747, 43.64288, 43.69814, 43.75325, 43.80821, 43.86302, 
    43.91768, 43.97219, 44.02655, 44.08075, 44.1348, 44.1887, 44.24245, 
    44.29604, 44.34947, 44.40275, 44.45587, 44.50883, 44.56164, 44.61429, 
    44.66678, 44.71911, 44.77128, 44.82329, 44.87514, 44.92683, 44.97836, 
    45.02972, 45.08091, 45.13195, 45.18282, 45.23352, 45.28407, 45.33443, 
    45.38464, 45.43468, 45.48455, 45.53425, 45.58378, 45.63314, 45.68233, 
    45.73136, 45.7802, 45.82888, 45.87738, 45.92571, 45.97387, 46.02185, 
    46.06966, 46.11728, 46.16474, 46.21201, 46.25911, 46.30603, 46.35277, 
    46.39933, 46.44571, 46.49192, 46.53793, 46.58377, 46.62943, 46.6749, 
    46.72018, 46.76529, 46.81021, 46.85494, 46.89949, 46.94385, 46.98802, 
    47.03201, 47.0758, 47.11941, 47.16283, 47.20605, 47.24909, 47.29193, 
    47.33459, 47.37704, 47.41931, 47.46138, 47.50326, 47.54494, 47.58643, 
    47.62772, 47.66882, 47.70971, 47.75041, 47.79091, 47.83121, 47.87131, 
    47.91121, 47.95091, 47.99041, 48.0297, 48.06879, 48.10768, 48.14636, 
    48.18484, 48.22312, 48.26119, 48.29905, 48.3367, 48.37415, 48.41139, 
    48.44842, 48.48524, 48.52185, 48.55826, 48.59445, 48.63042, 48.66619, 
    48.70175, 48.73709, 48.77221, 48.80713, 48.84182, 48.8763, 48.91057, 
    48.94462, 48.97845, 49.01207, 49.04546, 49.07864, 49.1116, 49.14433, 
    49.17685, 49.20914, 49.24122, 49.27307, 49.3047, 49.33611, 49.36729, 
    49.39825, 49.42898, 49.45949, 49.48977, 49.51982, 49.54965, 49.57925, 
    49.60863, 49.63777, 49.66669, 49.69537, 49.72383, 49.75206, 49.78005, 
    49.80781, 49.83535, 49.86264, 49.88971, 49.91654, 49.94314, 49.96951, 
    49.99563, 50.02153, 50.04718, 50.07261, 50.09779, 50.12274, 50.14745, 
    50.17192, 50.19616, 50.22015, 50.2439, 50.26742, 50.29069, 50.31372, 
    50.33652, 50.35907, 50.38138, 50.40344, 50.42527, 50.44685, 50.46818, 
    50.48928, 50.51012, 50.53072, 50.55108, 50.57119, 50.59106, 50.61068, 
    50.63005, 50.64917, 50.66805, 50.68668, 50.70506, 50.72319, 50.74107, 
    50.75871, 50.77609, 50.79322, 50.81011, 50.82674, 50.84312, 50.85925, 
    50.87513, 50.89075, 50.90613, 50.92125, 50.93612, 50.95073, 50.9651, 
    50.9792, 50.99305, 51.00665, 51.02, 51.03308, 51.04592, 51.0585, 
    51.07082, 51.08289, 51.0947, 51.10625, 51.11755, 51.12859, 51.13937, 
    51.1499, 51.16017, 51.17018, 51.17993, 51.18942, 51.19866, 51.20764, 
    51.21635, 51.22482, 51.23302, 51.24096, 51.24864, 51.25606, 51.26322, 
    51.27013, 51.27677, 51.28315, 51.28927, 51.29513, 51.30073, 51.30607, 
    51.31115, 51.31597, 51.32053, 51.32483, 51.32886, 51.33263, 51.33615, 
    51.3394, 51.34239, 51.34512, 51.34758, 51.34978, 51.35173, 51.35341, 
    51.35483, 51.35599, 51.35688, 51.35752, 51.35789, 51.358, 51.35785, 
    51.35743, 51.35676, 51.35582, 51.35462, 51.35316, 51.35144, 51.34945, 
    51.34721, 51.3447, 51.34193, 51.3389, 51.33561, 51.33205, 51.32824, 
    51.32416, 51.31982, 51.31523, 51.31037, 51.30524, 51.29987, 51.29422, 
    51.28832, 51.28216, 51.27573, 51.26905, 51.26211, 51.2549, 51.24744, 
    51.23972, 51.23174, 51.2235, 51.21499, 51.20623, 51.19722, 51.18794, 
    51.17841, 51.16861, 51.15856, 51.14825, 51.13768, 51.12686, 51.11578, 
    51.10444, 51.09285, 51.081, 51.06889, 51.05653, 51.04391, 51.03103, 
    51.0179, 51.00452, 50.99088, 50.97699, 50.96284, 50.94844, 50.93378, 
    50.91888, 50.90371, 50.8883, 50.87263, 50.85672, 50.84055, 50.82413, 
    50.80746, 50.79053, 50.77336, 50.75594, 50.73826, 50.72034, 50.70217, 
    50.68375, 50.66508, 50.64616, 50.627, 50.60759, 50.58793, 50.56803, 
    50.54788, 50.52748, 50.50684, 50.48595, 50.46482, 50.44345, 50.42183, 
    50.39997, 50.37786, 50.35552, 50.33293, 50.3101, 50.28703, 50.26371, 
    50.24016, 50.21637, 50.19234, 50.16807, 50.14356, 50.11881, 50.09382, 
    50.0686, 50.04314, 50.01745, 49.99152, 49.96535, 49.93895, 49.91231, 
    49.88544, 49.85834, 49.83101, 49.80344, 49.77564, 49.7476, 49.71935, 
    49.69085, 49.66213, 49.63317, 49.604, 49.57458, 49.54495, 49.51508, 
    49.48499, 49.45468, 49.42413, 49.39336, 49.36237, 49.33115, 49.29971, 
    49.26805, 49.23616, 49.20405, 49.17172, 49.13917, 49.1064, 49.0734, 
    49.04019, 49.00676, 48.97311, 48.93925, 48.90516, 48.87086, 48.83635, 
    48.80162, 48.76667, 48.73151, 48.69614, 48.66055, 48.62475, 48.58874, 
    48.55251, 48.51608, 48.47943, 48.44258, 48.40551, 48.36824, 48.33076, 
    48.29307, 48.25518, 48.21708, 48.17877, 48.14026, 48.10154, 48.06262, 
    48.0235, 47.98417, 47.94464, 47.90491, 47.86498, 47.82485, 47.78452, 
    47.74399, 47.70326,
  43.23319, 43.28985, 43.34637, 43.40274, 43.45897, 43.51505, 43.57099, 
    43.62678, 43.68243, 43.73792, 43.79327, 43.84846, 43.90351, 43.95841, 
    44.01316, 44.06775, 44.1222, 44.17649, 44.23063, 44.28461, 44.33844, 
    44.39212, 44.44564, 44.499, 44.55221, 44.60526, 44.65816, 44.71089, 
    44.76347, 44.81588, 44.86814, 44.92024, 44.97217, 45.02395, 45.07556, 
    45.12701, 45.17829, 45.22941, 45.28037, 45.33116, 45.38179, 45.43224, 
    45.48254, 45.53266, 45.58261, 45.6324, 45.68202, 45.73147, 45.78074, 
    45.82985, 45.87878, 45.92754, 45.97613, 46.02455, 46.07279, 46.12085, 
    46.16874, 46.21646, 46.264, 46.31136, 46.35854, 46.40554, 46.45237, 
    46.49902, 46.54548, 46.59176, 46.63787, 46.68379, 46.72953, 46.77508, 
    46.82045, 46.86564, 46.91064, 46.95546, 47.00008, 47.04453, 47.08878, 
    47.13285, 47.17673, 47.22042, 47.26392, 47.30723, 47.35035, 47.39327, 
    47.436, 47.47854, 47.52089, 47.56305, 47.605, 47.64677, 47.68833, 
    47.7297, 47.77087, 47.81185, 47.85263, 47.89321, 47.93359, 47.97376, 
    48.01374, 48.05352, 48.09309, 48.13247, 48.17163, 48.2106, 48.24936, 
    48.28792, 48.32627, 48.36441, 48.40235, 48.44008, 48.4776, 48.51492, 
    48.55202, 48.58892, 48.62561, 48.66208, 48.69835, 48.7344, 48.77024, 
    48.80587, 48.84128, 48.87648, 48.91146, 48.94623, 48.98078, 49.01512, 
    49.04924, 49.08314, 49.11683, 49.15029, 49.18354, 49.21656, 49.24937, 
    49.28196, 49.31432, 49.34646, 49.37838, 49.41008, 49.44155, 49.4728, 
    49.50382, 49.53462, 49.56519, 49.59554, 49.62566, 49.65555, 49.68522, 
    49.71465, 49.74386, 49.77284, 49.80159, 49.83011, 49.85839, 49.88645, 
    49.91427, 49.94186, 49.96922, 49.99635, 50.02324, 50.0499, 50.07632, 
    50.1025, 50.12846, 50.15417, 50.17965, 50.20489, 50.22989, 50.25466, 
    50.27919, 50.30347, 50.32752, 50.35133, 50.3749, 50.39822, 50.42131, 
    50.44415, 50.46675, 50.48911, 50.51123, 50.5331, 50.55473, 50.57611, 
    50.59725, 50.61815, 50.6388, 50.6592, 50.67936, 50.69927, 50.71893, 
    50.73835, 50.75751, 50.77644, 50.79511, 50.81353, 50.8317, 50.84963, 
    50.8673, 50.88473, 50.9019, 50.91882, 50.93549, 50.95191, 50.96808, 
    50.98399, 50.99966, 51.01506, 51.03022, 51.04512, 51.05977, 51.07417, 
    51.08831, 51.10219, 51.11582, 51.1292, 51.14232, 51.15518, 51.16779, 
    51.18014, 51.19224, 51.20407, 51.21566, 51.22698, 51.23804, 51.24886, 
    51.25941, 51.2697, 51.27973, 51.28951, 51.29902, 51.30828, 51.31728, 
    51.32602, 51.3345, 51.34272, 51.35068, 51.35838, 51.36582, 51.373, 
    51.37992, 51.38657, 51.39297, 51.39911, 51.40498, 51.4106, 51.41595, 
    51.42104, 51.42587, 51.43044, 51.43475, 51.43879, 51.44257, 51.44609, 
    51.44935, 51.45235, 51.45509, 51.45756, 51.45977, 51.46171, 51.4634, 
    51.46482, 51.46598, 51.46688, 51.46751, 51.46789, 51.468, 51.46785, 
    51.46743, 51.46675, 51.46582, 51.46461, 51.46315, 51.46142, 51.45943, 
    51.45718, 51.45467, 51.45189, 51.44886, 51.44555, 51.44199, 51.43817, 
    51.43408, 51.42973, 51.42513, 51.42025, 51.41512, 51.40973, 51.40407, 
    51.39816, 51.39198, 51.38554, 51.37884, 51.37188, 51.36466, 51.35718, 
    51.34944, 51.34143, 51.33318, 51.32465, 51.31587, 51.30684, 51.29753, 
    51.28798, 51.27816, 51.26809, 51.25776, 51.24716, 51.23631, 51.2252, 
    51.21384, 51.20222, 51.19034, 51.1782, 51.16581, 51.15316, 51.14026, 
    51.1271, 51.11369, 51.10001, 51.08609, 51.07191, 51.05747, 51.04278, 
    51.02784, 51.01265, 50.9972, 50.98149, 50.96554, 50.94933, 50.93287, 
    50.91616, 50.8992, 50.88199, 50.86452, 50.84681, 50.82885, 50.81063, 
    50.79217, 50.77346, 50.7545, 50.73529, 50.71584, 50.69614, 50.67619, 
    50.65599, 50.63555, 50.61486, 50.59393, 50.57275, 50.55132, 50.52966, 
    50.50774, 50.48559, 50.46319, 50.44056, 50.41767, 50.39455, 50.37119, 
    50.34758, 50.32373, 50.29965, 50.27532, 50.25076, 50.22596, 50.20091, 
    50.17564, 50.15012, 50.12437, 50.09838, 50.07215, 50.0457, 50.019, 
    49.99207, 49.96491, 49.93752, 49.90989, 49.88203, 49.85394, 49.82561, 
    49.79706, 49.76827, 49.73926, 49.71001, 49.68054, 49.65084, 49.62091, 
    49.59076, 49.56037, 49.52976, 49.49893, 49.46787, 49.43658, 49.40508, 
    49.37335, 49.34139, 49.30922, 49.27682, 49.24419, 49.21135, 49.1783, 
    49.14501, 49.11151, 49.07779, 49.04386, 49.0097, 48.97533, 48.94075, 
    48.90594, 48.87092, 48.83569, 48.80024, 48.76458, 48.72871, 48.69262, 
    48.65633, 48.61982, 48.5831, 48.54617, 48.50903, 48.47168, 48.43413, 
    48.39636, 48.35839, 48.32021, 48.28183, 48.24324, 48.20445, 48.16545, 
    48.12625, 48.08685, 48.04724, 48.00743, 47.96742, 47.92721, 47.8868, 
    47.84619, 47.80538,
  43.3274, 43.38415, 43.44075, 43.49721, 43.55353, 43.6097, 43.66572, 
    43.7216, 43.77733, 43.83291, 43.88834, 43.94363, 43.99876, 44.05375, 
    44.10858, 44.16326, 44.21779, 44.27217, 44.3264, 44.38047, 44.43439, 
    44.48815, 44.54176, 44.59521, 44.6485, 44.70164, 44.75462, 44.80744, 
    44.86011, 44.91261, 44.96495, 45.01714, 45.06916, 45.12102, 45.17272, 
    45.22425, 45.27562, 45.32683, 45.37787, 45.42875, 45.47946, 45.53001, 
    45.58038, 45.6306, 45.68064, 45.73051, 45.78021, 45.82975, 45.87911, 
    45.9283, 45.97732, 46.02617, 46.07484, 46.12334, 46.17167, 46.21982, 
    46.26779, 46.31559, 46.36321, 46.41066, 46.45793, 46.50502, 46.55193, 
    46.59866, 46.6452, 46.69157, 46.73776, 46.78376, 46.82959, 46.87523, 
    46.92068, 46.96595, 47.01104, 47.05593, 47.10065, 47.14517, 47.18951, 
    47.23366, 47.27762, 47.32139, 47.36497, 47.40836, 47.45156, 47.49457, 
    47.53738, 47.58001, 47.62244, 47.66467, 47.70671, 47.74855, 47.7902, 
    47.83165, 47.8729, 47.91396, 47.95481, 47.99547, 48.03593, 48.07619, 
    48.11624, 48.1561, 48.19575, 48.2352, 48.27445, 48.31349, 48.35233, 
    48.39096, 48.42939, 48.46761, 48.50562, 48.54343, 48.58103, 48.61842, 
    48.6556, 48.69257, 48.72933, 48.76588, 48.80222, 48.83834, 48.87426, 
    48.90996, 48.94545, 48.98072, 49.01577, 49.05061, 49.08524, 49.11965, 
    49.15384, 49.18781, 49.22157, 49.2551, 49.28842, 49.32151, 49.35439, 
    49.38704, 49.41947, 49.45168, 49.48367, 49.51543, 49.54697, 49.57829, 
    49.60938, 49.64024, 49.67088, 49.70129, 49.73148, 49.76144, 49.79116, 
    49.82066, 49.84994, 49.87898, 49.90779, 49.93637, 49.96472, 49.99283, 
    50.02072, 50.04837, 50.07579, 50.10297, 50.12992, 50.15664, 50.18312, 
    50.20937, 50.23537, 50.26115, 50.28668, 50.31198, 50.33704, 50.36185, 
    50.38644, 50.41078, 50.43488, 50.45874, 50.48236, 50.50574, 50.52888, 
    50.55177, 50.57442, 50.59684, 50.619, 50.64092, 50.6626, 50.68403, 
    50.70522, 50.72617, 50.74686, 50.76731, 50.78751, 50.80747, 50.82718, 
    50.84664, 50.86585, 50.88482, 50.90353, 50.92199, 50.94021, 50.95818, 
    50.97589, 50.99335, 51.01057, 51.02753, 51.04424, 51.0607, 51.0769, 
    51.09285, 51.10855, 51.124, 51.13919, 51.15413, 51.16881, 51.18324, 
    51.19741, 51.21133, 51.22499, 51.2384, 51.25154, 51.26444, 51.27708, 
    51.28946, 51.30158, 51.31345, 51.32506, 51.33641, 51.3475, 51.35833, 
    51.36891, 51.37923, 51.38928, 51.39908, 51.40862, 51.4179, 51.42692, 
    51.43568, 51.44418, 51.45242, 51.4604, 51.46812, 51.47557, 51.48277, 
    51.4897, 51.49638, 51.50279, 51.50894, 51.51483, 51.52046, 51.52583, 
    51.53093, 51.53577, 51.54035, 51.54467, 51.54872, 51.55251, 51.55604, 
    51.55931, 51.56231, 51.56505, 51.56753, 51.56975, 51.5717, 51.57339, 
    51.57481, 51.57598, 51.57688, 51.57751, 51.57789, 51.578, 51.57785, 
    51.57743, 51.57675, 51.57581, 51.57461, 51.57314, 51.57141, 51.56941, 
    51.56716, 51.56464, 51.56186, 51.55881, 51.5555, 51.55193, 51.5481, 
    51.544, 51.53964, 51.53502, 51.53014, 51.52499, 51.51959, 51.51392, 
    51.50799, 51.5018, 51.49534, 51.48862, 51.48165, 51.47441, 51.46692, 
    51.45915, 51.45113, 51.44285, 51.43431, 51.42551, 51.41645, 51.40713, 
    51.39755, 51.38771, 51.37761, 51.36725, 51.35664, 51.34576, 51.33463, 
    51.32324, 51.31159, 51.29968, 51.28752, 51.2751, 51.26242, 51.24949, 
    51.23629, 51.22285, 51.20914, 51.19518, 51.18097, 51.1665, 51.15178, 
    51.1368, 51.12157, 51.10608, 51.09035, 51.07435, 51.05811, 51.04161, 
    51.02486, 51.00786, 50.99061, 50.97311, 50.95535, 50.93735, 50.91909, 
    50.90059, 50.88183, 50.86283, 50.84358, 50.82408, 50.80433, 50.78434, 
    50.76409, 50.7436, 50.72287, 50.70189, 50.68066, 50.65919, 50.63747, 
    50.61551, 50.59331, 50.57086, 50.54817, 50.52523, 50.50206, 50.47864, 
    50.45498, 50.43108, 50.40694, 50.38256, 50.35794, 50.33309, 50.30799, 
    50.28266, 50.25708, 50.23127, 50.20523, 50.17895, 50.15243, 50.12568, 
    50.09869, 50.07147, 50.04401, 50.01632, 49.9884, 49.96025, 49.93186, 
    49.90325, 49.8744, 49.84532, 49.81601, 49.78648, 49.75671, 49.72672, 
    49.6965, 49.66605, 49.63538, 49.60448, 49.57335, 49.542, 49.51043, 
    49.47863, 49.4466, 49.41436, 49.38189, 49.3492, 49.31629, 49.28316, 
    49.24981, 49.21624, 49.18245, 49.14845, 49.11422, 49.07978, 49.04512, 
    49.01024, 48.97515, 48.93985, 48.90433, 48.86859, 48.83265, 48.79649, 
    48.76011, 48.72353, 48.68674, 48.64973, 48.61252, 48.5751, 48.53746, 
    48.49963, 48.46158, 48.42332, 48.38486, 48.3462, 48.30733, 48.26825, 
    48.22897, 48.18949, 48.14981, 48.10992, 48.06983, 48.02954, 47.98905, 
    47.94836, 47.90747,
  43.42155, 43.47839, 43.53508, 43.59163, 43.64803, 43.70429, 43.7604, 
    43.81636, 43.87218, 43.92785, 43.98337, 44.03874, 44.09396, 44.14903, 
    44.20395, 44.25872, 44.31334, 44.36781, 44.42212, 44.47628, 44.53028, 
    44.58413, 44.63783, 44.69136, 44.74475, 44.79797, 44.85104, 44.90395, 
    44.9567, 45.00929, 45.06172, 45.11399, 45.1661, 45.21804, 45.26983, 
    45.32145, 45.37291, 45.4242, 45.47533, 45.52629, 45.57709, 45.62772, 
    45.67819, 45.72849, 45.77861, 45.82857, 45.87836, 45.92798, 45.97743, 
    46.02671, 46.07581, 46.12474, 46.1735, 46.22209, 46.2705, 46.31874, 
    46.3668, 46.41468, 46.46239, 46.50992, 46.55727, 46.60445, 46.65144, 
    46.69825, 46.74489, 46.79134, 46.83761, 46.8837, 46.92961, 46.97533, 
    47.02087, 47.06622, 47.11139, 47.15638, 47.20117, 47.24578, 47.2902, 
    47.33443, 47.37848, 47.42233, 47.46599, 47.50946, 47.55275, 47.59584, 
    47.63873, 47.68143, 47.72395, 47.76626, 47.80838, 47.8503, 47.89203, 
    47.93356, 47.9749, 48.01603, 48.05696, 48.0977, 48.13824, 48.17858, 
    48.21871, 48.25864, 48.29838, 48.33791, 48.37723, 48.41635, 48.45527, 
    48.49398, 48.53248, 48.57078, 48.60887, 48.64675, 48.68443, 48.72189, 
    48.75915, 48.7962, 48.83303, 48.86966, 48.90607, 48.94227, 48.97825, 
    49.01403, 49.04959, 49.08493, 49.12006, 49.15497, 49.18967, 49.22415, 
    49.25841, 49.29245, 49.32628, 49.35989, 49.39327, 49.42644, 49.45938, 
    49.4921, 49.5246, 49.55688, 49.58894, 49.62077, 49.65238, 49.68376, 
    49.71492, 49.74585, 49.77655, 49.80703, 49.83728, 49.8673, 49.89709, 
    49.92666, 49.95599, 49.9851, 50.01397, 50.04261, 50.07102, 50.0992, 
    50.12715, 50.15486, 50.18234, 50.20958, 50.23659, 50.26337, 50.28991, 
    50.31621, 50.34228, 50.3681, 50.3937, 50.41905, 50.44416, 50.46904, 
    50.49368, 50.51807, 50.54223, 50.56614, 50.58982, 50.61325, 50.63644, 
    50.65938, 50.68209, 50.70455, 50.72676, 50.74874, 50.77046, 50.79194, 
    50.81318, 50.83417, 50.85492, 50.87541, 50.89566, 50.91566, 50.93542, 
    50.95492, 50.97418, 50.99319, 51.01194, 51.03045, 51.04871, 51.06672, 
    51.08447, 51.10197, 51.11923, 51.13623, 51.15298, 51.16947, 51.18571, 
    51.20171, 51.21744, 51.23292, 51.24815, 51.26312, 51.27784, 51.2923, 
    51.30651, 51.32046, 51.33415, 51.34759, 51.36077, 51.3737, 51.38636, 
    51.39877, 51.41092, 51.42282, 51.43446, 51.44583, 51.45695, 51.46781, 
    51.47841, 51.48875, 51.49883, 51.50866, 51.51822, 51.52752, 51.53656, 
    51.54534, 51.55386, 51.56212, 51.57012, 51.57785, 51.58533, 51.59254, 
    51.59949, 51.60619, 51.61261, 51.61878, 51.62468, 51.63032, 51.6357, 
    51.64082, 51.64567, 51.65026, 51.65459, 51.65865, 51.66245, 51.66599, 
    51.66926, 51.67228, 51.67502, 51.67751, 51.67973, 51.68168, 51.68338, 
    51.68481, 51.68597, 51.68687, 51.68752, 51.68789, 51.688, 51.68785, 
    51.68743, 51.68675, 51.68581, 51.6846, 51.68313, 51.68139, 51.67939, 
    51.67713, 51.67461, 51.67181, 51.66876, 51.66545, 51.66187, 51.65802, 
    51.65392, 51.64955, 51.64492, 51.64003, 51.63487, 51.62945, 51.62376, 
    51.61782, 51.61161, 51.60514, 51.59841, 51.59142, 51.58416, 51.57665, 
    51.56887, 51.56083, 51.55253, 51.54397, 51.53515, 51.52607, 51.51672, 
    51.50712, 51.49726, 51.48713, 51.47675, 51.46611, 51.45521, 51.44405, 
    51.43263, 51.42096, 51.40902, 51.39683, 51.38438, 51.37167, 51.3587, 
    51.34548, 51.332, 51.31827, 51.30428, 51.29003, 51.27553, 51.26077, 
    51.24576, 51.23049, 51.21497, 51.19919, 51.18316, 51.16688, 51.15034, 
    51.13356, 51.11652, 51.09922, 51.08168, 51.06388, 51.04584, 51.02754, 
    51.00899, 50.9902, 50.97115, 50.95185, 50.93231, 50.91251, 50.89248, 
    50.87218, 50.85165, 50.83087, 50.80984, 50.78856, 50.76704, 50.74528, 
    50.72327, 50.70101, 50.67851, 50.65577, 50.63279, 50.60956, 50.58609, 
    50.56237, 50.53842, 50.51423, 50.4898, 50.46512, 50.44021, 50.41505, 
    50.38966, 50.36404, 50.33817, 50.31207, 50.28572, 50.25915, 50.23234, 
    50.20529, 50.17801, 50.15049, 50.12274, 50.09476, 50.06654, 50.0381, 
    50.00942, 49.98051, 49.95137, 49.922, 49.8924, 49.86257, 49.83251, 
    49.80222, 49.77171, 49.74097, 49.71, 49.67881, 49.64739, 49.61575, 
    49.58389, 49.55179, 49.51948, 49.48694, 49.45419, 49.42121, 49.388, 
    49.35458, 49.32095, 49.28709, 49.25301, 49.21871, 49.1842, 49.14946, 
    49.11452, 49.07935, 49.04398, 49.00838, 48.97258, 48.93655, 48.90032, 
    48.86388, 48.82722, 48.79035, 48.75327, 48.71598, 48.67848, 48.64077, 
    48.60286, 48.56474, 48.52641, 48.48787, 48.44912, 48.41018, 48.37102, 
    48.33167, 48.29211, 48.25234, 48.21238, 48.17221, 48.13184, 48.09127, 
    48.0505, 48.00954,
  43.51566, 43.57258, 43.62936, 43.686, 43.74249, 43.79883, 43.85503, 
    43.91108, 43.96698, 44.02274, 44.07834, 44.1338, 44.18911, 44.24427, 
    44.29927, 44.35413, 44.40884, 44.46339, 44.51779, 44.57203, 44.62613, 
    44.68006, 44.73384, 44.78747, 44.84094, 44.89425, 44.94741, 45.0004, 
    45.05324, 45.10592, 45.15844, 45.21079, 45.26299, 45.31502, 45.36689, 
    45.4186, 45.47015, 45.52153, 45.57274, 45.62379, 45.67468, 45.7254, 
    45.77595, 45.82633, 45.87654, 45.92659, 45.97647, 46.02617, 46.07571, 
    46.12507, 46.17426, 46.22328, 46.27213, 46.3208, 46.36929, 46.41761, 
    46.46576, 46.51373, 46.56152, 46.60914, 46.65658, 46.70384, 46.75092, 
    46.79782, 46.84454, 46.89107, 46.93743, 46.9836, 47.02959, 47.0754, 
    47.12102, 47.16646, 47.21171, 47.25677, 47.30165, 47.34635, 47.39085, 
    47.43517, 47.47929, 47.52323, 47.56697, 47.61053, 47.6539, 47.69707, 
    47.74004, 47.78283, 47.82542, 47.86782, 47.91002, 47.95202, 47.99383, 
    48.03544, 48.07685, 48.11807, 48.15909, 48.1999, 48.24052, 48.28094, 
    48.32115, 48.36116, 48.40097, 48.44058, 48.47998, 48.51918, 48.55817, 
    48.59696, 48.63554, 48.67392, 48.71209, 48.75005, 48.7878, 48.82534, 
    48.86267, 48.89979, 48.9367, 48.9734, 49.00989, 49.04616, 49.08222, 
    49.11807, 49.1537, 49.18912, 49.22432, 49.25931, 49.29408, 49.32863, 
    49.36296, 49.39708, 49.43097, 49.46465, 49.4981, 49.53134, 49.56435, 
    49.59715, 49.62972, 49.66206, 49.69419, 49.72609, 49.75776, 49.78921, 
    49.82043, 49.85143, 49.8822, 49.91274, 49.94306, 49.97314, 50.003, 
    50.03263, 50.06203, 50.0912, 50.12014, 50.14884, 50.17731, 50.20555, 
    50.23356, 50.26133, 50.28887, 50.31618, 50.34325, 50.37008, 50.39668, 
    50.42304, 50.44917, 50.47505, 50.5007, 50.52611, 50.55128, 50.57621, 
    50.6009, 50.62535, 50.64956, 50.67353, 50.69726, 50.72074, 50.74398, 
    50.76698, 50.78974, 50.81225, 50.83451, 50.85654, 50.87831, 50.89985, 
    50.92113, 50.94217, 50.96296, 50.9835, 51.0038, 51.02385, 51.04365, 
    51.0632, 51.0825, 51.10155, 51.12035, 51.1389, 51.1572, 51.17525, 
    51.19305, 51.21059, 51.22788, 51.24492, 51.26171, 51.27824, 51.29453, 
    51.31055, 51.32632, 51.34184, 51.35711, 51.37211, 51.38686, 51.40136, 
    51.4156, 51.42958, 51.44331, 51.45678, 51.46999, 51.48295, 51.49564, 
    51.50808, 51.52026, 51.53218, 51.54385, 51.55525, 51.5664, 51.57729, 
    51.58791, 51.59827, 51.60838, 51.61823, 51.62781, 51.63713, 51.6462, 
    51.655, 51.66354, 51.67182, 51.67984, 51.68759, 51.69508, 51.70231, 
    51.70928, 51.71599, 51.72243, 51.72861, 51.73453, 51.74018, 51.74557, 
    51.7507, 51.75557, 51.76017, 51.76451, 51.76858, 51.77239, 51.77594, 
    51.77922, 51.78224, 51.78499, 51.78748, 51.78971, 51.79167, 51.79337, 
    51.7948, 51.79597, 51.79687, 51.79751, 51.79789, 51.798, 51.79785, 
    51.79743, 51.79675, 51.7958, 51.79459, 51.79311, 51.79137, 51.78937, 
    51.78711, 51.78457, 51.78178, 51.77872, 51.77539, 51.7718, 51.76795, 
    51.76384, 51.75946, 51.75481, 51.74991, 51.74474, 51.73931, 51.73361, 
    51.72765, 51.72143, 51.71495, 51.7082, 51.70119, 51.69392, 51.68638, 
    51.67859, 51.67052, 51.6622, 51.65363, 51.64478, 51.63568, 51.62631, 
    51.61669, 51.6068, 51.59665, 51.58625, 51.57558, 51.56465, 51.55347, 
    51.54202, 51.53032, 51.51835, 51.50613, 51.49365, 51.48092, 51.46792, 
    51.45467, 51.44115, 51.42739, 51.41336, 51.39908, 51.38455, 51.36975, 
    51.35471, 51.33941, 51.32384, 51.30803, 51.29197, 51.27565, 51.25907, 
    51.24224, 51.22517, 51.20783, 51.19025, 51.17241, 51.15432, 51.13598, 
    51.11739, 51.09855, 51.07946, 51.06012, 51.04053, 51.02069, 51.00061, 
    50.98027, 50.95969, 50.93886, 50.91778, 50.89646, 50.87489, 50.85307, 
    50.83101, 50.8087, 50.78616, 50.76336, 50.74033, 50.71704, 50.69352, 
    50.66975, 50.64575, 50.6215, 50.59701, 50.57228, 50.54731, 50.52211, 
    50.49666, 50.47097, 50.44505, 50.41888, 50.39249, 50.36585, 50.33898, 
    50.31187, 50.28453, 50.25695, 50.22915, 50.2011, 50.17282, 50.14431, 
    50.11557, 50.0866, 50.0574, 50.02796, 49.99829, 49.9684, 49.93828, 
    49.90793, 49.87735, 49.84654, 49.81551, 49.78425, 49.75277, 49.72105, 
    49.68912, 49.65696, 49.62458, 49.59198, 49.55915, 49.5261, 49.49283, 
    49.45934, 49.42562, 49.39169, 49.35754, 49.32318, 49.28859, 49.25379, 
    49.21877, 49.18353, 49.14808, 49.11242, 49.07653, 49.04044, 49.00413, 
    48.96761, 48.93088, 48.89393, 48.85678, 48.81941, 48.78184, 48.74405, 
    48.70606, 48.66786, 48.62946, 48.59084, 48.55202, 48.51299, 48.47376, 
    48.43433, 48.39469, 48.35485, 48.3148, 48.27456, 48.23411, 48.19346, 
    48.15261, 48.11156,
  43.60971, 43.66672, 43.72359, 43.78031, 43.83688, 43.89331, 43.9496, 
    44.00574, 44.06173, 44.11757, 44.17326, 44.22881, 44.28421, 44.33945, 
    44.39455, 44.44949, 44.50428, 44.55892, 44.61341, 44.66774, 44.72192, 
    44.77594, 44.82981, 44.88353, 44.93708, 44.99048, 45.04372, 45.09681, 
    45.14973, 45.2025, 45.2551, 45.30754, 45.35983, 45.41195, 45.46391, 
    45.51571, 45.56734, 45.6188, 45.67011, 45.72124, 45.77222, 45.82302, 
    45.87366, 45.92413, 45.97443, 46.02456, 46.07452, 46.12432, 46.17394, 
    46.22339, 46.27267, 46.32177, 46.3707, 46.41946, 46.46804, 46.51645, 
    46.56468, 46.61274, 46.66062, 46.70832, 46.75584, 46.80318, 46.85035, 
    46.89734, 46.94414, 46.99076, 47.0372, 47.08346, 47.12954, 47.17543, 
    47.22113, 47.26665, 47.31199, 47.35714, 47.4021, 47.44688, 47.49147, 
    47.53587, 47.58007, 47.62409, 47.66792, 47.71156, 47.755, 47.79826, 
    47.84132, 47.88419, 47.92686, 47.96934, 48.01162, 48.05371, 48.0956, 
    48.13729, 48.17878, 48.22008, 48.26117, 48.30207, 48.34277, 48.38326, 
    48.42356, 48.46365, 48.50354, 48.54322, 48.5827, 48.62198, 48.66105, 
    48.69992, 48.73857, 48.77703, 48.81527, 48.85331, 48.89114, 48.92875, 
    48.96616, 49.00336, 49.04034, 49.07712, 49.11368, 49.15003, 49.18616, 
    49.22209, 49.25779, 49.29329, 49.32856, 49.36362, 49.39846, 49.43308, 
    49.46749, 49.50167, 49.53564, 49.56939, 49.60292, 49.63622, 49.66931, 
    49.70217, 49.73481, 49.76722, 49.79942, 49.83138, 49.86312, 49.89464, 
    49.92593, 49.957, 49.98783, 50.01844, 50.04882, 50.07897, 50.10889, 
    50.13859, 50.16805, 50.19728, 50.22628, 50.25505, 50.28358, 50.31189, 
    50.33995, 50.36779, 50.39539, 50.42276, 50.44989, 50.47678, 50.50344, 
    50.52985, 50.55604, 50.58198, 50.60769, 50.63315, 50.65838, 50.68337, 
    50.70811, 50.73262, 50.75689, 50.78091, 50.80469, 50.82823, 50.85152, 
    50.87457, 50.89738, 50.91994, 50.94226, 50.96433, 50.98616, 51.00774, 
    51.02907, 51.05016, 51.071, 51.09159, 51.11193, 51.13202, 51.15187, 
    51.17146, 51.19081, 51.2099, 51.22875, 51.24734, 51.26569, 51.28378, 
    51.30161, 51.3192, 51.33653, 51.35361, 51.37044, 51.38701, 51.40333, 
    51.4194, 51.4352, 51.45076, 51.46606, 51.4811, 51.49588, 51.51041, 
    51.52469, 51.5387, 51.55246, 51.56596, 51.57921, 51.59219, 51.60492, 
    51.61739, 51.6296, 51.64155, 51.65324, 51.66467, 51.67585, 51.68676, 
    51.69741, 51.7078, 51.71793, 51.72779, 51.7374, 51.74675, 51.75583, 
    51.76466, 51.77322, 51.78152, 51.78955, 51.79733, 51.80484, 51.81208, 
    51.81907, 51.82579, 51.83225, 51.83844, 51.84438, 51.85004, 51.85545, 
    51.86059, 51.86547, 51.87008, 51.87442, 51.87851, 51.88233, 51.88588, 
    51.88917, 51.8922, 51.89496, 51.89746, 51.89968, 51.90165, 51.90335, 
    51.90479, 51.90596, 51.90687, 51.90751, 51.90789, 51.908, 51.90784, 
    51.90743, 51.90674, 51.9058, 51.90458, 51.9031, 51.90136, 51.89935, 
    51.89708, 51.89454, 51.89174, 51.88867, 51.88534, 51.88174, 51.87788, 
    51.87376, 51.86937, 51.86471, 51.85979, 51.85461, 51.84917, 51.84346, 
    51.83748, 51.83125, 51.82475, 51.81798, 51.81096, 51.80367, 51.79611, 
    51.7883, 51.78022, 51.77188, 51.76328, 51.75441, 51.74529, 51.7359, 
    51.72625, 51.71634, 51.70617, 51.69574, 51.68505, 51.6741, 51.66288, 
    51.65141, 51.63968, 51.62769, 51.61544, 51.60292, 51.59016, 51.57713, 
    51.56385, 51.5503, 51.5365, 51.52245, 51.50813, 51.49356, 51.47874, 
    51.46365, 51.44831, 51.43272, 51.41687, 51.40076, 51.38441, 51.36779, 
    51.35093, 51.33381, 51.31643, 51.29881, 51.28093, 51.2628, 51.24442, 
    51.22578, 51.2069, 51.18776, 51.16838, 51.14875, 51.12886, 51.10873, 
    51.08834, 51.06771, 51.04684, 51.02571, 51.00434, 50.98272, 50.96085, 
    50.93874, 50.91639, 50.89379, 50.87094, 50.84785, 50.82452, 50.80094, 
    50.77712, 50.75306, 50.72876, 50.70422, 50.67943, 50.65441, 50.62914, 
    50.60364, 50.57789, 50.55191, 50.52569, 50.49923, 50.47254, 50.44561, 
    50.41844, 50.39104, 50.3634, 50.33553, 50.30743, 50.27909, 50.25051, 
    50.22171, 50.19267, 50.16341, 50.13391, 50.10418, 50.07422, 50.04403, 
    50.01361, 49.98297, 49.9521, 49.921, 49.88967, 49.85812, 49.82634, 
    49.79434, 49.76211, 49.72966, 49.69698, 49.66409, 49.63097, 49.59763, 
    49.56406, 49.53028, 49.49628, 49.46206, 49.42762, 49.39296, 49.35809, 
    49.32299, 49.28769, 49.25216, 49.21642, 49.18047, 49.14429, 49.10791, 
    49.07132, 49.03451, 48.99749, 48.96026, 48.92282, 48.88517, 48.84731, 
    48.80924, 48.77096, 48.73248, 48.69378, 48.65488, 48.61578, 48.57647, 
    48.53696, 48.49724, 48.45732, 48.4172, 48.37687, 48.33634, 48.29562, 
    48.25469, 48.21356,
  43.70371, 43.7608, 43.81776, 43.87457, 43.93123, 43.98775, 44.04412, 
    44.10034, 44.15642, 44.21235, 44.26814, 44.32376, 44.37925, 44.43458, 
    44.48977, 44.5448, 44.59968, 44.6544, 44.70898, 44.7634, 44.81767, 
    44.87178, 44.92574, 44.97953, 45.03318, 45.08667, 45.14, 45.19316, 
    45.24618, 45.29903, 45.35172, 45.40425, 45.45662, 45.50883, 45.56088, 
    45.61276, 45.66448, 45.71603, 45.76743, 45.81865, 45.86971, 45.9206, 
    45.97132, 46.02188, 46.07227, 46.12249, 46.17254, 46.22242, 46.27213, 
    46.32166, 46.37103, 46.42022, 46.46923, 46.51808, 46.56675, 46.61524, 
    46.66356, 46.7117, 46.75967, 46.80745, 46.85506, 46.90249, 46.94974, 
    46.99681, 47.0437, 47.09041, 47.13694, 47.18328, 47.22944, 47.27541, 
    47.32121, 47.36681, 47.41223, 47.45747, 47.50251, 47.54737, 47.59204, 
    47.63652, 47.68082, 47.72492, 47.76883, 47.81255, 47.85608, 47.89942, 
    47.94256, 47.98551, 48.02827, 48.07082, 48.11319, 48.15536, 48.19733, 
    48.2391, 48.28068, 48.32205, 48.36323, 48.40421, 48.44498, 48.48556, 
    48.52593, 48.5661, 48.60607, 48.64584, 48.68539, 48.72475, 48.7639, 
    48.80285, 48.84158, 48.88011, 48.91843, 48.95655, 48.99445, 49.03214, 
    49.06963, 49.1069, 49.14396, 49.18081, 49.21745, 49.25387, 49.29008, 
    49.32608, 49.36186, 49.39742, 49.43277, 49.4679, 49.50282, 49.53751, 
    49.57199, 49.60625, 49.64029, 49.67411, 49.7077, 49.74108, 49.77423, 
    49.80717, 49.83987, 49.87236, 49.90462, 49.93666, 49.96847, 50.00005, 
    50.03141, 50.06254, 50.09344, 50.12412, 50.15456, 50.18478, 50.21477, 
    50.24453, 50.27405, 50.30335, 50.33241, 50.36124, 50.38984, 50.41821, 
    50.44633, 50.47423, 50.50189, 50.52932, 50.55651, 50.58346, 50.61018, 
    50.63665, 50.6629, 50.6889, 50.71466, 50.74018, 50.76547, 50.79051, 
    50.81532, 50.83988, 50.8642, 50.88827, 50.91211, 50.9357, 50.95905, 
    50.98215, 51.00501, 51.02762, 51.04999, 51.07211, 51.09399, 51.11562, 
    51.137, 51.15813, 51.17902, 51.19966, 51.22005, 51.24019, 51.26008, 
    51.27972, 51.29911, 51.31825, 51.33714, 51.35578, 51.37416, 51.39229, 
    51.41018, 51.4278, 51.44518, 51.4623, 51.47916, 51.49577, 51.51213, 
    51.52823, 51.54408, 51.55967, 51.575, 51.59008, 51.6049, 51.61946, 
    51.63377, 51.64782, 51.66161, 51.67515, 51.68842, 51.70144, 51.7142, 
    51.72669, 51.73893, 51.75091, 51.76263, 51.77409, 51.78529, 51.79623, 
    51.8069, 51.81732, 51.82747, 51.83736, 51.84699, 51.85636, 51.86547, 
    51.87431, 51.88289, 51.89121, 51.89927, 51.90706, 51.91459, 51.92185, 
    51.92886, 51.93559, 51.94207, 51.94828, 51.95422, 51.9599, 51.96532, 
    51.97047, 51.97536, 51.97998, 51.98434, 51.98844, 51.99227, 51.99583, 
    51.99913, 52.00216, 52.00493, 52.00743, 52.00967, 52.01164, 52.01334, 
    52.01478, 52.01596, 52.01687, 52.01751, 52.01789, 52.018, 52.01785, 
    52.01743, 52.01674, 52.01579, 52.01457, 52.01309, 52.01134, 52.00933, 
    52.00705, 52.00451, 52.0017, 51.99862, 51.99529, 51.99168, 51.98781, 
    51.98367, 51.97927, 51.97461, 51.96968, 51.96448, 51.95902, 51.9533, 
    51.94731, 51.94106, 51.93454, 51.92776, 51.92072, 51.91341, 51.90584, 
    51.89801, 51.88991, 51.88155, 51.87293, 51.86404, 51.8549, 51.84549, 
    51.83582, 51.82588, 51.81569, 51.80523, 51.79451, 51.78354, 51.77229, 
    51.7608, 51.74903, 51.73701, 51.72474, 51.7122, 51.6994, 51.68634, 
    51.67302, 51.65945, 51.64561, 51.63153, 51.61718, 51.60257, 51.58771, 
    51.57259, 51.55722, 51.54159, 51.5257, 51.50956, 51.49316, 51.47651, 
    51.4596, 51.44244, 51.42503, 51.40736, 51.38944, 51.37127, 51.35284, 
    51.33417, 51.31524, 51.29606, 51.27663, 51.25695, 51.23702, 51.21684, 
    51.19641, 51.17574, 51.15481, 51.13363, 51.11221, 51.09055, 51.06863, 
    51.04647, 51.02406, 51.00141, 50.97851, 50.95537, 50.93198, 50.90835, 
    50.88448, 50.86036, 50.83601, 50.81141, 50.78657, 50.76149, 50.73616, 
    50.7106, 50.6848, 50.65876, 50.63248, 50.60597, 50.57921, 50.55222, 
    50.52499, 50.49753, 50.46983, 50.4419, 50.41373, 50.38533, 50.3567, 
    50.32783, 50.29873, 50.2694, 50.23983, 50.21004, 50.18002, 50.14977, 
    50.11928, 50.08857, 50.05763, 50.02646, 49.99507, 49.96345, 49.9316, 
    49.89953, 49.86724, 49.83472, 49.80197, 49.769, 49.73582, 49.7024, 
    49.66877, 49.63492, 49.60085, 49.56655, 49.53204, 49.49731, 49.46236, 
    49.42719, 49.39181, 49.35621, 49.3204, 49.28437, 49.24813, 49.21167, 
    49.175, 49.13811, 49.10102, 49.06371, 49.0262, 48.98847, 48.95053, 
    48.91238, 48.87403, 48.83547, 48.7967, 48.75772, 48.71854, 48.67915, 
    48.63956, 48.59976, 48.55976, 48.51956, 48.47915, 48.43855, 48.39774, 
    48.35673, 48.31552,
  43.79765, 43.85483, 43.91187, 43.96877, 44.02552, 44.08212, 44.13858, 
    44.1949, 44.25106, 44.30708, 44.36295, 44.41867, 44.47424, 44.52966, 
    44.58493, 44.64005, 44.69502, 44.74984, 44.8045, 44.859, 44.91336, 
    44.96756, 45.0216, 45.07549, 45.12922, 45.1828, 45.23621, 45.28947, 
    45.34257, 45.39551, 45.44829, 45.50091, 45.55337, 45.60567, 45.6578, 
    45.70977, 45.76158, 45.81322, 45.8647, 45.91601, 45.96716, 46.01814, 
    46.06895, 46.11959, 46.17007, 46.22037, 46.27051, 46.32047, 46.37027, 
    46.41989, 46.46934, 46.51862, 46.56773, 46.61666, 46.66541, 46.71399, 
    46.7624, 46.81062, 46.85868, 46.90655, 46.95424, 47.00176, 47.0491, 
    47.09625, 47.14322, 47.19002, 47.23663, 47.28306, 47.3293, 47.37536, 
    47.42124, 47.46693, 47.51244, 47.55775, 47.60288, 47.64783, 47.69258, 
    47.73715, 47.78152, 47.82571, 47.86971, 47.91351, 47.95712, 48.00054, 
    48.04377, 48.0868, 48.12963, 48.17228, 48.21472, 48.25697, 48.29903, 
    48.34088, 48.38254, 48.42399, 48.46525, 48.50631, 48.54716, 48.58782, 
    48.62827, 48.66853, 48.70857, 48.74842, 48.78806, 48.82749, 48.86672, 
    48.90574, 48.94455, 48.98316, 49.02156, 49.05975, 49.09773, 49.13551, 
    49.17307, 49.21041, 49.24755, 49.28448, 49.32119, 49.35769, 49.39397, 
    49.43004, 49.4659, 49.50154, 49.53696, 49.57216, 49.60715, 49.64192, 
    49.67647, 49.7108, 49.74491, 49.7788, 49.81247, 49.84592, 49.87914, 
    49.91214, 49.94492, 49.97747, 50.0098, 50.04191, 50.07379, 50.10544, 
    50.13686, 50.16806, 50.19903, 50.22977, 50.26029, 50.29057, 50.32063, 
    50.35044, 50.38004, 50.4094, 50.43852, 50.46742, 50.49608, 50.52451, 
    50.5527, 50.58066, 50.60838, 50.63586, 50.66312, 50.69013, 50.7169, 
    50.74344, 50.76974, 50.7958, 50.82162, 50.8472, 50.87254, 50.89764, 
    50.9225, 50.94712, 50.97149, 50.99562, 51.01951, 51.04316, 51.06656, 
    51.08971, 51.11263, 51.13529, 51.15771, 51.17988, 51.20181, 51.22349, 
    51.24492, 51.2661, 51.28704, 51.30772, 51.32816, 51.34835, 51.36829, 
    51.38797, 51.40741, 51.42659, 51.44552, 51.4642, 51.48263, 51.5008, 
    51.51873, 51.5364, 51.55381, 51.57097, 51.58788, 51.60453, 51.62092, 
    51.63706, 51.65294, 51.66857, 51.68394, 51.69905, 51.71391, 51.72851, 
    51.74285, 51.75694, 51.77076, 51.78432, 51.79763, 51.81068, 51.82347, 
    51.83599, 51.84826, 51.86027, 51.87202, 51.8835, 51.89473, 51.90569, 
    51.91639, 51.92683, 51.93701, 51.94693, 51.95658, 51.96597, 51.9751, 
    51.98396, 51.99257, 52.0009, 52.00898, 52.01679, 52.02434, 52.03162, 
    52.03864, 52.04539, 52.05188, 52.05811, 52.06407, 52.06976, 52.0752, 
    52.08036, 52.08526, 52.08989, 52.09426, 52.09837, 52.1022, 52.10577, 
    52.10908, 52.11212, 52.11489, 52.1174, 52.11965, 52.12162, 52.12333, 
    52.12477, 52.12595, 52.12687, 52.12751, 52.12789, 52.128, 52.12785, 
    52.12743, 52.12674, 52.12579, 52.12457, 52.12308, 52.12133, 52.11931, 
    52.11702, 52.11448, 52.11166, 52.10858, 52.10523, 52.10162, 52.09774, 
    52.09359, 52.08918, 52.0845, 52.07956, 52.07435, 52.06888, 52.06314, 
    52.05714, 52.05087, 52.04434, 52.03755, 52.03049, 52.02316, 52.01557, 
    52.00772, 51.9996, 51.99122, 51.98258, 51.97367, 51.9645, 51.95507, 
    51.94538, 51.93542, 51.9252, 51.91472, 51.90397, 51.89297, 51.8817, 
    51.87017, 51.85839, 51.84634, 51.83403, 51.82146, 51.80863, 51.79554, 
    51.7822, 51.76859, 51.75472, 51.7406, 51.72622, 51.71158, 51.69668, 
    51.68153, 51.66611, 51.65045, 51.63453, 51.61834, 51.60191, 51.58522, 
    51.56827, 51.55107, 51.53362, 51.51591, 51.49795, 51.47973, 51.46127, 
    51.44254, 51.42357, 51.40435, 51.38487, 51.36515, 51.34517, 51.32494, 
    51.30447, 51.28374, 51.26277, 51.24155, 51.22008, 51.19836, 51.17639, 
    51.15418, 51.13172, 51.10902, 51.08607, 51.06287, 51.03943, 51.01575, 
    50.99183, 50.96766, 50.94324, 50.91859, 50.89369, 50.86855, 50.84317, 
    50.81755, 50.79169, 50.7656, 50.73926, 50.71268, 50.68587, 50.65882, 
    50.63153, 50.60401, 50.57625, 50.54826, 50.52002, 50.49156, 50.46286, 
    50.43393, 50.40477, 50.37537, 50.34575, 50.31588, 50.2858, 50.25548, 
    50.22493, 50.19415, 50.16314, 50.13191, 50.10045, 50.06876, 50.03685, 
    50.0047, 49.97234, 49.93975, 49.90694, 49.8739, 49.84064, 49.80716, 
    49.77345, 49.73953, 49.70538, 49.67102, 49.63643, 49.60163, 49.56661, 
    49.53137, 49.49591, 49.46024, 49.42435, 49.38825, 49.35193, 49.3154, 
    49.27865, 49.24169, 49.20452, 49.16714, 49.12954, 49.09174, 49.05373, 
    49.0155, 48.97707, 48.93843, 48.89958, 48.86053, 48.82127, 48.7818, 
    48.74213, 48.70225, 48.66217, 48.62189, 48.5814, 48.54072, 48.49983, 
    48.45874, 48.41745,
  43.89154, 43.94881, 44.00594, 44.06292, 44.11975, 44.17645, 44.233, 
    44.2894, 44.34565, 44.40176, 44.45771, 44.51352, 44.56918, 44.62469, 
    44.68005, 44.73525, 44.79031, 44.84521, 44.89996, 44.95456, 45.009, 
    45.06329, 45.11742, 45.1714, 45.22522, 45.27888, 45.33238, 45.38573, 
    45.43892, 45.49195, 45.54482, 45.59752, 45.65007, 45.70245, 45.75467, 
    45.80673, 45.85862, 45.91035, 45.96192, 46.01332, 46.06455, 46.11562, 
    46.16652, 46.21725, 46.26781, 46.31821, 46.36843, 46.41848, 46.46836, 
    46.51808, 46.56762, 46.61698, 46.66617, 46.71519, 46.76403, 46.8127, 
    46.86119, 46.9095, 46.95764, 47.0056, 47.05338, 47.10098, 47.1484, 
    47.19564, 47.24271, 47.28959, 47.33628, 47.38279, 47.42912, 47.47527, 
    47.52123, 47.56701, 47.6126, 47.658, 47.70322, 47.74825, 47.79308, 
    47.83773, 47.88219, 47.92646, 47.97054, 48.01443, 48.05812, 48.10163, 
    48.14494, 48.18805, 48.23097, 48.27369, 48.31622, 48.35855, 48.40069, 
    48.44262, 48.48436, 48.5259, 48.56724, 48.60838, 48.64931, 48.69005, 
    48.73058, 48.77092, 48.81104, 48.85097, 48.89069, 48.9302, 48.96951, 
    49.00861, 49.0475, 49.08619, 49.12466, 49.16293, 49.20099, 49.23883, 
    49.27647, 49.3139, 49.35111, 49.38811, 49.4249, 49.46148, 49.49784, 
    49.53398, 49.56991, 49.60562, 49.64112, 49.6764, 49.71146, 49.7463, 
    49.78092, 49.81533, 49.84951, 49.88347, 49.91721, 49.95073, 49.98402, 
    50.0171, 50.04995, 50.08257, 50.11497, 50.14714, 50.17909, 50.21081, 
    50.2423, 50.27357, 50.3046, 50.33541, 50.36599, 50.39634, 50.42646, 
    50.45635, 50.486, 50.51543, 50.54462, 50.57357, 50.6023, 50.63079, 
    50.65905, 50.68707, 50.71485, 50.7424, 50.76971, 50.79678, 50.82362, 
    50.85021, 50.87657, 50.90269, 50.92857, 50.95421, 50.97961, 51.00476, 
    51.02967, 51.05435, 51.07878, 51.10297, 51.12691, 51.1506, 51.17406, 
    51.19727, 51.22023, 51.24295, 51.26542, 51.28764, 51.30962, 51.33135, 
    51.35283, 51.37406, 51.39505, 51.41578, 51.43626, 51.4565, 51.47648, 
    51.49621, 51.51569, 51.53492, 51.5539, 51.57262, 51.59109, 51.60931, 
    51.62727, 51.64499, 51.66244, 51.67964, 51.69658, 51.71328, 51.72971, 
    51.74588, 51.76181, 51.77747, 51.79288, 51.80803, 51.82292, 51.83755, 
    51.85193, 51.86604, 51.8799, 51.8935, 51.90684, 51.91991, 51.93273, 
    51.94529, 51.95759, 51.96962, 51.9814, 51.99291, 52.00417, 52.01516, 
    52.02588, 52.03635, 52.04655, 52.05649, 52.06617, 52.07558, 52.08473, 
    52.09362, 52.10224, 52.1106, 52.11869, 52.12652, 52.13409, 52.14139, 
    52.14842, 52.15519, 52.1617, 52.16794, 52.17391, 52.17962, 52.18507, 
    52.19024, 52.19516, 52.1998, 52.20418, 52.20829, 52.21214, 52.21572, 
    52.21904, 52.22208, 52.22486, 52.22738, 52.22963, 52.23161, 52.23332, 
    52.23477, 52.23595, 52.23686, 52.23751, 52.23789, 52.238, 52.23785, 
    52.23742, 52.23674, 52.23578, 52.23456, 52.23307, 52.23131, 52.22929, 
    52.227, 52.22444, 52.22162, 52.21853, 52.21517, 52.21155, 52.20766, 
    52.20351, 52.19909, 52.1944, 52.18944, 52.18422, 52.17874, 52.17299, 
    52.16697, 52.16069, 52.15414, 52.14733, 52.14025, 52.13291, 52.1253, 
    52.11743, 52.10929, 52.10089, 52.09223, 52.0833, 52.07411, 52.06466, 
    52.05494, 52.04495, 52.03471, 52.0242, 52.01344, 52.0024, 51.99111, 
    51.97955, 51.96774, 51.95566, 51.94332, 51.93072, 51.91786, 51.90474, 
    51.89137, 51.87773, 51.86383, 51.84967, 51.83525, 51.82058, 51.80565, 
    51.79046, 51.77501, 51.7593, 51.74334, 51.72713, 51.71065, 51.69392, 
    51.67694, 51.65969, 51.6422, 51.62445, 51.60645, 51.58819, 51.56968, 
    51.55091, 51.5319, 51.51263, 51.49311, 51.47334, 51.45331, 51.43304, 
    51.41252, 51.39174, 51.37072, 51.34945, 51.32793, 51.30616, 51.28415, 
    51.26188, 51.23937, 51.21662, 51.19361, 51.17036, 51.14687, 51.12313, 
    51.09916, 51.07493, 51.05046, 51.02575, 51.0008, 50.97561, 50.95017, 
    50.92449, 50.89857, 50.87242, 50.84602, 50.81939, 50.79251, 50.7654, 
    50.73805, 50.71047, 50.68265, 50.65459, 50.6263, 50.59777, 50.56901, 
    50.54002, 50.51079, 50.48133, 50.45163, 50.42171, 50.39156, 50.36117, 
    50.33055, 50.29971, 50.26864, 50.23734, 50.20581, 50.17405, 50.14207, 
    50.10986, 50.07742, 50.04476, 50.01188, 49.97877, 49.94544, 49.91189, 
    49.87811, 49.84412, 49.8099, 49.77546, 49.7408, 49.70592, 49.67083, 
    49.63552, 49.59999, 49.56424, 49.52828, 49.4921, 49.45571, 49.4191, 
    49.38227, 49.34524, 49.30799, 49.27053, 49.23286, 49.19498, 49.15689, 
    49.11859, 49.08008, 49.04136, 49.00243, 48.9633, 48.92396, 48.88441, 
    48.84467, 48.80471, 48.76455, 48.72419, 48.68362, 48.64285, 48.60188, 
    48.56071, 48.51934,
  43.98537, 44.04272, 44.09994, 44.15701, 44.21394, 44.27072, 44.32735, 
    44.38384, 44.44018, 44.49638, 44.55242, 44.60832, 44.66407, 44.71966, 
    44.77511, 44.8304, 44.88555, 44.94054, 44.99538, 45.05006, 45.10459, 
    45.15897, 45.21319, 45.26725, 45.32116, 45.37491, 45.4285, 45.48194, 
    45.53521, 45.58833, 45.64128, 45.69408, 45.74672, 45.79919, 45.8515, 
    45.90364, 45.95562, 46.00744, 46.0591, 46.11058, 46.1619, 46.21306, 
    46.26405, 46.31487, 46.36552, 46.416, 46.46631, 46.51645, 46.56642, 
    46.61621, 46.66584, 46.71529, 46.76457, 46.81367, 46.86261, 46.91136, 
    46.95994, 47.00834, 47.05656, 47.10461, 47.15248, 47.20016, 47.24767, 
    47.295, 47.34214, 47.38911, 47.43589, 47.48249, 47.52891, 47.57514, 
    47.62119, 47.66705, 47.71272, 47.75821, 47.80351, 47.84862, 47.89355, 
    47.93828, 47.98283, 48.02718, 48.07134, 48.11531, 48.15909, 48.20267, 
    48.24607, 48.28926, 48.33227, 48.37508, 48.41769, 48.4601, 48.50232, 
    48.54433, 48.58615, 48.62777, 48.66919, 48.71041, 48.75143, 48.79225, 
    48.83286, 48.87328, 48.91348, 48.95348, 48.99328, 49.03288, 49.07226, 
    49.11144, 49.15041, 49.18917, 49.22773, 49.26608, 49.30421, 49.34214, 
    49.37985, 49.41735, 49.45465, 49.49173, 49.52859, 49.56524, 49.60167, 
    49.63789, 49.6739, 49.70969, 49.74525, 49.78061, 49.81574, 49.85065, 
    49.88535, 49.91983, 49.95408, 49.98812, 50.02193, 50.05552, 50.08888, 
    50.12203, 50.15495, 50.18764, 50.22011, 50.25235, 50.28437, 50.31615, 
    50.34772, 50.37905, 50.41016, 50.44103, 50.47168, 50.50209, 50.53228, 
    50.56223, 50.59195, 50.62144, 50.6507, 50.67971, 50.7085, 50.73706, 
    50.76537, 50.79346, 50.8213, 50.84891, 50.87628, 50.90342, 50.93031, 
    50.95697, 50.98339, 51.00956, 51.0355, 51.0612, 51.08665, 51.11187, 
    51.13684, 51.16156, 51.18605, 51.21029, 51.23429, 51.25804, 51.28155, 
    51.30481, 51.32783, 51.3506, 51.37312, 51.39539, 51.41742, 51.4392, 
    51.46073, 51.48201, 51.50304, 51.52383, 51.54436, 51.56464, 51.58467, 
    51.60445, 51.62397, 51.64325, 51.66227, 51.68103, 51.69955, 51.71781, 
    51.73581, 51.75357, 51.77106, 51.7883, 51.80529, 51.82202, 51.83849, 
    51.85471, 51.87066, 51.88636, 51.90181, 51.91699, 51.93192, 51.94659, 
    51.961, 51.97515, 51.98904, 52.00267, 52.01604, 52.02915, 52.042, 
    52.05458, 52.06691, 52.07898, 52.09078, 52.10232, 52.1136, 52.12461, 
    52.13537, 52.14586, 52.15609, 52.16605, 52.17575, 52.18519, 52.19436, 
    52.20327, 52.21191, 52.22029, 52.2284, 52.23625, 52.24384, 52.25115, 
    52.25821, 52.26499, 52.27151, 52.27777, 52.28376, 52.28948, 52.29494, 
    52.30013, 52.30505, 52.30971, 52.3141, 52.31822, 52.32208, 52.32567, 
    52.32899, 52.33205, 52.33483, 52.33735, 52.33961, 52.34159, 52.34331, 
    52.34476, 52.34594, 52.34686, 52.34751, 52.34789, 52.348, 52.34784, 
    52.34742, 52.34673, 52.34577, 52.34455, 52.34306, 52.34129, 52.33927, 
    52.33697, 52.33441, 52.33158, 52.32848, 52.32512, 52.32149, 52.31759, 
    52.31342, 52.30899, 52.30429, 52.29932, 52.29409, 52.28859, 52.28283, 
    52.2768, 52.2705, 52.26394, 52.25711, 52.25001, 52.24265, 52.23503, 
    52.22713, 52.21898, 52.21056, 52.20187, 52.19292, 52.18371, 52.17423, 
    52.16449, 52.15449, 52.14422, 52.13369, 52.12289, 52.11183, 52.10051, 
    52.08893, 52.07708, 52.06498, 52.05261, 52.03998, 52.02709, 52.01394, 
    52.00053, 51.98686, 51.97293, 51.95874, 51.94429, 51.92958, 51.91461, 
    51.89938, 51.8839, 51.86816, 51.85216, 51.8359, 51.81939, 51.80262, 
    51.78559, 51.76831, 51.75077, 51.73298, 51.71494, 51.69664, 51.67808, 
    51.65928, 51.64021, 51.6209, 51.60133, 51.58152, 51.56145, 51.54113, 
    51.52055, 51.49973, 51.47866, 51.45734, 51.43577, 51.41396, 51.39189, 
    51.36957, 51.34701, 51.3242, 51.30115, 51.27785, 51.2543, 51.23051, 
    51.20647, 51.18219, 51.15767, 51.1329, 51.10789, 51.08264, 51.05715, 
    51.03141, 51.00544, 50.97923, 50.95277, 50.92607, 50.89914, 50.87197, 
    50.84456, 50.81691, 50.78903, 50.76091, 50.73256, 50.70396, 50.67514, 
    50.64608, 50.61679, 50.58727, 50.55751, 50.52752, 50.4973, 50.46684, 
    50.43616, 50.40525, 50.37411, 50.34274, 50.31114, 50.27932, 50.24726, 
    50.21498, 50.18248, 50.14975, 50.1168, 50.08362, 50.05022, 50.01659, 
    49.98275, 49.94868, 49.91439, 49.87988, 49.84515, 49.8102, 49.77503, 
    49.73964, 49.70404, 49.66822, 49.63218, 49.59592, 49.55946, 49.52277, 
    49.48587, 49.44876, 49.41144, 49.3739, 49.33615, 49.29819, 49.26003, 
    49.22165, 49.18306, 49.14426, 49.10526, 49.06604, 49.02663, 48.987, 
    48.94717, 48.90714, 48.86689, 48.82645, 48.7858, 48.74496, 48.70391, 
    48.66265, 48.6212,
  44.07914, 44.13659, 44.19389, 44.25105, 44.30807, 44.36493, 44.42166, 
    44.47823, 44.53466, 44.59095, 44.64708, 44.70306, 44.7589, 44.81458, 
    44.87012, 44.9255, 44.98073, 45.03581, 45.09074, 45.14551, 45.20013, 
    45.25459, 45.3089, 45.36306, 45.41705, 45.47089, 45.52457, 45.57809, 
    45.63146, 45.68466, 45.73771, 45.79059, 45.84331, 45.89587, 45.94827, 
    46.0005, 46.05257, 46.10448, 46.15622, 46.2078, 46.25921, 46.31045, 
    46.36153, 46.41243, 46.46317, 46.51374, 46.56414, 46.61437, 46.66442, 
    46.71431, 46.76402, 46.81356, 46.86293, 46.91212, 46.96114, 47.00998, 
    47.05864, 47.10713, 47.15544, 47.20358, 47.25153, 47.2993, 47.3469, 
    47.39431, 47.44154, 47.48859, 47.53546, 47.58215, 47.62865, 47.67496, 
    47.7211, 47.76704, 47.81281, 47.85838, 47.90376, 47.94896, 47.99397, 
    48.03879, 48.08342, 48.12786, 48.1721, 48.21616, 48.26002, 48.30369, 
    48.34716, 48.39045, 48.43353, 48.47642, 48.51912, 48.56161, 48.60391, 
    48.64601, 48.68791, 48.72961, 48.77111, 48.81242, 48.85352, 48.89441, 
    48.93511, 48.9756, 49.01589, 49.05597, 49.09585, 49.13552, 49.17499, 
    49.21424, 49.2533, 49.29214, 49.33077, 49.36919, 49.40741, 49.44541, 
    49.4832, 49.52079, 49.55815, 49.59531, 49.63225, 49.66897, 49.70548, 
    49.74178, 49.77786, 49.81372, 49.84937, 49.88479, 49.92, 49.95499, 
    49.98976, 50.0243, 50.05863, 50.09274, 50.12662, 50.16028, 50.19372, 
    50.22694, 50.25993, 50.29269, 50.32523, 50.35754, 50.38963, 50.42148, 
    50.45311, 50.48451, 50.51569, 50.54663, 50.57734, 50.60782, 50.63807, 
    50.66809, 50.69788, 50.72743, 50.75675, 50.78584, 50.81469, 50.84331, 
    50.87169, 50.89983, 50.92774, 50.95541, 50.98284, 51.01004, 51.03699, 
    51.06371, 51.09019, 51.11642, 51.14242, 51.16817, 51.19369, 51.21896, 
    51.24398, 51.26877, 51.29331, 51.31761, 51.34166, 51.36547, 51.38903, 
    51.41234, 51.43541, 51.45823, 51.48081, 51.50313, 51.52521, 51.54704, 
    51.56862, 51.58995, 51.61103, 51.63186, 51.65244, 51.67277, 51.69284, 
    51.71267, 51.73224, 51.75156, 51.77063, 51.78944, 51.80799, 51.8263, 
    51.84435, 51.86214, 51.87968, 51.89696, 51.91398, 51.93075, 51.94727, 
    51.96352, 51.97952, 51.99525, 52.01073, 52.02596, 52.04092, 52.05562, 
    52.07006, 52.08425, 52.09817, 52.11184, 52.12524, 52.13838, 52.15126, 
    52.16388, 52.17623, 52.18832, 52.20016, 52.21173, 52.22303, 52.23407, 
    52.24485, 52.25537, 52.26562, 52.27561, 52.28533, 52.29479, 52.30399, 
    52.31292, 52.32158, 52.32998, 52.33811, 52.34598, 52.35358, 52.36092, 
    52.36799, 52.37479, 52.38133, 52.3876, 52.3936, 52.39934, 52.40481, 
    52.41001, 52.41495, 52.41962, 52.42402, 52.42815, 52.43201, 52.43561, 
    52.43894, 52.44201, 52.4448, 52.44733, 52.44958, 52.45158, 52.4533, 
    52.45475, 52.45594, 52.45686, 52.4575, 52.45789, 52.458, 52.45784, 
    52.45742, 52.45673, 52.45577, 52.45454, 52.45304, 52.45128, 52.44925, 
    52.44695, 52.44438, 52.44154, 52.43843, 52.43506, 52.43142, 52.42751, 
    52.42334, 52.4189, 52.41418, 52.40921, 52.40396, 52.39845, 52.39267, 
    52.38662, 52.38031, 52.37373, 52.36689, 52.35978, 52.3524, 52.34475, 
    52.33684, 52.32867, 52.32022, 52.31152, 52.30255, 52.29331, 52.28381, 
    52.27405, 52.26402, 52.25372, 52.24316, 52.23235, 52.22126, 52.20991, 
    52.1983, 52.18643, 52.17429, 52.1619, 52.14924, 52.13631, 52.12313, 
    52.10969, 52.09599, 52.08202, 52.06779, 52.05331, 52.03857, 52.02356, 
    52.0083, 51.99278, 51.977, 51.96096, 51.94467, 51.92812, 51.91131, 
    51.89424, 51.87692, 51.85934, 51.84151, 51.82342, 51.80508, 51.78648, 
    51.76763, 51.74852, 51.72916, 51.70955, 51.68969, 51.66957, 51.6492, 
    51.62859, 51.60772, 51.58659, 51.56522, 51.54361, 51.52174, 51.49962, 
    51.47725, 51.45464, 51.43178, 51.40867, 51.38531, 51.36172, 51.33787, 
    51.31378, 51.28944, 51.26487, 51.24004, 51.21498, 51.18967, 51.16412, 
    51.13832, 51.11229, 51.08601, 51.0595, 51.03275, 51.00575, 50.97852, 
    50.95105, 50.92334, 50.89539, 50.86721, 50.83879, 50.81014, 50.78125, 
    50.75213, 50.72277, 50.69318, 50.66336, 50.6333, 50.60302, 50.5725, 
    50.54175, 50.51077, 50.47956, 50.44812, 50.41646, 50.38456, 50.35244, 
    50.3201, 50.28752, 50.25472, 50.22169, 50.18845, 50.15497, 50.12128, 
    50.08736, 50.05322, 50.01886, 49.98427, 49.94947, 49.91444, 49.8792, 
    49.84374, 49.80806, 49.77216, 49.73605, 49.69972, 49.66318, 49.62642, 
    49.58944, 49.55225, 49.51485, 49.47724, 49.43941, 49.40138, 49.36313, 
    49.32467, 49.28601, 49.24713, 49.20805, 49.16876, 49.12926, 49.08955, 
    49.04964, 49.00953, 48.96921, 48.92868, 48.88796, 48.84703, 48.8059, 
    48.76456, 48.72303,
  44.17286, 44.2304, 44.28779, 44.34504, 44.40214, 44.4591, 44.51591, 
    44.57257, 44.62909, 44.68546, 44.74168, 44.79775, 44.85368, 44.90945, 
    44.96507, 45.02055, 45.07586, 45.13103, 45.18605, 45.24091, 45.29562, 
    45.35017, 45.40456, 45.45881, 45.51289, 45.56682, 45.62059, 45.6742, 
    45.72765, 45.78094, 45.83408, 45.88705, 45.93986, 45.99251, 46.04499, 
    46.09732, 46.14948, 46.20147, 46.2533, 46.30497, 46.35646, 46.40779, 
    46.45896, 46.50995, 46.56078, 46.61143, 46.66192, 46.71224, 46.76238, 
    46.81236, 46.86216, 46.91179, 46.96124, 47.01052, 47.05962, 47.10855, 
    47.1573, 47.20588, 47.25428, 47.30249, 47.35054, 47.3984, 47.44608, 
    47.49358, 47.5409, 47.58804, 47.63499, 47.68176, 47.72835, 47.77475, 
    47.82097, 47.867, 47.91285, 47.95851, 48.00398, 48.04926, 48.09435, 
    48.13926, 48.18397, 48.22849, 48.27283, 48.31696, 48.36091, 48.40466, 
    48.44822, 48.49159, 48.53476, 48.57773, 48.62051, 48.66309, 48.70547, 
    48.74765, 48.78963, 48.83142, 48.873, 48.91438, 48.95557, 48.99654, 
    49.03732, 49.07789, 49.11826, 49.15842, 49.19838, 49.23814, 49.27768, 
    49.31702, 49.35615, 49.39507, 49.43378, 49.47229, 49.51058, 49.54866, 
    49.58653, 49.62418, 49.66163, 49.69886, 49.73588, 49.77268, 49.80927, 
    49.84564, 49.88179, 49.91773, 49.95345, 49.98895, 50.02423, 50.05929, 
    50.09414, 50.12876, 50.16316, 50.19734, 50.23129, 50.26503, 50.29853, 
    50.33182, 50.36488, 50.39771, 50.43032, 50.4627, 50.49486, 50.52679, 
    50.55849, 50.58995, 50.6212, 50.65221, 50.68299, 50.71354, 50.74385, 
    50.77394, 50.80379, 50.83341, 50.86279, 50.89194, 50.92086, 50.94954, 
    50.97798, 51.00619, 51.03416, 51.06189, 51.08939, 51.11664, 51.14366, 
    51.17044, 51.19697, 51.22327, 51.24932, 51.27514, 51.3007, 51.32603, 
    51.35112, 51.37596, 51.40055, 51.42491, 51.44902, 51.47288, 51.49649, 
    51.51986, 51.54298, 51.56586, 51.58849, 51.61086, 51.63299, 51.65487, 
    51.6765, 51.69788, 51.71901, 51.73989, 51.76052, 51.78089, 51.80102, 
    51.82088, 51.8405, 51.85987, 51.87898, 51.89783, 51.91644, 51.93478, 
    51.95287, 51.97071, 51.98829, 52.00561, 52.02267, 52.03948, 52.05603, 
    52.07233, 52.08836, 52.10414, 52.11965, 52.13491, 52.14991, 52.16465, 
    52.17913, 52.19334, 52.2073, 52.221, 52.23443, 52.2476, 52.26051, 
    52.27316, 52.28555, 52.29767, 52.30953, 52.32113, 52.33246, 52.34353, 
    52.35434, 52.36488, 52.37515, 52.38517, 52.39491, 52.40439, 52.41361, 
    52.42256, 52.43125, 52.43967, 52.44782, 52.45571, 52.46333, 52.47068, 
    52.47777, 52.48459, 52.49114, 52.49743, 52.50344, 52.50919, 52.51468, 
    52.51989, 52.52484, 52.52952, 52.53393, 52.53808, 52.54195, 52.54556, 
    52.5489, 52.55197, 52.55477, 52.5573, 52.55957, 52.56156, 52.56329, 
    52.56474, 52.56593, 52.56685, 52.5675, 52.56789, 52.568, 52.56784, 
    52.56742, 52.56673, 52.56576, 52.56453, 52.56303, 52.56126, 52.55922, 
    52.55692, 52.55434, 52.5515, 52.54839, 52.54501, 52.54136, 52.53744, 
    52.53325, 52.5288, 52.52408, 52.51909, 52.51383, 52.5083, 52.50251, 
    52.49645, 52.49012, 52.48352, 52.47667, 52.46954, 52.46214, 52.45448, 
    52.44655, 52.43835, 52.42989, 52.42116, 52.41217, 52.40291, 52.39339, 
    52.3836, 52.37355, 52.36323, 52.35264, 52.3418, 52.33068, 52.31931, 
    52.30767, 52.29577, 52.2836, 52.27118, 52.25849, 52.24554, 52.23232, 
    52.21885, 52.20511, 52.19111, 52.17685, 52.16233, 52.14755, 52.13251, 
    52.11721, 52.10166, 52.08584, 52.06977, 52.05343, 52.03684, 52.01999, 
    52.00288, 51.98552, 51.9679, 51.95003, 51.9319, 51.91351, 51.89487, 
    51.87597, 51.85682, 51.83742, 51.81776, 51.79785, 51.77769, 51.75727, 
    51.7366, 51.71569, 51.69452, 51.6731, 51.65143, 51.62951, 51.60734, 
    51.58492, 51.56226, 51.53934, 51.51618, 51.49277, 51.46912, 51.44522, 
    51.42107, 51.39668, 51.37205, 51.34717, 51.32204, 51.29668, 51.27107, 
    51.24522, 51.21912, 51.19279, 51.16621, 51.1394, 51.11235, 51.08505, 
    51.05752, 51.02975, 51.00174, 50.9735, 50.94502, 50.9163, 50.88735, 
    50.85816, 50.82874, 50.79908, 50.7692, 50.73907, 50.70872, 50.67813, 
    50.64732, 50.61627, 50.58499, 50.55349, 50.52175, 50.48979, 50.4576, 
    50.42518, 50.39254, 50.35966, 50.32657, 50.29325, 50.2597, 50.22594, 
    50.19194, 50.15773, 50.12329, 50.08864, 50.05376, 50.01867, 49.98335, 
    49.94781, 49.91206, 49.87609, 49.8399, 49.80349, 49.76687, 49.73003, 
    49.69299, 49.65572, 49.61824, 49.58055, 49.54265, 49.50453, 49.46621, 
    49.42767, 49.38893, 49.34997, 49.31081, 49.27144, 49.23186, 49.19207, 
    49.15208, 49.11189, 49.07149, 49.03088, 48.99007, 48.94907, 48.90785, 
    48.86644, 48.82482,
  44.26653, 44.32415, 44.38163, 44.43896, 44.49615, 44.5532, 44.6101, 
    44.66685, 44.72346, 44.77991, 44.83623, 44.89239, 44.9484, 45.00426, 
    45.05997, 45.11554, 45.17094, 45.2262, 45.2813, 45.33625, 45.39105, 
    45.44569, 45.50018, 45.5545, 45.60868, 45.6627, 45.71655, 45.77026, 
    45.8238, 45.87718, 45.9304, 45.98346, 46.03636, 46.0891, 46.14167, 
    46.19408, 46.24633, 46.29841, 46.35033, 46.40208, 46.45367, 46.50509, 
    46.55634, 46.60743, 46.65834, 46.70908, 46.75966, 46.81006, 46.8603, 
    46.91036, 46.96025, 47.00996, 47.0595, 47.10887, 47.15806, 47.20708, 
    47.25592, 47.30458, 47.35307, 47.40137, 47.4495, 47.49745, 47.54522, 
    47.5928, 47.64021, 47.68744, 47.73447, 47.78133, 47.82801, 47.8745, 
    47.9208, 47.96692, 48.01285, 48.05859, 48.10415, 48.14952, 48.1947, 
    48.23969, 48.28448, 48.32909, 48.37351, 48.41773, 48.46177, 48.5056, 
    48.54924, 48.59269, 48.63594, 48.679, 48.72186, 48.76453, 48.80699, 
    48.84925, 48.89132, 48.93319, 48.97485, 49.01632, 49.05758, 49.09864, 
    49.1395, 49.18015, 49.2206, 49.26085, 49.30088, 49.34072, 49.38034, 
    49.41976, 49.45897, 49.49797, 49.53676, 49.57534, 49.61371, 49.65187, 
    49.68982, 49.72755, 49.76508, 49.80238, 49.83948, 49.87636, 49.91302, 
    49.94947, 49.9857, 50.02171, 50.05751, 50.09308, 50.12844, 50.16357, 
    50.19849, 50.23318, 50.26766, 50.30191, 50.33594, 50.36974, 50.40332, 
    50.43668, 50.46981, 50.50272, 50.5354, 50.56785, 50.60007, 50.63207, 
    50.66384, 50.69538, 50.72668, 50.75776, 50.78861, 50.81923, 50.84961, 
    50.87976, 50.90968, 50.93937, 50.96881, 50.99803, 51.02701, 51.05575, 
    51.08426, 51.11253, 51.14056, 51.16836, 51.19592, 51.22323, 51.25031, 
    51.27715, 51.30374, 51.3301, 51.35621, 51.38208, 51.40771, 51.4331, 
    51.45824, 51.48314, 51.50779, 51.5322, 51.55636, 51.58028, 51.60395, 
    51.62737, 51.65054, 51.67347, 51.69615, 51.71858, 51.74076, 51.76269, 
    51.78437, 51.8058, 51.82698, 51.84791, 51.86858, 51.88901, 51.90918, 
    51.92909, 51.94876, 51.96817, 51.98732, 52.00622, 52.02487, 52.04326, 
    52.06139, 52.07927, 52.09689, 52.11425, 52.13136, 52.1482, 52.16479, 
    52.18113, 52.1972, 52.21301, 52.22857, 52.24386, 52.2589, 52.27367, 
    52.28818, 52.30243, 52.31643, 52.33015, 52.34362, 52.35682, 52.36977, 
    52.38245, 52.39486, 52.40701, 52.4189, 52.43053, 52.44189, 52.45298, 
    52.46381, 52.47438, 52.48468, 52.49472, 52.50449, 52.51399, 52.52323, 
    52.53221, 52.54091, 52.54935, 52.55753, 52.56543, 52.57307, 52.58044, 
    52.58755, 52.59438, 52.60095, 52.60725, 52.61329, 52.61905, 52.62455, 
    52.62978, 52.63474, 52.63943, 52.64385, 52.648, 52.65189, 52.6555, 
    52.65885, 52.66193, 52.66473, 52.66727, 52.66954, 52.67154, 52.67327, 
    52.67474, 52.67593, 52.67685, 52.6775, 52.67789, 52.678, 52.67784, 
    52.67742, 52.67672, 52.67576, 52.67452, 52.67302, 52.67125, 52.6692, 
    52.66689, 52.66431, 52.66146, 52.65834, 52.65495, 52.65129, 52.64737, 
    52.64317, 52.6387, 52.63397, 52.62897, 52.6237, 52.61816, 52.61235, 
    52.60627, 52.59993, 52.59332, 52.58644, 52.57929, 52.57188, 52.5642, 
    52.55625, 52.54803, 52.53955, 52.5308, 52.52179, 52.51251, 52.50296, 
    52.49315, 52.48307, 52.47273, 52.46212, 52.45124, 52.44011, 52.4287, 
    52.41704, 52.40511, 52.39291, 52.38046, 52.36774, 52.35475, 52.34151, 
    52.328, 52.31423, 52.3002, 52.2859, 52.27135, 52.25653, 52.24146, 
    52.22612, 52.21053, 52.19468, 52.17856, 52.16219, 52.14556, 52.12867, 
    52.11152, 52.09412, 52.07646, 52.05854, 52.04036, 52.02193, 52.00325, 
    51.98431, 51.96511, 51.94566, 51.92596, 51.906, 51.88579, 51.86533, 
    51.84462, 51.82365, 51.80243, 51.78096, 51.75924, 51.73727, 51.71505, 
    51.69258, 51.66986, 51.6469, 51.62368, 51.60022, 51.57651, 51.55256, 
    51.52835, 51.50391, 51.47921, 51.45428, 51.4291, 51.40368, 51.37801, 
    51.3521, 51.32594, 51.29955, 51.27291, 51.24604, 51.21893, 51.19157, 
    51.16398, 51.13614, 51.10807, 51.07977, 51.05122, 51.02244, 50.99342, 
    50.96417, 50.93468, 50.90496, 50.87501, 50.84482, 50.8144, 50.78375, 
    50.75286, 50.72175, 50.6904, 50.65883, 50.62703, 50.59499, 50.56273, 
    50.53024, 50.49753, 50.46459, 50.43142, 50.39803, 50.36441, 50.33057, 
    50.29651, 50.26222, 50.22771, 50.19298, 50.15803, 50.12286, 50.08747, 
    50.05186, 50.01603, 49.97998, 49.94372, 49.90723, 49.87054, 49.83363, 
    49.7965, 49.75916, 49.7216, 49.68383, 49.64585, 49.60766, 49.56925, 
    49.53064, 49.49181, 49.45278, 49.41354, 49.37409, 49.33443, 49.29456, 
    49.25449, 49.21422, 49.17374, 49.13305, 49.09216, 49.05107, 49.00977, 
    48.96828, 48.92658,
  44.36013, 44.41785, 44.47541, 44.53284, 44.59011, 44.64725, 44.70424, 
    44.76108, 44.81777, 44.87432, 44.93072, 44.98697, 45.04307, 45.09902, 
    45.15482, 45.21047, 45.26597, 45.32131, 45.37651, 45.43155, 45.48643, 
    45.54116, 45.59573, 45.65015, 45.70441, 45.75852, 45.81247, 45.86626, 
    45.91989, 45.97336, 46.02667, 46.07982, 46.13281, 46.18563, 46.2383, 
    46.2908, 46.34314, 46.39531, 46.44731, 46.49915, 46.55083, 46.60234, 
    46.65368, 46.70485, 46.75585, 46.80669, 46.85735, 46.90784, 46.95816, 
    47.00831, 47.05829, 47.10809, 47.15772, 47.20718, 47.25646, 47.30556, 
    47.35449, 47.40324, 47.45181, 47.50021, 47.54842, 47.59646, 47.64431, 
    47.69199, 47.73948, 47.78679, 47.83392, 47.88086, 47.92762, 47.9742, 
    48.02059, 48.0668, 48.11281, 48.15864, 48.20428, 48.24974, 48.295, 
    48.34008, 48.38496, 48.42965, 48.47416, 48.51846, 48.56258, 48.6065, 
    48.65023, 48.69376, 48.7371, 48.78024, 48.82318, 48.86593, 48.90848, 
    48.95082, 48.99297, 49.03492, 49.07667, 49.11822, 49.15956, 49.20071, 
    49.24165, 49.28238, 49.32291, 49.36324, 49.40335, 49.44327, 49.48297, 
    49.52247, 49.56176, 49.60084, 49.63971, 49.67837, 49.71682, 49.75506, 
    49.79308, 49.8309, 49.8685, 49.90588, 49.94305, 49.98001, 50.01675, 
    50.05327, 50.08958, 50.12566, 50.16153, 50.19719, 50.23262, 50.26783, 
    50.30282, 50.33759, 50.37214, 50.40646, 50.44056, 50.47444, 50.50809, 
    50.54152, 50.57472, 50.6077, 50.64045, 50.67297, 50.70527, 50.73733, 
    50.76917, 50.80078, 50.83215, 50.8633, 50.89421, 50.9249, 50.95535, 
    50.98557, 51.01555, 51.0453, 51.07482, 51.1041, 51.13314, 51.16195, 
    51.19052, 51.21885, 51.24695, 51.27481, 51.30243, 51.3298, 51.35694, 
    51.38384, 51.4105, 51.43691, 51.46309, 51.48901, 51.5147, 51.54015, 
    51.56535, 51.5903, 51.61501, 51.63947, 51.66369, 51.68766, 51.71139, 
    51.73486, 51.75809, 51.78107, 51.80381, 51.82629, 51.84852, 51.8705, 
    51.89223, 51.91371, 51.93494, 51.95592, 51.97664, 51.99711, 52.01733, 
    52.03729, 52.057, 52.07646, 52.09566, 52.1146, 52.13329, 52.15173, 
    52.1699, 52.18782, 52.20548, 52.22289, 52.24004, 52.25692, 52.27355, 
    52.28992, 52.30603, 52.32188, 52.33748, 52.35281, 52.36788, 52.38269, 
    52.39724, 52.41152, 52.42554, 52.43931, 52.4528, 52.46604, 52.47902, 
    52.49172, 52.50417, 52.51635, 52.52827, 52.53992, 52.55131, 52.56243, 
    52.57329, 52.58388, 52.59421, 52.60427, 52.61406, 52.62359, 52.63285, 
    52.64185, 52.65058, 52.65904, 52.66723, 52.67516, 52.68281, 52.6902, 
    52.69732, 52.70418, 52.71076, 52.71708, 52.72313, 52.7289, 52.73442, 
    52.73966, 52.74463, 52.74933, 52.75377, 52.75793, 52.76182, 52.76545, 
    52.7688, 52.77189, 52.7747, 52.77725, 52.77952, 52.78153, 52.78326, 
    52.78473, 52.78592, 52.78685, 52.7875, 52.78788, 52.788, 52.78784, 
    52.78741, 52.78672, 52.78575, 52.78452, 52.78301, 52.78123, 52.77918, 
    52.77686, 52.77428, 52.77142, 52.76829, 52.76489, 52.76123, 52.75729, 
    52.75308, 52.74861, 52.74386, 52.73885, 52.73356, 52.72801, 52.72219, 
    52.7161, 52.70974, 52.70311, 52.69622, 52.68905, 52.68162, 52.67392, 
    52.66595, 52.65771, 52.64921, 52.64044, 52.63141, 52.6221, 52.61253, 
    52.6027, 52.59259, 52.58223, 52.57159, 52.56069, 52.54953, 52.5381, 
    52.5264, 52.51444, 52.50222, 52.48973, 52.47698, 52.46397, 52.45069, 
    52.43715, 52.42334, 52.40928, 52.39495, 52.38036, 52.36551, 52.3504, 
    52.33503, 52.3194, 52.3035, 52.28735, 52.27094, 52.25427, 52.23734, 
    52.22015, 52.20271, 52.18501, 52.16704, 52.14883, 52.13035, 52.11162, 
    52.09264, 52.0734, 52.0539, 52.03415, 52.01415, 51.99389, 51.97338, 
    51.95261, 51.9316, 51.91033, 51.88881, 51.86704, 51.84502, 51.82275, 
    51.80022, 51.77745, 51.75444, 51.73117, 51.70765, 51.68389, 51.65988, 
    51.63562, 51.61112, 51.58637, 51.56137, 51.53614, 51.51065, 51.48493, 
    51.45896, 51.43275, 51.4063, 51.3796, 51.35266, 51.32549, 51.29807, 
    51.27042, 51.24252, 51.21439, 51.18602, 51.15741, 51.12856, 51.09948, 
    51.07016, 51.04061, 51.01083, 50.9808, 50.95055, 50.92006, 50.88934, 
    50.85839, 50.82721, 50.79579, 50.76415, 50.73228, 50.70017, 50.66784, 
    50.63528, 50.6025, 50.56948, 50.53625, 50.50278, 50.46909, 50.43518, 
    50.40105, 50.36668, 50.3321, 50.2973, 50.26227, 50.22703, 50.19156, 
    50.15588, 50.11997, 50.08385, 50.04751, 50.01095, 49.97418, 49.93719, 
    49.89998, 49.86256, 49.82493, 49.78708, 49.74902, 49.71075, 49.67227, 
    49.63358, 49.59467, 49.55556, 49.51624, 49.4767, 49.43697, 49.39702, 
    49.35687, 49.31651, 49.27595, 49.23518, 49.19421, 49.15304, 49.11166, 
    49.07008, 49.0283,
  44.45369, 44.51148, 44.56914, 44.62665, 44.68402, 44.74124, 44.79832, 
    44.85525, 44.91203, 44.96867, 45.02515, 45.08149, 45.13768, 45.19373, 
    45.24961, 45.30535, 45.36094, 45.41637, 45.47165, 45.52678, 45.58176, 
    45.63657, 45.69124, 45.74575, 45.8001, 45.85429, 45.90833, 45.96221, 
    46.01593, 46.06949, 46.12289, 46.17612, 46.2292, 46.28212, 46.33487, 
    46.38746, 46.43989, 46.49215, 46.54424, 46.59617, 46.64794, 46.69954, 
    46.75097, 46.80222, 46.85332, 46.90424, 46.95499, 47.00557, 47.05598, 
    47.10622, 47.15628, 47.20618, 47.25589, 47.30544, 47.3548, 47.404, 
    47.45301, 47.50185, 47.55051, 47.599, 47.6473, 47.69542, 47.74337, 
    47.79113, 47.83871, 47.8861, 47.93332, 47.98035, 48.0272, 48.07386, 
    48.12034, 48.16663, 48.21273, 48.25865, 48.30438, 48.34992, 48.39527, 
    48.44043, 48.4854, 48.53018, 48.57476, 48.61916, 48.66336, 48.70736, 
    48.75117, 48.79479, 48.83821, 48.88144, 48.92447, 48.9673, 49.00993, 
    49.05236, 49.09459, 49.13662, 49.17846, 49.22009, 49.26151, 49.30273, 
    49.34376, 49.38457, 49.42519, 49.46559, 49.50579, 49.54578, 49.58557, 
    49.62515, 49.66452, 49.70368, 49.74263, 49.78137, 49.8199, 49.85821, 
    49.89632, 49.93421, 49.97189, 50.00935, 50.0466, 50.08363, 50.12045, 
    50.15705, 50.19343, 50.22959, 50.26554, 50.30127, 50.33677, 50.37206, 
    50.40712, 50.44197, 50.47659, 50.51099, 50.54516, 50.57911, 50.61283, 
    50.64634, 50.67961, 50.71266, 50.74548, 50.77807, 50.81044, 50.84257, 
    50.87448, 50.90615, 50.9376, 50.96882, 50.9998, 51.03055, 51.06107, 
    51.09135, 51.1214, 51.15122, 51.1808, 51.21015, 51.23926, 51.26813, 
    51.29676, 51.32516, 51.35332, 51.38124, 51.40892, 51.43636, 51.46356, 
    51.49052, 51.51723, 51.54371, 51.56994, 51.59593, 51.62168, 51.64718, 
    51.67244, 51.69745, 51.72222, 51.74674, 51.77101, 51.79504, 51.81882, 
    51.84235, 51.86563, 51.88866, 51.91145, 51.93398, 51.95626, 51.9783, 
    52.00008, 52.02161, 52.04289, 52.06392, 52.08469, 52.10521, 52.12547, 
    52.14548, 52.16524, 52.18474, 52.20399, 52.22298, 52.24171, 52.26019, 
    52.2784, 52.29637, 52.31407, 52.33152, 52.34871, 52.36563, 52.38231, 
    52.39871, 52.41486, 52.43075, 52.44638, 52.46175, 52.47686, 52.4917, 
    52.50628, 52.5206, 52.53466, 52.54845, 52.56199, 52.57526, 52.58826, 
    52.601, 52.61348, 52.62569, 52.63763, 52.64931, 52.66073, 52.67188, 
    52.68277, 52.69338, 52.70374, 52.71382, 52.72364, 52.73319, 52.74247, 
    52.75149, 52.76024, 52.76872, 52.77693, 52.78488, 52.79255, 52.79996, 
    52.8071, 52.81397, 52.82057, 52.8269, 52.83297, 52.83876, 52.84428, 
    52.84954, 52.85452, 52.85924, 52.86368, 52.86786, 52.87176, 52.87539, 
    52.87876, 52.88185, 52.88467, 52.88722, 52.8895, 52.89151, 52.89325, 
    52.89472, 52.89592, 52.89684, 52.8975, 52.89788, 52.898, 52.89784, 
    52.89742, 52.89672, 52.89575, 52.8945, 52.89299, 52.89121, 52.88916, 
    52.88684, 52.88424, 52.88138, 52.87824, 52.87484, 52.87116, 52.86721, 
    52.863, 52.85851, 52.85375, 52.84872, 52.84343, 52.83786, 52.83203, 
    52.82592, 52.81955, 52.8129, 52.80599, 52.79881, 52.79136, 52.78364, 
    52.77565, 52.7674, 52.75887, 52.75008, 52.74102, 52.7317, 52.7221, 
    52.71224, 52.70211, 52.69172, 52.68106, 52.67014, 52.65894, 52.64748, 
    52.63576, 52.62377, 52.61152, 52.599, 52.58622, 52.57317, 52.55986, 
    52.54629, 52.53246, 52.51836, 52.50399, 52.48937, 52.47448, 52.45934, 
    52.44393, 52.42826, 52.41233, 52.39613, 52.37968, 52.36297, 52.346, 
    52.32878, 52.31129, 52.29354, 52.27554, 52.25728, 52.23876, 52.21999, 
    52.20096, 52.18167, 52.16213, 52.14233, 52.12228, 52.10198, 52.08142, 
    52.0606, 52.03954, 52.01822, 51.99665, 51.97483, 51.95276, 51.93044, 
    51.90786, 51.88504, 51.86197, 51.83864, 51.81507, 51.79125, 51.76719, 
    51.74287, 51.71832, 51.69351, 51.66846, 51.64316, 51.61762, 51.59184, 
    51.56581, 51.53954, 51.51303, 51.48627, 51.45927, 51.43203, 51.40456, 
    51.37684, 51.34888, 51.32069, 51.29225, 51.26358, 51.23467, 51.20552, 
    51.17614, 51.14652, 51.11666, 51.08658, 51.05626, 51.0257, 50.99492, 
    50.96389, 50.93264, 50.90116, 50.86945, 50.83751, 50.80533, 50.77293, 
    50.7403, 50.70745, 50.67436, 50.64105, 50.60752, 50.57375, 50.53977, 
    50.50556, 50.47113, 50.43647, 50.40159, 50.36649, 50.33117, 50.29563, 
    50.25987, 50.22389, 50.18769, 50.15127, 50.11464, 50.07779, 50.04072, 
    50.00344, 49.96594, 49.92823, 49.8903, 49.85217, 49.81382, 49.77525, 
    49.73648, 49.6975, 49.65831, 49.6189, 49.57929, 49.53947, 49.49945, 
    49.45921, 49.41877, 49.37813, 49.33728, 49.29623, 49.25497, 49.21351, 
    49.17185, 49.12999,
  44.54718, 44.60506, 44.66281, 44.72041, 44.77787, 44.83518, 44.89234, 
    44.94936, 45.00623, 45.06296, 45.11954, 45.17596, 45.23224, 45.28837, 
    45.34435, 45.40018, 45.45585, 45.51138, 45.56675, 45.62197, 45.67703, 
    45.73194, 45.78669, 45.84129, 45.89573, 45.95001, 46.00414, 46.05811, 
    46.11192, 46.16557, 46.21906, 46.27238, 46.32555, 46.37856, 46.4314, 
    46.48407, 46.53659, 46.58894, 46.64112, 46.69315, 46.745, 46.79668, 
    46.8482, 46.89955, 46.95073, 47.00174, 47.05259, 47.10326, 47.15376, 
    47.20408, 47.25423, 47.30421, 47.35402, 47.40365, 47.45311, 47.50239, 
    47.55149, 47.60042, 47.64917, 47.69774, 47.74613, 47.79434, 47.84237, 
    47.89022, 47.93789, 47.98537, 48.03268, 48.0798, 48.12673, 48.17348, 
    48.22004, 48.26642, 48.31261, 48.35862, 48.40443, 48.45006, 48.49549, 
    48.54074, 48.5858, 48.63066, 48.67533, 48.71981, 48.7641, 48.80819, 
    48.85209, 48.89579, 48.93929, 48.9826, 49.02571, 49.06863, 49.11134, 
    49.15386, 49.19617, 49.23829, 49.2802, 49.32191, 49.36342, 49.40473, 
    49.44584, 49.48673, 49.52743, 49.56791, 49.6082, 49.64827, 49.68814, 
    49.72779, 49.76725, 49.80648, 49.84552, 49.88433, 49.92294, 49.96134, 
    49.99952, 50.03749, 50.07525, 50.11279, 50.15012, 50.18723, 50.22412, 
    50.2608, 50.29725, 50.33349, 50.36951, 50.40532, 50.4409, 50.47626, 
    50.5114, 50.54632, 50.58101, 50.61549, 50.64973, 50.68375, 50.71755, 
    50.75113, 50.78447, 50.81759, 50.85049, 50.88315, 50.91558, 50.94779, 
    50.97977, 51.01151, 51.04303, 51.07431, 51.10537, 51.13618, 51.16677, 
    51.19712, 51.22724, 51.25712, 51.28677, 51.31618, 51.34535, 51.37429, 
    51.40299, 51.43145, 51.45967, 51.48766, 51.5154, 51.5429, 51.57016, 
    51.59718, 51.62396, 51.65049, 51.67679, 51.70284, 51.72864, 51.7542, 
    51.77952, 51.80458, 51.82941, 51.85398, 51.87831, 51.9024, 51.92623, 
    51.94982, 51.97316, 51.99624, 52.01908, 52.04167, 52.064, 52.08609, 
    52.10792, 52.1295, 52.15083, 52.1719, 52.19273, 52.21329, 52.2336, 
    52.25366, 52.27347, 52.29301, 52.31231, 52.33134, 52.35012, 52.36864, 
    52.3869, 52.40491, 52.42265, 52.44014, 52.45737, 52.47434, 52.49105, 
    52.5075, 52.52369, 52.53961, 52.55528, 52.57068, 52.58583, 52.60071, 
    52.61533, 52.62968, 52.64377, 52.6576, 52.67117, 52.68446, 52.6975, 
    52.71027, 52.72278, 52.73502, 52.74699, 52.75871, 52.77015, 52.78133, 
    52.79224, 52.80288, 52.81326, 52.82337, 52.83321, 52.84278, 52.85209, 
    52.86113, 52.8699, 52.8784, 52.88663, 52.8946, 52.90229, 52.90972, 
    52.91688, 52.92376, 52.93038, 52.93673, 52.94281, 52.94862, 52.95415, 
    52.95942, 52.96442, 52.96914, 52.97359, 52.97778, 52.98169, 52.98534, 
    52.98871, 52.99181, 52.99464, 52.9972, 52.99948, 53.0015, 53.00324, 
    53.00471, 53.00591, 53.00684, 53.0075, 53.00788, 53.008, 53.00784, 
    53.00741, 53.00671, 53.00574, 53.0045, 53.00298, 53.00119, 52.99914, 
    52.99681, 52.99421, 52.99134, 52.98819, 52.98478, 52.98109, 52.97714, 
    52.97291, 52.96841, 52.96364, 52.9586, 52.95329, 52.94772, 52.94186, 
    52.93575, 52.92935, 52.92269, 52.91576, 52.90857, 52.9011, 52.89336, 
    52.88535, 52.87708, 52.86853, 52.85972, 52.85064, 52.84129, 52.83167, 
    52.82178, 52.81163, 52.80121, 52.79053, 52.77958, 52.76836, 52.75687, 
    52.74512, 52.7331, 52.72082, 52.70827, 52.69546, 52.68238, 52.66904, 
    52.65543, 52.64156, 52.62743, 52.61303, 52.59837, 52.58345, 52.56826, 
    52.55282, 52.53711, 52.52114, 52.50491, 52.48842, 52.47167, 52.45466, 
    52.43739, 52.41986, 52.40208, 52.38403, 52.36573, 52.34716, 52.32835, 
    52.30927, 52.28994, 52.27035, 52.25051, 52.23041, 52.21006, 52.18945, 
    52.16859, 52.14747, 52.1261, 52.10448, 52.08261, 52.06049, 52.03811, 
    52.01548, 51.99261, 51.96948, 51.94611, 51.92248, 51.89861, 51.87449, 
    51.85012, 51.8255, 51.80064, 51.77553, 51.75018, 51.72458, 51.69873, 
    51.67265, 51.64631, 51.61974, 51.59292, 51.56586, 51.53857, 51.51102, 
    51.48325, 51.45522, 51.42696, 51.39846, 51.36973, 51.34075, 51.31154, 
    51.28209, 51.25241, 51.22249, 51.19233, 51.16195, 51.13132, 51.10047, 
    51.06938, 51.03806, 51.00651, 50.97472, 50.94271, 50.91047, 50.878, 
    50.8453, 50.81237, 50.77921, 50.74583, 50.71222, 50.67839, 50.64433, 
    50.61005, 50.57554, 50.54081, 50.50586, 50.47068, 50.43529, 50.39967, 
    50.36383, 50.32778, 50.2915, 50.25501, 50.2183, 50.18137, 50.14423, 
    50.10686, 50.06929, 50.0315, 49.9935, 49.95528, 49.91685, 49.87821, 
    49.83936, 49.80029, 49.76102, 49.72153, 49.68184, 49.64194, 49.60184, 
    49.56152, 49.521, 49.48028, 49.43935, 49.39821, 49.35687, 49.31533, 
    49.27359, 49.23164,
  44.64061, 44.69859, 44.75642, 44.81411, 44.87166, 44.92906, 44.98631, 
    45.04342, 45.10038, 45.1572, 45.21386, 45.27038, 45.32675, 45.38297, 
    45.43903, 45.49495, 45.55072, 45.60633, 45.66179, 45.71709, 45.77225, 
    45.82725, 45.88209, 45.93678, 45.99131, 46.04568, 46.0999, 46.15395, 
    46.20785, 46.26159, 46.31517, 46.36859, 46.42184, 46.47494, 46.52787, 
    46.58064, 46.63324, 46.68568, 46.73796, 46.79007, 46.84201, 46.89378, 
    46.94539, 46.99683, 47.0481, 47.0992, 47.15013, 47.20089, 47.25148, 
    47.30189, 47.35213, 47.40221, 47.4521, 47.50182, 47.55136, 47.60073, 
    47.64993, 47.69894, 47.74778, 47.79644, 47.84492, 47.89322, 47.94133, 
    47.98927, 48.03703, 48.0846, 48.13199, 48.1792, 48.22622, 48.27306, 
    48.31971, 48.36617, 48.41245, 48.45854, 48.50444, 48.55016, 48.59568, 
    48.64101, 48.68615, 48.7311, 48.77586, 48.82042, 48.8648, 48.90897, 
    48.95295, 48.99674, 49.04033, 49.08372, 49.12692, 49.16992, 49.21272, 
    49.25532, 49.29772, 49.33992, 49.38191, 49.42371, 49.4653, 49.50669, 
    49.54788, 49.58886, 49.62963, 49.6702, 49.71057, 49.75072, 49.79067, 
    49.83041, 49.86994, 49.90926, 49.94837, 49.98727, 50.02596, 50.06443, 
    50.1027, 50.14074, 50.17858, 50.2162, 50.2536, 50.29079, 50.32776, 
    50.36451, 50.40105, 50.43737, 50.47346, 50.50934, 50.545, 50.58044, 
    50.61565, 50.65064, 50.68541, 50.71996, 50.75428, 50.78838, 50.82225, 
    50.8559, 50.88931, 50.9225, 50.95547, 50.9882, 51.02071, 51.05299, 
    51.08503, 51.11685, 51.14843, 51.17979, 51.21091, 51.24179, 51.27245, 
    51.30287, 51.33305, 51.363, 51.39272, 51.42219, 51.45143, 51.48043, 
    51.5092, 51.53772, 51.56601, 51.59405, 51.62186, 51.64943, 51.67675, 
    51.70383, 51.73067, 51.75726, 51.78362, 51.80973, 51.83559, 51.86121, 
    51.88658, 51.91171, 51.93659, 51.96122, 51.98561, 52.00975, 52.03364, 
    52.05728, 52.08067, 52.10381, 52.1267, 52.14934, 52.17173, 52.19386, 
    52.21575, 52.23738, 52.25876, 52.27988, 52.30075, 52.32137, 52.34173, 
    52.36184, 52.38168, 52.40128, 52.42062, 52.4397, 52.45852, 52.47709, 
    52.49539, 52.51344, 52.53123, 52.54876, 52.56603, 52.58304, 52.59978, 
    52.61628, 52.6325, 52.64847, 52.66417, 52.67962, 52.69479, 52.70971, 
    52.72436, 52.73875, 52.75288, 52.76674, 52.78034, 52.79367, 52.80674, 
    52.81954, 52.83208, 52.84435, 52.85635, 52.86809, 52.87956, 52.89077, 
    52.9017, 52.91238, 52.92278, 52.93291, 52.94278, 52.95238, 52.9617, 
    52.97077, 52.97956, 52.98808, 52.99633, 53.00432, 53.01203, 53.01948, 
    53.02665, 53.03356, 53.04019, 53.04655, 53.05265, 53.05847, 53.06402, 
    53.0693, 53.07431, 53.07904, 53.08351, 53.08771, 53.09163, 53.09528, 
    53.09866, 53.10177, 53.1046, 53.10717, 53.10946, 53.11148, 53.11323, 
    53.1147, 53.11591, 53.11684, 53.1175, 53.11789, 53.118, 53.11784, 
    53.11741, 53.11671, 53.11573, 53.11449, 53.11297, 53.11118, 53.10912, 
    53.10678, 53.10417, 53.1013, 53.09814, 53.09472, 53.09103, 53.08706, 
    53.08282, 53.07831, 53.07353, 53.06848, 53.06316, 53.05756, 53.0517, 
    53.04557, 53.03916, 53.03248, 53.02554, 53.01832, 53.01083, 53.00307, 
    52.99505, 52.98675, 52.97819, 52.96935, 52.96025, 52.95087, 52.94123, 
    52.93133, 52.92115, 52.91071, 52.89999, 52.88901, 52.87777, 52.86625, 
    52.85447, 52.84243, 52.83011, 52.81753, 52.80469, 52.79158, 52.77821, 
    52.76456, 52.75066, 52.7365, 52.72206, 52.70737, 52.69241, 52.67719, 
    52.66171, 52.64596, 52.62995, 52.61369, 52.59715, 52.58036, 52.56331, 
    52.546, 52.52843, 52.5106, 52.49251, 52.47416, 52.45556, 52.4367, 
    52.41758, 52.3982, 52.37856, 52.35867, 52.33853, 52.31812, 52.29747, 
    52.27656, 52.25539, 52.23397, 52.2123, 52.19038, 52.1682, 52.14577, 
    52.1231, 52.10017, 52.07698, 52.05355, 52.02987, 52.00595, 51.98177, 
    51.95734, 51.93267, 51.90775, 51.88258, 51.85717, 51.83151, 51.80561, 
    51.77946, 51.75307, 51.72644, 51.69956, 51.67244, 51.64508, 51.61748, 
    51.58963, 51.56155, 51.53323, 51.50466, 51.47586, 51.44682, 51.41755, 
    51.38803, 51.35828, 51.32829, 51.29807, 51.26762, 51.23692, 51.206, 
    51.17484, 51.14346, 51.11183, 51.07998, 51.0479, 51.01558, 50.98304, 
    50.95027, 50.91727, 50.88404, 50.85059, 50.81691, 50.783, 50.74887, 
    50.71451, 50.67993, 50.64512, 50.6101, 50.57484, 50.53938, 50.50368, 
    50.46777, 50.43164, 50.39529, 50.35872, 50.32193, 50.28492, 50.2477, 
    50.21026, 50.17261, 50.13474, 50.09666, 50.05836, 50.01985, 49.98113, 
    49.9422, 49.90305, 49.8637, 49.82414, 49.78437, 49.74438, 49.7042, 
    49.6638, 49.6232, 49.58239, 49.54137, 49.50016, 49.45874, 49.41711, 
    49.37528, 49.33326,
  44.73399, 44.79205, 44.84998, 44.90776, 44.96539, 45.02288, 45.08022, 
    45.13742, 45.19447, 45.25137, 45.30813, 45.36474, 45.4212, 45.4775, 
    45.53366, 45.58966, 45.64552, 45.70123, 45.75677, 45.81217, 45.86741, 
    45.9225, 45.97743, 46.03221, 46.08683, 46.14129, 46.1956, 46.24975, 
    46.30373, 46.35756, 46.41123, 46.46474, 46.51809, 46.57127, 46.62429, 
    46.67715, 46.72984, 46.78237, 46.83474, 46.88694, 46.93897, 46.99083, 
    47.04253, 47.09406, 47.14542, 47.19661, 47.24763, 47.29848, 47.34915, 
    47.39966, 47.44999, 47.50015, 47.55013, 47.59994, 47.64957, 47.69904, 
    47.74831, 47.79742, 47.84634, 47.89509, 47.94366, 47.99205, 48.04025, 
    48.08828, 48.13612, 48.18378, 48.23126, 48.27856, 48.32567, 48.37259, 
    48.41933, 48.46588, 48.51225, 48.55842, 48.60441, 48.65021, 48.69582, 
    48.74124, 48.78647, 48.8315, 48.87635, 48.921, 48.96545, 49.00972, 
    49.05379, 49.09766, 49.14133, 49.18481, 49.22809, 49.27118, 49.31406, 
    49.35674, 49.39923, 49.44151, 49.48359, 49.52547, 49.56715, 49.60862, 
    49.64989, 49.69095, 49.73181, 49.77246, 49.8129, 49.85314, 49.89317, 
    49.93299, 49.9726, 50.012, 50.05119, 50.09018, 50.12894, 50.1675, 
    50.20584, 50.24397, 50.28188, 50.31958, 50.35706, 50.39433, 50.43137, 
    50.4682, 50.50482, 50.54121, 50.57739, 50.61334, 50.64907, 50.68459, 
    50.71988, 50.75494, 50.78979, 50.82441, 50.8588, 50.89297, 50.92692, 
    50.96064, 50.99413, 51.02739, 51.06043, 51.09324, 51.12581, 51.15816, 
    51.19028, 51.22216, 51.25382, 51.28524, 51.31643, 51.34739, 51.37811, 
    51.40859, 51.43885, 51.46886, 51.49864, 51.52818, 51.55749, 51.58656, 
    51.61539, 51.64397, 51.67233, 51.70044, 51.7283, 51.75593, 51.78332, 
    51.81046, 51.83736, 51.86402, 51.89043, 51.9166, 51.94252, 51.9682, 
    51.99363, 52.01882, 52.04375, 52.06845, 52.09289, 52.11708, 52.14103, 
    52.16472, 52.18817, 52.21136, 52.23431, 52.257, 52.27944, 52.30163, 
    52.32357, 52.34525, 52.36668, 52.38785, 52.40877, 52.42944, 52.44984, 
    52.47, 52.48989, 52.50954, 52.52892, 52.54805, 52.56691, 52.58552, 
    52.60387, 52.62196, 52.63979, 52.65737, 52.67468, 52.69173, 52.70852, 
    52.72505, 52.74131, 52.75732, 52.77306, 52.78854, 52.80376, 52.81871, 
    52.8334, 52.84782, 52.86198, 52.87588, 52.88951, 52.90287, 52.91597, 
    52.92881, 52.94137, 52.95367, 52.96571, 52.97747, 52.98898, 53.00021, 
    53.01117, 53.02187, 53.0323, 53.04245, 53.05235, 53.06197, 53.07132, 
    53.0804, 53.08921, 53.09776, 53.10603, 53.11404, 53.12177, 53.12923, 
    53.13643, 53.14335, 53.15, 53.15638, 53.16248, 53.16832, 53.17389, 
    53.17918, 53.1842, 53.18895, 53.19342, 53.19763, 53.20156, 53.20522, 
    53.20861, 53.21173, 53.21457, 53.21714, 53.21944, 53.22146, 53.22322, 
    53.2247, 53.2259, 53.22684, 53.2275, 53.22789, 53.228, 53.22784, 
    53.22741, 53.22671, 53.22573, 53.22448, 53.22296, 53.22116, 53.21909, 
    53.21675, 53.21414, 53.21125, 53.2081, 53.20466, 53.20096, 53.19698, 
    53.19273, 53.18822, 53.18342, 53.17836, 53.17302, 53.16742, 53.16154, 
    53.15538, 53.14896, 53.14227, 53.13531, 53.12807, 53.12056, 53.11279, 
    53.10474, 53.09643, 53.08784, 53.07898, 53.06986, 53.06046, 53.0508, 
    53.04087, 53.03066, 53.02019, 53.00945, 52.99845, 52.98717, 52.97563, 
    52.96382, 52.95174, 52.9394, 52.92679, 52.91392, 52.90078, 52.88737, 
    52.8737, 52.85976, 52.84556, 52.83109, 52.81636, 52.80136, 52.78611, 
    52.77059, 52.7548, 52.73876, 52.72245, 52.70588, 52.68905, 52.67196, 
    52.65461, 52.63699, 52.61912, 52.60099, 52.5826, 52.56395, 52.54504, 
    52.52587, 52.50645, 52.48677, 52.46683, 52.44663, 52.42619, 52.40548, 
    52.38452, 52.3633, 52.34184, 52.32011, 52.29814, 52.27591, 52.25343, 
    52.23069, 52.20771, 52.18448, 52.16099, 52.13726, 52.11327, 52.08904, 
    52.06456, 52.03983, 52.01485, 51.98962, 51.96415, 51.93844, 51.91248, 
    51.88627, 51.85982, 51.83312, 51.80618, 51.779, 51.75158, 51.72391, 
    51.696, 51.66785, 51.63947, 51.61084, 51.58197, 51.55287, 51.52353, 
    51.49395, 51.46413, 51.43407, 51.40379, 51.37326, 51.3425, 51.31151, 
    51.28028, 51.24883, 51.21714, 51.18521, 51.15306, 51.12067, 51.08806, 
    51.05522, 51.02214, 50.98885, 50.95532, 50.92157, 50.88758, 50.85338, 
    50.81895, 50.78429, 50.74941, 50.71431, 50.67899, 50.64344, 50.60767, 
    50.57168, 50.53547, 50.49904, 50.46239, 50.42553, 50.38845, 50.35115, 
    50.31363, 50.2759, 50.23795, 50.19979, 50.16141, 50.12282, 50.08402, 
    50.04501, 50.00579, 49.96635, 49.92671, 49.88685, 49.84679, 49.80652, 
    49.76604, 49.72536, 49.68447, 49.64337, 49.60207, 49.56057, 49.51886, 
    49.47695, 49.43483,
  44.8273, 44.88546, 44.94347, 45.00134, 45.05906, 45.11664, 45.17408, 
    45.23136, 45.2885, 45.3455, 45.40234, 45.45904, 45.51559, 45.57198, 
    45.62823, 45.68433, 45.74027, 45.79606, 45.8517, 45.90719, 45.96252, 
    46.0177, 46.07272, 46.12759, 46.1823, 46.23685, 46.29125, 46.34549, 
    46.39956, 46.45348, 46.50724, 46.56084, 46.61428, 46.66755, 46.72066, 
    46.77361, 46.82639, 46.87901, 46.93147, 46.98375, 47.03588, 47.08783, 
    47.13962, 47.19123, 47.24269, 47.29396, 47.34507, 47.39601, 47.44678, 
    47.49738, 47.54779, 47.59804, 47.64812, 47.69802, 47.74774, 47.79729, 
    47.84666, 47.89585, 47.94486, 47.9937, 48.04235, 48.09083, 48.13913, 
    48.18724, 48.23518, 48.28292, 48.33049, 48.37787, 48.42507, 48.47208, 
    48.51891, 48.56555, 48.612, 48.65826, 48.70434, 48.75023, 48.79592, 
    48.84143, 48.88674, 48.93187, 48.9768, 49.02153, 49.06607, 49.11042, 
    49.15458, 49.19854, 49.24229, 49.28586, 49.32923, 49.37239, 49.41536, 
    49.45813, 49.5007, 49.54306, 49.58523, 49.62719, 49.66895, 49.71051, 
    49.75186, 49.79301, 49.83395, 49.87468, 49.91521, 49.95553, 49.99564, 
    50.03554, 50.07523, 50.11472, 50.15399, 50.19305, 50.2319, 50.27053, 
    50.30895, 50.34716, 50.38515, 50.42293, 50.46049, 50.49783, 50.53496, 
    50.57187, 50.60856, 50.64503, 50.68128, 50.71731, 50.75312, 50.78871, 
    50.82407, 50.85922, 50.89414, 50.92883, 50.9633, 50.99755, 51.03156, 
    51.06536, 51.09892, 51.13226, 51.16536, 51.19824, 51.23089, 51.26331, 
    51.2955, 51.32746, 51.35918, 51.39067, 51.42193, 51.45295, 51.48375, 
    51.5143, 51.54462, 51.5747, 51.60455, 51.63416, 51.66353, 51.69266, 
    51.72156, 51.75021, 51.77863, 51.8068, 51.83473, 51.86242, 51.88987, 
    51.91708, 51.94404, 51.97076, 51.99723, 52.02346, 52.04944, 52.07518, 
    52.10067, 52.12591, 52.15091, 52.17566, 52.20016, 52.22441, 52.24841, 
    52.27216, 52.29566, 52.31891, 52.3419, 52.36465, 52.38715, 52.40939, 
    52.43137, 52.45311, 52.47459, 52.49581, 52.51678, 52.53749, 52.55795, 
    52.57815, 52.59809, 52.61778, 52.63721, 52.65638, 52.6753, 52.69395, 
    52.71235, 52.73048, 52.74836, 52.76597, 52.78332, 52.80042, 52.81725, 
    52.83381, 52.85012, 52.86616, 52.88194, 52.89746, 52.91271, 52.9277, 
    52.94242, 52.95689, 52.97108, 52.98501, 52.99867, 53.01207, 53.0252, 
    53.03807, 53.05066, 53.063, 53.07506, 53.08685, 53.09838, 53.10964, 
    53.12063, 53.13136, 53.14181, 53.15199, 53.16191, 53.17155, 53.18093, 
    53.19004, 53.19887, 53.20744, 53.21573, 53.22375, 53.23151, 53.23899, 
    53.2462, 53.25314, 53.2598, 53.2662, 53.27232, 53.27817, 53.28375, 
    53.28905, 53.29409, 53.29885, 53.30334, 53.30756, 53.3115, 53.31517, 
    53.31857, 53.32169, 53.32454, 53.32711, 53.32942, 53.33145, 53.33321, 
    53.33469, 53.3359, 53.33683, 53.33749, 53.33788, 53.338, 53.33784, 
    53.33741, 53.3367, 53.33572, 53.33447, 53.33294, 53.33115, 53.32907, 
    53.32673, 53.3241, 53.32121, 53.31805, 53.31461, 53.31089, 53.30691, 
    53.30265, 53.29811, 53.29331, 53.28823, 53.28289, 53.27726, 53.27137, 
    53.26521, 53.25877, 53.25206, 53.24508, 53.23782, 53.2303, 53.2225, 
    53.21444, 53.2061, 53.19749, 53.18861, 53.17947, 53.17005, 53.16036, 
    53.1504, 53.14017, 53.12968, 53.11891, 53.10788, 53.09658, 53.08501, 
    53.07317, 53.06106, 53.04869, 53.03605, 53.02314, 53.00997, 52.99653, 
    52.98282, 52.96885, 52.95462, 52.94011, 52.92535, 52.91032, 52.89502, 
    52.87946, 52.86364, 52.84756, 52.83121, 52.8146, 52.79773, 52.78059, 
    52.7632, 52.74554, 52.72763, 52.70945, 52.69102, 52.67232, 52.65337, 
    52.63416, 52.61469, 52.59496, 52.57497, 52.55473, 52.53423, 52.51348, 
    52.49247, 52.4712, 52.44968, 52.42791, 52.40588, 52.3836, 52.36107, 
    52.33828, 52.31525, 52.29196, 52.26842, 52.24463, 52.22058, 52.1963, 
    52.17176, 52.14697, 52.12194, 52.09665, 52.07112, 52.04535, 52.01933, 
    51.99306, 51.96655, 51.93979, 51.91279, 51.88554, 51.85806, 51.83033, 
    51.80236, 51.77415, 51.74569, 51.717, 51.68807, 51.6589, 51.62949, 
    51.59984, 51.56996, 51.53984, 51.50948, 51.47889, 51.44806, 51.417, 
    51.38571, 51.35418, 51.32242, 51.29042, 51.2582, 51.22574, 51.19306, 
    51.16014, 51.127, 51.09363, 51.06002, 51.0262, 50.99215, 50.95786, 
    50.92336, 50.88863, 50.85368, 50.8185, 50.7831, 50.74747, 50.71163, 
    50.67556, 50.63927, 50.60277, 50.56604, 50.5291, 50.49194, 50.45456, 
    50.41697, 50.37915, 50.34113, 50.30289, 50.26443, 50.22577, 50.18688, 
    50.14779, 50.10848, 50.06897, 50.02924, 49.98931, 49.94916, 49.90881, 
    49.86825, 49.82748, 49.78651, 49.74533, 49.70395, 49.66236, 49.62057, 
    49.57858, 49.53638,
  44.92057, 44.97881, 45.03691, 45.09487, 45.15268, 45.21035, 45.26787, 
    45.32525, 45.38248, 45.43956, 45.49649, 45.55328, 45.60992, 45.66641, 
    45.72274, 45.77893, 45.83496, 45.89085, 45.94658, 46.00216, 46.05758, 
    46.11285, 46.16796, 46.22292, 46.27771, 46.33236, 46.38684, 46.44117, 
    46.49534, 46.54935, 46.6032, 46.65689, 46.71041, 46.76377, 46.81698, 
    46.87002, 46.92289, 46.9756, 47.02814, 47.08052, 47.13274, 47.18478, 
    47.23666, 47.28836, 47.3399, 47.39127, 47.44247, 47.4935, 47.54436, 
    47.59504, 47.64555, 47.69589, 47.74605, 47.79604, 47.84586, 47.89549, 
    47.94495, 47.99423, 48.04333, 48.09226, 48.14101, 48.18957, 48.23796, 
    48.28616, 48.33418, 48.38202, 48.42967, 48.47714, 48.52443, 48.57153, 
    48.61844, 48.66517, 48.71171, 48.75806, 48.80423, 48.8502, 48.89598, 
    48.94158, 48.98698, 49.03219, 49.07721, 49.12203, 49.16666, 49.21109, 
    49.25533, 49.29937, 49.34322, 49.38687, 49.43032, 49.47358, 49.51663, 
    49.55948, 49.60213, 49.64458, 49.68683, 49.72888, 49.77073, 49.81236, 
    49.8538, 49.89503, 49.93605, 49.97687, 50.01748, 50.05788, 50.09807, 
    50.13806, 50.17783, 50.2174, 50.25675, 50.29589, 50.33482, 50.37353, 
    50.41203, 50.45032, 50.48839, 50.52625, 50.56389, 50.60131, 50.63852, 
    50.6755, 50.71227, 50.74882, 50.78515, 50.82125, 50.85714, 50.89281, 
    50.92825, 50.96347, 50.99846, 51.03323, 51.06778, 51.10209, 51.13618, 
    51.17005, 51.20369, 51.2371, 51.27028, 51.30323, 51.33595, 51.36844, 
    51.4007, 51.43273, 51.46452, 51.49608, 51.52741, 51.5585, 51.58936, 
    51.61999, 51.65037, 51.68052, 51.71044, 51.74011, 51.76955, 51.79875, 
    51.82771, 51.85643, 51.88491, 51.91314, 51.94114, 51.96889, 51.99641, 
    52.02367, 52.0507, 52.07748, 52.10401, 52.1303, 52.15634, 52.18214, 
    52.20769, 52.23299, 52.25805, 52.28285, 52.30741, 52.33171, 52.35577, 
    52.37958, 52.40313, 52.42644, 52.44949, 52.47229, 52.49483, 52.51713, 
    52.53917, 52.56096, 52.58249, 52.60376, 52.62478, 52.64554, 52.66605, 
    52.6863, 52.70629, 52.72602, 52.7455, 52.76472, 52.78367, 52.80237, 
    52.82081, 52.83899, 52.85691, 52.87457, 52.89196, 52.90909, 52.92596, 
    52.94257, 52.95892, 52.975, 52.99082, 53.00637, 53.02166, 53.03669, 
    53.05145, 53.06594, 53.08017, 53.09414, 53.10783, 53.12127, 53.13443, 
    53.14732, 53.15995, 53.17231, 53.18441, 53.19623, 53.20779, 53.21907, 
    53.23009, 53.24084, 53.25132, 53.26153, 53.27147, 53.28114, 53.29054, 
    53.29967, 53.30853, 53.31711, 53.32543, 53.33347, 53.34124, 53.34874, 
    53.35597, 53.36293, 53.36961, 53.37602, 53.38216, 53.38802, 53.39362, 
    53.39893, 53.40398, 53.40875, 53.41325, 53.41748, 53.42143, 53.42511, 
    53.42852, 53.43165, 53.43451, 53.43709, 53.4394, 53.44143, 53.44319, 
    53.44468, 53.44589, 53.44683, 53.44749, 53.44788, 53.448, 53.44784, 
    53.44741, 53.4467, 53.44572, 53.44446, 53.44293, 53.44113, 53.43905, 
    53.4367, 53.43407, 53.43117, 53.42799, 53.42455, 53.42083, 53.41683, 
    53.41256, 53.40802, 53.4032, 53.39811, 53.39275, 53.38711, 53.3812, 
    53.37502, 53.36857, 53.36184, 53.35484, 53.34757, 53.34003, 53.33221, 
    53.32413, 53.31577, 53.30714, 53.29824, 53.28907, 53.27963, 53.26992, 
    53.25993, 53.24968, 53.23916, 53.22837, 53.21731, 53.20598, 53.19438, 
    53.18251, 53.17038, 53.15797, 53.1453, 53.13236, 53.11916, 53.10568, 
    53.09195, 53.07794, 53.06367, 53.04913, 53.03433, 53.01926, 53.00393, 
    52.98833, 52.97247, 52.95635, 52.93996, 52.92331, 52.9064, 52.88923, 
    52.87179, 52.85409, 52.83613, 52.81791, 52.79943, 52.78069, 52.76169, 
    52.74244, 52.72292, 52.70314, 52.68311, 52.66282, 52.64227, 52.62147, 
    52.60041, 52.57909, 52.55753, 52.5357, 52.51362, 52.49129, 52.4687, 
    52.44586, 52.42277, 52.39943, 52.37583, 52.35198, 52.32789, 52.30354, 
    52.27895, 52.2541, 52.22901, 52.20366, 52.17808, 52.15224, 52.12616, 
    52.09983, 52.07326, 52.04644, 52.01937, 51.99207, 51.96452, 51.93673, 
    51.9087, 51.88042, 51.8519, 51.82314, 51.79415, 51.76491, 51.73544, 
    51.70572, 51.67577, 51.64558, 51.61516, 51.5845, 51.5536, 51.52247, 
    51.4911, 51.45951, 51.42768, 51.39561, 51.36332, 51.33079, 51.29803, 
    51.26505, 51.23183, 51.19838, 51.16471, 51.13081, 51.09668, 51.06232, 
    51.02774, 50.99294, 50.95791, 50.92266, 50.88718, 50.85148, 50.81556, 
    50.77942, 50.74305, 50.70647, 50.66967, 50.63264, 50.59541, 50.55795, 
    50.52028, 50.48238, 50.44428, 50.40596, 50.36742, 50.32867, 50.28971, 
    50.25054, 50.21115, 50.17155, 50.13174, 50.09173, 50.0515, 50.01107, 
    49.97042, 49.92958, 49.88852, 49.84726, 49.80579, 49.76412, 49.72224, 
    49.68016, 49.63788,
  45.01376, 45.0721, 45.13029, 45.18834, 45.24624, 45.304, 45.36161, 
    45.41908, 45.47639, 45.53357, 45.59059, 45.64747, 45.7042, 45.76077, 
    45.8172, 45.87348, 45.9296, 45.98558, 46.0414, 46.09706, 46.15258, 
    46.20794, 46.26314, 46.31818, 46.37308, 46.42781, 46.48239, 46.5368, 
    46.59106, 46.64516, 46.6991, 46.75288, 46.8065, 46.85995, 46.91324, 
    46.96637, 47.01934, 47.07214, 47.12477, 47.17724, 47.22954, 47.28168, 
    47.33364, 47.38544, 47.43707, 47.48853, 47.53982, 47.59094, 47.64189, 
    47.69266, 47.74326, 47.79369, 47.84394, 47.89402, 47.94392, 47.99365, 
    48.0432, 48.09257, 48.14176, 48.19078, 48.23961, 48.28827, 48.33674, 
    48.38503, 48.43314, 48.48107, 48.52881, 48.57637, 48.62374, 48.67093, 
    48.71793, 48.76475, 48.81138, 48.85782, 48.90407, 48.95013, 48.996, 
    49.04168, 49.08717, 49.13247, 49.17757, 49.22248, 49.2672, 49.31172, 
    49.35604, 49.40017, 49.44411, 49.48784, 49.53138, 49.57471, 49.61786, 
    49.66079, 49.70353, 49.74607, 49.7884, 49.83053, 49.87246, 49.91418, 
    49.9557, 49.99701, 50.03812, 50.07902, 50.11971, 50.1602, 50.20047, 
    50.24054, 50.2804, 50.32004, 50.35947, 50.3987, 50.43771, 50.4765, 
    50.51508, 50.55345, 50.5916, 50.62954, 50.66726, 50.70476, 50.74204, 
    50.77911, 50.81595, 50.85258, 50.88898, 50.92517, 50.96114, 50.99688, 
    51.03239, 51.06769, 51.10276, 51.1376, 51.17222, 51.20662, 51.24078, 
    51.27472, 51.30843, 51.34192, 51.37517, 51.40819, 51.44098, 51.47355, 
    51.50587, 51.53798, 51.56984, 51.60147, 51.63287, 51.66403, 51.69496, 
    51.72565, 51.75611, 51.78632, 51.81631, 51.84605, 51.87555, 51.90482, 
    51.93384, 51.96263, 51.99117, 52.01947, 52.04753, 52.07535, 52.10292, 
    52.13026, 52.15734, 52.18418, 52.21078, 52.23713, 52.26323, 52.28909, 
    52.3147, 52.34006, 52.36517, 52.39003, 52.41465, 52.43901, 52.46312, 
    52.48699, 52.5106, 52.53396, 52.55706, 52.57992, 52.60252, 52.62486, 
    52.64695, 52.66879, 52.69037, 52.7117, 52.73277, 52.75358, 52.77414, 
    52.79443, 52.81447, 52.83425, 52.85378, 52.87304, 52.89204, 52.91079, 
    52.92927, 52.94749, 52.96545, 52.98315, 53.00059, 53.01777, 53.03468, 
    53.05132, 53.06771, 53.08383, 53.09969, 53.11528, 53.13061, 53.14567, 
    53.16047, 53.175, 53.18926, 53.20326, 53.21699, 53.23045, 53.24365, 
    53.25658, 53.26924, 53.28163, 53.29375, 53.30561, 53.31719, 53.32851, 
    53.33955, 53.35033, 53.36083, 53.37107, 53.38103, 53.39072, 53.40015, 
    53.4093, 53.41818, 53.42678, 53.43512, 53.44318, 53.45097, 53.45849, 
    53.46574, 53.47271, 53.47941, 53.48584, 53.49199, 53.49787, 53.50348, 
    53.50881, 53.51387, 53.51865, 53.52317, 53.5274, 53.53136, 53.53505, 
    53.53847, 53.54161, 53.54447, 53.54706, 53.54937, 53.55141, 53.55318, 
    53.55467, 53.55589, 53.55683, 53.55749, 53.55788, 53.558, 53.55784, 
    53.55741, 53.5567, 53.55571, 53.55445, 53.55292, 53.55111, 53.54903, 
    53.54667, 53.54404, 53.54113, 53.53794, 53.53449, 53.53076, 53.52675, 
    53.52247, 53.51792, 53.51309, 53.50799, 53.50261, 53.49696, 53.49104, 
    53.48484, 53.47837, 53.47163, 53.46461, 53.45732, 53.44976, 53.44193, 
    53.43382, 53.42544, 53.41679, 53.40787, 53.39867, 53.38921, 53.37947, 
    53.36946, 53.35919, 53.34864, 53.33782, 53.32673, 53.31538, 53.30375, 
    53.29185, 53.27969, 53.26725, 53.25455, 53.24158, 53.22834, 53.21484, 
    53.20106, 53.18702, 53.17272, 53.15814, 53.14331, 53.1282, 53.11283, 
    53.0972, 53.0813, 53.06514, 53.04871, 53.03202, 53.01506, 52.99785, 
    52.98037, 52.96263, 52.94463, 52.92636, 52.90784, 52.88905, 52.87001, 
    52.8507, 52.83114, 52.81132, 52.79124, 52.7709, 52.75031, 52.72945, 
    52.70834, 52.68697, 52.66535, 52.64347, 52.62135, 52.59896, 52.57632, 
    52.55342, 52.53028, 52.50688, 52.48323, 52.45933, 52.43517, 52.41077, 
    52.38612, 52.36121, 52.33606, 52.31066, 52.28502, 52.25912, 52.23298, 
    52.20659, 52.17995, 52.15307, 52.12595, 52.09858, 52.07096, 52.04311, 
    52.01501, 51.98667, 51.95809, 51.92927, 51.9002, 51.8709, 51.84136, 
    51.81158, 51.78156, 51.7513, 51.72081, 51.69008, 51.65912, 51.62792, 
    51.59648, 51.56482, 51.53291, 51.50078, 51.46841, 51.43581, 51.40298, 
    51.36992, 51.33663, 51.30311, 51.26937, 51.23539, 51.20119, 51.16676, 
    51.1321, 51.09723, 51.06212, 51.02679, 50.99124, 50.95546, 50.91946, 
    50.88324, 50.8468, 50.81014, 50.77326, 50.73616, 50.69884, 50.6613, 
    50.62355, 50.58558, 50.54739, 50.509, 50.47038, 50.43155, 50.39251, 
    50.35325, 50.31378, 50.27411, 50.23421, 50.19411, 50.15381, 50.11329, 
    50.07256, 50.03163, 49.99049, 49.94915, 49.9076, 49.86584, 49.82388, 
    49.78172, 49.73935,
  45.1069, 45.16533, 45.22361, 45.28175, 45.33974, 45.39759, 45.45529, 
    45.51284, 45.57026, 45.62752, 45.68463, 45.7416, 45.79842, 45.85508, 
    45.9116, 45.96797, 46.02419, 46.08025, 46.13616, 46.19192, 46.24752, 
    46.30297, 46.35826, 46.4134, 46.46838, 46.5232, 46.57787, 46.63238, 
    46.68673, 46.74092, 46.79495, 46.84882, 46.90253, 46.95607, 47.00945, 
    47.06268, 47.11573, 47.16862, 47.22134, 47.2739, 47.3263, 47.37852, 
    47.43058, 47.48247, 47.53419, 47.58574, 47.63712, 47.68833, 47.73936, 
    47.79023, 47.84092, 47.89144, 47.94178, 47.99195, 48.04194, 48.09176, 
    48.1414, 48.19086, 48.24014, 48.28925, 48.33817, 48.38691, 48.43547, 
    48.48386, 48.53205, 48.58007, 48.6279, 48.67555, 48.72301, 48.77029, 
    48.81738, 48.86429, 48.911, 48.95753, 49.00387, 49.05002, 49.09598, 
    49.14175, 49.18732, 49.23271, 49.2779, 49.3229, 49.3677, 49.4123, 
    49.45672, 49.50093, 49.54495, 49.58878, 49.6324, 49.67582, 49.71904, 
    49.76207, 49.80489, 49.84751, 49.88993, 49.93215, 49.97416, 50.01596, 
    50.05757, 50.09896, 50.14016, 50.18114, 50.22191, 50.26248, 50.30284, 
    50.34299, 50.38293, 50.42265, 50.46217, 50.50147, 50.54056, 50.57944, 
    50.6181, 50.65655, 50.69478, 50.7328, 50.7706, 50.80818, 50.84554, 
    50.88268, 50.91961, 50.95631, 50.9928, 51.02906, 51.0651, 51.10092, 
    51.13651, 51.17188, 51.20703, 51.24195, 51.27664, 51.31111, 51.34535, 
    51.37936, 51.41315, 51.4467, 51.48003, 51.51313, 51.54599, 51.57863, 
    51.61103, 51.6432, 51.67514, 51.70684, 51.7383, 51.76954, 51.80053, 
    51.8313, 51.86182, 51.89211, 51.92215, 51.95197, 51.98154, 52.01087, 
    52.03996, 52.06881, 52.09742, 52.12579, 52.15391, 52.18179, 52.20943, 
    52.23682, 52.26397, 52.29087, 52.31753, 52.34394, 52.37011, 52.39602, 
    52.42169, 52.44711, 52.47228, 52.4972, 52.52187, 52.5463, 52.57047, 
    52.59438, 52.61805, 52.64146, 52.66462, 52.68753, 52.71019, 52.73258, 
    52.75473, 52.77662, 52.79825, 52.81963, 52.84074, 52.86161, 52.88221, 
    52.90256, 52.92265, 52.94247, 52.96204, 52.98135, 53.0004, 53.01919, 
    53.03772, 53.05599, 53.07399, 53.09173, 53.10921, 53.12643, 53.14338, 
    53.16007, 53.17649, 53.19266, 53.20855, 53.22418, 53.23955, 53.25465, 
    53.26948, 53.28405, 53.29834, 53.31238, 53.32614, 53.33964, 53.35287, 
    53.36583, 53.37852, 53.39094, 53.40309, 53.41498, 53.42659, 53.43793, 
    53.44901, 53.45981, 53.47034, 53.4806, 53.49059, 53.50031, 53.50975, 
    53.51892, 53.52783, 53.53646, 53.54481, 53.55289, 53.56071, 53.56824, 
    53.57551, 53.5825, 53.58921, 53.59566, 53.60183, 53.60772, 53.61334, 
    53.61869, 53.62376, 53.62856, 53.63308, 53.63733, 53.6413, 53.645, 
    53.64842, 53.65157, 53.65443, 53.65703, 53.65935, 53.6614, 53.66317, 
    53.66466, 53.66588, 53.66682, 53.66749, 53.66788, 53.668, 53.66784, 
    53.6674, 53.66669, 53.66571, 53.66444, 53.66291, 53.66109, 53.659, 
    53.65664, 53.654, 53.65108, 53.6479, 53.64443, 53.64069, 53.63667, 
    53.63238, 53.62782, 53.62297, 53.61786, 53.61247, 53.60681, 53.60087, 
    53.59466, 53.58817, 53.58141, 53.57438, 53.56707, 53.55949, 53.55164, 
    53.54351, 53.53511, 53.52644, 53.51749, 53.50828, 53.49879, 53.48903, 
    53.479, 53.46869, 53.45812, 53.44727, 53.43616, 53.42477, 53.41312, 
    53.40119, 53.38899, 53.37653, 53.3638, 53.35079, 53.33752, 53.32398, 
    53.31018, 53.2961, 53.28176, 53.26715, 53.25228, 53.23714, 53.22173, 
    53.20605, 53.19012, 53.17392, 53.15745, 53.14072, 53.12372, 53.10646, 
    53.08894, 53.07116, 53.05312, 53.03481, 53.01624, 52.99741, 52.97832, 
    52.95897, 52.93935, 52.91949, 52.89936, 52.87897, 52.85832, 52.83742, 
    52.81626, 52.79485, 52.77317, 52.75124, 52.72906, 52.70662, 52.68393, 
    52.66098, 52.63778, 52.61432, 52.59062, 52.56666, 52.54245, 52.51799, 
    52.49327, 52.46832, 52.4431, 52.41764, 52.39194, 52.36598, 52.33978, 
    52.31333, 52.28663, 52.25969, 52.2325, 52.20507, 52.17739, 52.14948, 
    52.12132, 52.09291, 52.06426, 52.03537, 52.00624, 51.97688, 51.94727, 
    51.91742, 51.88733, 51.85701, 51.82645, 51.79565, 51.76461, 51.73334, 
    51.70184, 51.6701, 51.63813, 51.60592, 51.57348, 51.54081, 51.50791, 
    51.47478, 51.44141, 51.40782, 51.374, 51.33995, 51.30567, 51.27117, 
    51.23644, 51.20148, 51.1663, 51.13089, 51.09526, 51.05941, 51.02334, 
    50.98704, 50.95052, 50.91378, 50.87682, 50.83965, 50.80225, 50.76463, 
    50.7268, 50.68875, 50.65048, 50.612, 50.5733, 50.53439, 50.49527, 
    50.45593, 50.41638, 50.37662, 50.33665, 50.29647, 50.25608, 50.21548, 
    50.17467, 50.13365, 50.09243, 50.051, 50.00937, 49.96753, 49.92548, 
    49.88324, 49.84078,
  45.19999, 45.2585, 45.31687, 45.3751, 45.43318, 45.49112, 45.54891, 
    45.60656, 45.66405, 45.72141, 45.77861, 45.83567, 45.89258, 45.94934, 
    46.00594, 46.0624, 46.11871, 46.17486, 46.23086, 46.28671, 46.34241, 
    46.39795, 46.45333, 46.50856, 46.56363, 46.61855, 46.67331, 46.7279, 
    46.78234, 46.83662, 46.89074, 46.94471, 46.9985, 47.05214, 47.10561, 
    47.15892, 47.21207, 47.26505, 47.31787, 47.37052, 47.423, 47.47532, 
    47.52747, 47.57944, 47.63126, 47.6829, 47.73437, 47.78567, 47.8368, 
    47.88775, 47.93853, 47.98914, 48.03957, 48.08983, 48.13991, 48.18982, 
    48.23955, 48.2891, 48.33847, 48.38766, 48.43668, 48.48551, 48.53416, 
    48.58264, 48.63092, 48.67903, 48.72695, 48.77469, 48.82224, 48.86961, 
    48.91679, 48.96378, 49.01059, 49.0572, 49.10363, 49.14986, 49.19591, 
    49.24177, 49.28743, 49.3329, 49.37818, 49.42327, 49.46816, 49.51285, 
    49.55735, 49.60165, 49.64576, 49.68967, 49.73338, 49.77689, 49.82019, 
    49.8633, 49.90621, 49.94892, 49.99142, 50.03373, 50.07582, 50.11771, 
    50.1594, 50.20088, 50.24215, 50.28322, 50.32408, 50.36473, 50.40517, 
    50.4454, 50.48542, 50.52523, 50.56483, 50.60422, 50.64339, 50.68235, 
    50.72109, 50.75962, 50.79793, 50.83603, 50.87391, 50.91156, 50.94901, 
    50.98623, 51.02323, 51.06002, 51.09658, 51.13292, 51.16904, 51.20493, 
    51.2406, 51.27605, 51.31127, 51.34627, 51.38103, 51.41558, 51.4499, 
    51.48398, 51.51784, 51.55147, 51.58487, 51.61804, 51.65098, 51.68369, 
    51.71616, 51.7484, 51.78041, 51.81218, 51.84372, 51.87502, 51.90609, 
    51.93692, 51.96751, 51.99787, 52.02798, 52.05786, 52.0875, 52.1169, 
    52.14606, 52.17497, 52.20364, 52.23208, 52.26027, 52.28821, 52.31591, 
    52.34337, 52.37058, 52.39754, 52.42426, 52.45074, 52.47696, 52.50294, 
    52.52867, 52.55415, 52.57938, 52.60435, 52.62909, 52.65356, 52.67779, 
    52.70177, 52.72549, 52.74896, 52.77217, 52.79514, 52.81784, 52.84029, 
    52.86249, 52.88443, 52.90612, 52.92754, 52.94871, 52.96962, 52.99028, 
    53.01067, 53.03081, 53.05069, 53.0703, 53.08966, 53.10876, 53.12759, 
    53.14616, 53.16447, 53.18252, 53.20031, 53.21783, 53.23509, 53.25208, 
    53.26881, 53.28528, 53.30148, 53.31741, 53.33308, 53.34848, 53.36362, 
    53.37849, 53.39309, 53.40742, 53.42149, 53.43529, 53.44882, 53.46208, 
    53.47507, 53.4878, 53.50025, 53.51243, 53.52435, 53.53599, 53.54736, 
    53.55846, 53.56929, 53.57985, 53.59013, 53.60014, 53.60989, 53.61935, 
    53.62855, 53.63748, 53.64613, 53.6545, 53.66261, 53.67044, 53.67799, 
    53.68528, 53.69228, 53.69902, 53.70547, 53.71166, 53.71757, 53.72321, 
    53.72857, 53.73365, 53.73846, 53.74299, 53.74725, 53.75123, 53.75494, 
    53.75837, 53.76152, 53.7644, 53.76701, 53.76933, 53.77138, 53.77316, 
    53.77465, 53.77588, 53.77682, 53.77749, 53.77788, 53.778, 53.77784, 
    53.7774, 53.77669, 53.7757, 53.77444, 53.77289, 53.77108, 53.76898, 
    53.76661, 53.76397, 53.76104, 53.75784, 53.75437, 53.75062, 53.74659, 
    53.74229, 53.73772, 53.73286, 53.72773, 53.72233, 53.71665, 53.7107, 
    53.70447, 53.69797, 53.69119, 53.68414, 53.67682, 53.66922, 53.66134, 
    53.6532, 53.64478, 53.63608, 53.62712, 53.61788, 53.60836, 53.59858, 
    53.58852, 53.57819, 53.56759, 53.55672, 53.54558, 53.53416, 53.52248, 
    53.51052, 53.49829, 53.4858, 53.47303, 53.46, 53.4467, 53.43312, 
    53.41928, 53.40517, 53.3908, 53.37615, 53.36124, 53.34607, 53.33062, 
    53.31491, 53.29893, 53.28269, 53.26618, 53.24941, 53.23238, 53.21508, 
    53.19751, 53.17968, 53.16159, 53.14324, 53.12463, 53.10575, 53.08662, 
    53.06722, 53.04756, 53.02764, 53.00747, 52.98703, 52.96634, 52.94538, 
    52.92417, 52.9027, 52.88098, 52.859, 52.83676, 52.81427, 52.79152, 
    52.76852, 52.74526, 52.72175, 52.69799, 52.67398, 52.64971, 52.62519, 
    52.60042, 52.5754, 52.55013, 52.52461, 52.49884, 52.47283, 52.44656, 
    52.42006, 52.3933, 52.36629, 52.33904, 52.31155, 52.28381, 52.25583, 
    52.2276, 52.19913, 52.17041, 52.14146, 52.11226, 52.08283, 52.05315, 
    52.02324, 51.99308, 51.96269, 51.93206, 51.90119, 51.87009, 51.83875, 
    51.80717, 51.77536, 51.74332, 51.71104, 51.67853, 51.64579, 51.61281, 
    51.57961, 51.54617, 51.5125, 51.47861, 51.44448, 51.41013, 51.37555, 
    51.34074, 51.30571, 51.27045, 51.23497, 51.19927, 51.16334, 51.12719, 
    51.09081, 51.05421, 51.0174, 50.98036, 50.9431, 50.90562, 50.86793, 
    50.83001, 50.79188, 50.75354, 50.71497, 50.6762, 50.63721, 50.598, 
    50.55858, 50.51895, 50.47911, 50.43905, 50.39879, 50.35831, 50.31763, 
    50.27674, 50.23564, 50.19433, 50.15282, 50.1111, 50.06918, 50.02705, 
    49.98471, 49.94218,
  45.293, 45.35161, 45.41007, 45.46838, 45.52656, 45.58459, 45.64247, 
    45.70021, 45.7578, 45.81524, 45.87254, 45.92968, 45.98668, 46.04353, 
    46.10023, 46.15678, 46.21317, 46.26942, 46.32551, 46.38145, 46.43724, 
    46.49287, 46.54834, 46.60366, 46.65882, 46.71383, 46.76868, 46.82337, 
    46.8779, 46.93227, 46.98648, 47.04053, 47.09443, 47.14816, 47.20172, 
    47.25512, 47.30836, 47.36143, 47.41434, 47.46708, 47.51965, 47.57206, 
    47.6243, 47.67637, 47.72827, 47.78, 47.83157, 47.88295, 47.93417, 
    47.98522, 48.03609, 48.08679, 48.13731, 48.18766, 48.23783, 48.28783, 
    48.33765, 48.38729, 48.43676, 48.48604, 48.53514, 48.58407, 48.63281, 
    48.68137, 48.72975, 48.77794, 48.82595, 48.87378, 48.92142, 48.96888, 
    49.01614, 49.06323, 49.11012, 49.15683, 49.20334, 49.24967, 49.2958, 
    49.34175, 49.3875, 49.43306, 49.47842, 49.5236, 49.56858, 49.61336, 
    49.65794, 49.70234, 49.74652, 49.79052, 49.83432, 49.87791, 49.92131, 
    49.9645, 50.0075, 50.05029, 50.09288, 50.13527, 50.17744, 50.21942, 
    50.2612, 50.30276, 50.34412, 50.38527, 50.42621, 50.46695, 50.50747, 
    50.54778, 50.58789, 50.62778, 50.66746, 50.70693, 50.74618, 50.78522, 
    50.82404, 50.86265, 50.90105, 50.93922, 50.97718, 51.01492, 51.05244, 
    51.08974, 51.12683, 51.16369, 51.20033, 51.23675, 51.27295, 51.30892, 
    51.34467, 51.38019, 51.41549, 51.45056, 51.4854, 51.52002, 51.55442, 
    51.58858, 51.62251, 51.65622, 51.68969, 51.72293, 51.75594, 51.78872, 
    51.82127, 51.85358, 51.88566, 51.9175, 51.94911, 51.98048, 52.01162, 
    52.04252, 52.07318, 52.10361, 52.13379, 52.16374, 52.19344, 52.22291, 
    52.25213, 52.28112, 52.30986, 52.33835, 52.3666, 52.39462, 52.42238, 
    52.4499, 52.47717, 52.5042, 52.53098, 52.55752, 52.5838, 52.60984, 
    52.63563, 52.66117, 52.68646, 52.71149, 52.73628, 52.76082, 52.7851, 
    52.80914, 52.83291, 52.85644, 52.87971, 52.90273, 52.92549, 52.94799, 
    52.97024, 52.99223, 53.01397, 53.03545, 53.05667, 53.07763, 53.09834, 
    53.11878, 53.13897, 53.15889, 53.17855, 53.19796, 53.2171, 53.23598, 
    53.2546, 53.27295, 53.29105, 53.30887, 53.32644, 53.34374, 53.36077, 
    53.37754, 53.39405, 53.41029, 53.42627, 53.44197, 53.45741, 53.47258, 
    53.48749, 53.50213, 53.5165, 53.5306, 53.54443, 53.55799, 53.57129, 
    53.58432, 53.59707, 53.60955, 53.62177, 53.63371, 53.64538, 53.65678, 
    53.66791, 53.67876, 53.68935, 53.69966, 53.7097, 53.71946, 53.72896, 
    53.73818, 53.74712, 53.75579, 53.76419, 53.77232, 53.78017, 53.78774, 
    53.79504, 53.80207, 53.80882, 53.81529, 53.8215, 53.82742, 53.83307, 
    53.83844, 53.84354, 53.84836, 53.8529, 53.85717, 53.86116, 53.86488, 
    53.86832, 53.87148, 53.87437, 53.87698, 53.87931, 53.88137, 53.88314, 
    53.88465, 53.88587, 53.88682, 53.88749, 53.88788, 53.888, 53.88784, 
    53.8874, 53.88669, 53.8857, 53.88443, 53.88288, 53.88106, 53.87896, 
    53.87658, 53.87393, 53.871, 53.86779, 53.86431, 53.86055, 53.85651, 
    53.8522, 53.84761, 53.84275, 53.83761, 53.83219, 53.8265, 53.82053, 
    53.81429, 53.80777, 53.80098, 53.79391, 53.78656, 53.77894, 53.77105, 
    53.76288, 53.75444, 53.74573, 53.73674, 53.72747, 53.71794, 53.70813, 
    53.69805, 53.68769, 53.67706, 53.66616, 53.65499, 53.64355, 53.63184, 
    53.61985, 53.6076, 53.59507, 53.58227, 53.56921, 53.55587, 53.54226, 
    53.52839, 53.51424, 53.49983, 53.48515, 53.4702, 53.45499, 53.43951, 
    53.42376, 53.40774, 53.39146, 53.37491, 53.3581, 53.34102, 53.32368, 
    53.30607, 53.2882, 53.27007, 53.25167, 53.23301, 53.21409, 53.19491, 
    53.17546, 53.15576, 53.13579, 53.11557, 53.09508, 53.07433, 53.05333, 
    53.03207, 53.01055, 52.98877, 52.96674, 52.94445, 52.9219, 52.8991, 
    52.87605, 52.85273, 52.82917, 52.80535, 52.78128, 52.75695, 52.73238, 
    52.70755, 52.68247, 52.65715, 52.63157, 52.60574, 52.57966, 52.55334, 
    52.52676, 52.49994, 52.47288, 52.44556, 52.418, 52.3902, 52.36215, 
    52.33386, 52.30532, 52.27655, 52.24753, 52.21827, 52.18876, 52.15902, 
    52.12904, 52.09881, 52.06835, 52.03765, 52.00671, 51.97554, 51.94413, 
    51.91248, 51.8806, 51.84848, 51.81614, 51.78355, 51.75074, 51.71769, 
    51.68441, 51.6509, 51.61716, 51.58319, 51.54899, 51.51456, 51.47991, 
    51.44503, 51.40992, 51.37458, 51.33902, 51.30324, 51.26723, 51.231, 
    51.19455, 51.15788, 51.12098, 51.08386, 51.04652, 51.00897, 50.97119, 
    50.9332, 50.89499, 50.85656, 50.81792, 50.77906, 50.73999, 50.7007, 
    50.6612, 50.62148, 50.58156, 50.54142, 50.50108, 50.46052, 50.41975, 
    50.37877, 50.33759, 50.2962, 50.2546, 50.2128, 50.17079, 50.12857, 
    50.08615, 50.04353,
  45.38596, 45.44466, 45.50321, 45.56161, 45.61988, 45.67799, 45.73597, 
    45.7938, 45.85148, 45.90901, 45.9664, 46.02364, 46.08073, 46.13766, 
    46.19445, 46.25109, 46.30758, 46.36392, 46.4201, 46.47613, 46.53201, 
    46.58773, 46.6433, 46.69871, 46.75396, 46.80906, 46.864, 46.91878, 
    46.9734, 47.02787, 47.08217, 47.13631, 47.19029, 47.24411, 47.29777, 
    47.35126, 47.40459, 47.45775, 47.51075, 47.56358, 47.61625, 47.66875, 
    47.72108, 47.77324, 47.82523, 47.87706, 47.92871, 47.98019, 48.0315, 
    48.08264, 48.1336, 48.18439, 48.235, 48.28544, 48.33571, 48.3858, 
    48.4357, 48.48544, 48.53499, 48.58437, 48.63356, 48.68257, 48.73141, 
    48.78006, 48.82853, 48.87681, 48.92491, 48.97282, 49.02056, 49.0681, 
    49.11546, 49.16263, 49.20961, 49.25641, 49.30301, 49.34943, 49.39565, 
    49.44168, 49.48753, 49.53317, 49.57863, 49.62389, 49.66895, 49.71382, 
    49.7585, 49.80297, 49.84725, 49.89133, 49.93521, 49.9789, 50.02238, 
    50.06566, 50.10875, 50.15162, 50.1943, 50.23677, 50.27903, 50.3211, 
    50.36295, 50.4046, 50.44604, 50.48728, 50.52831, 50.56913, 50.60973, 
    50.65013, 50.69032, 50.73029, 50.77005, 50.8096, 50.84894, 50.88806, 
    50.92697, 50.96566, 51.00413, 51.04239, 51.08043, 51.11825, 51.15585, 
    51.19323, 51.23039, 51.26733, 51.30405, 51.34055, 51.37682, 51.41287, 
    51.4487, 51.4843, 51.51968, 51.55482, 51.58975, 51.62444, 51.65891, 
    51.69315, 51.72715, 51.76093, 51.79448, 51.8278, 51.86088, 51.89373, 
    51.92635, 51.95874, 51.99089, 52.0228, 52.05449, 52.08593, 52.11713, 
    52.1481, 52.17884, 52.20933, 52.23958, 52.2696, 52.29937, 52.3289, 
    52.35819, 52.38724, 52.41605, 52.44461, 52.47293, 52.501, 52.52883, 
    52.55642, 52.58375, 52.61084, 52.63769, 52.66428, 52.69063, 52.71673, 
    52.74258, 52.76818, 52.79353, 52.81862, 52.84347, 52.86806, 52.8924, 
    52.91649, 52.94033, 52.96391, 52.98723, 53.0103, 53.03312, 53.05568, 
    53.07798, 53.10003, 53.12181, 53.14334, 53.16462, 53.18563, 53.20639, 
    53.22688, 53.24711, 53.26709, 53.2868, 53.30625, 53.32544, 53.34436, 
    53.36303, 53.38142, 53.39956, 53.41743, 53.43504, 53.45238, 53.46946, 
    53.48627, 53.50282, 53.5191, 53.53511, 53.55086, 53.56634, 53.58155, 
    53.59649, 53.61116, 53.62557, 53.63971, 53.65357, 53.66717, 53.6805, 
    53.69355, 53.70634, 53.71885, 53.7311, 53.74307, 53.75477, 53.7662, 
    53.77736, 53.78824, 53.79885, 53.80919, 53.81925, 53.82904, 53.83856, 
    53.8478, 53.85677, 53.86546, 53.87388, 53.88203, 53.88989, 53.89749, 
    53.90481, 53.91185, 53.91862, 53.92511, 53.93132, 53.93726, 53.94293, 
    53.94831, 53.95342, 53.95826, 53.96281, 53.96709, 53.9711, 53.97482, 
    53.97827, 53.98144, 53.98433, 53.98695, 53.98929, 53.99135, 53.99313, 
    53.99464, 53.99586, 53.99681, 53.99749, 53.99788, 53.998, 53.99784, 
    53.9974, 53.99669, 53.99569, 53.99442, 53.99287, 53.99104, 53.98894, 
    53.98655, 53.98389, 53.98096, 53.97774, 53.97425, 53.97048, 53.96643, 
    53.96211, 53.95751, 53.95263, 53.94748, 53.94205, 53.93634, 53.93036, 
    53.9241, 53.91756, 53.91076, 53.90367, 53.89631, 53.88867, 53.88076, 
    53.87257, 53.86411, 53.85537, 53.84636, 53.83707, 53.82751, 53.81768, 
    53.80757, 53.79719, 53.78653, 53.77561, 53.76441, 53.75294, 53.74119, 
    53.72918, 53.71689, 53.70433, 53.69151, 53.67841, 53.66504, 53.6514, 
    53.63749, 53.62331, 53.60886, 53.59414, 53.57916, 53.5639, 53.54839, 
    53.5326, 53.51654, 53.50022, 53.48363, 53.46678, 53.44966, 53.43227, 
    53.41462, 53.39671, 53.37853, 53.36009, 53.34138, 53.32242, 53.30319, 
    53.2837, 53.26394, 53.24393, 53.22366, 53.20312, 53.18232, 53.16127, 
    53.13996, 53.11839, 53.09656, 53.07447, 53.05213, 53.02953, 53.00667, 
    52.98356, 52.96019, 52.93657, 52.9127, 52.88857, 52.86419, 52.83955, 
    52.81467, 52.78953, 52.76414, 52.73851, 52.71262, 52.68648, 52.66009, 
    52.63346, 52.60658, 52.57944, 52.55207, 52.52444, 52.49658, 52.46846, 
    52.44011, 52.41151, 52.38266, 52.35357, 52.32425, 52.29467, 52.26486, 
    52.23481, 52.20452, 52.17399, 52.14322, 52.11221, 52.08097, 52.04949, 
    52.01777, 51.98582, 51.95363, 51.92121, 51.88855, 51.85566, 51.82254, 
    51.78919, 51.7556, 51.72179, 51.68774, 51.65347, 51.61897, 51.58424, 
    51.54928, 51.5141, 51.47868, 51.44305, 51.40719, 51.3711, 51.33479, 
    51.29826, 51.26151, 51.22453, 51.18734, 51.14992, 51.11228, 51.07442, 
    51.03635, 50.99806, 50.95955, 50.92083, 50.88189, 50.84273, 50.80336, 
    50.76378, 50.72398, 50.68398, 50.64376, 50.60332, 50.56268, 50.52183, 
    50.48077, 50.4395, 50.39803, 50.35635, 50.31446, 50.27236, 50.23006, 
    50.18756, 50.14485,
  45.47886, 45.53764, 45.59628, 45.65478, 45.71313, 45.77134, 45.82941, 
    45.88733, 45.9451, 46.00272, 46.0602, 46.11753, 46.17471, 46.23174, 
    46.28862, 46.34535, 46.40193, 46.45836, 46.51463, 46.57076, 46.62672, 
    46.68254, 46.73819, 46.7937, 46.84904, 46.90423, 46.95926, 47.01414, 
    47.06885, 47.12341, 47.1778, 47.23204, 47.28611, 47.34002, 47.39376, 
    47.44735, 47.50077, 47.55402, 47.60712, 47.66004, 47.7128, 47.76539, 
    47.81781, 47.87006, 47.92215, 47.97406, 48.0258, 48.07738, 48.12878, 
    48.18, 48.23106, 48.28194, 48.33265, 48.38317, 48.43353, 48.48371, 
    48.53371, 48.58353, 48.63318, 48.68264, 48.73193, 48.78103, 48.82996, 
    48.8787, 48.92725, 48.97563, 49.02382, 49.07183, 49.11965, 49.16728, 
    49.21473, 49.26199, 49.30906, 49.35595, 49.40264, 49.44914, 49.49546, 
    49.54158, 49.58751, 49.63324, 49.67879, 49.72414, 49.76929, 49.81425, 
    49.85901, 49.90357, 49.94794, 49.99211, 50.03608, 50.07985, 50.12342, 
    50.16679, 50.20995, 50.25291, 50.29568, 50.33823, 50.38058, 50.42273, 
    50.46468, 50.50641, 50.54794, 50.58926, 50.63037, 50.67127, 50.71196, 
    50.75244, 50.79271, 50.83277, 50.87262, 50.91225, 50.95167, 50.99087, 
    51.02986, 51.06863, 51.10719, 51.14552, 51.18364, 51.22155, 51.25923, 
    51.29669, 51.33393, 51.37095, 51.40775, 51.44432, 51.48067, 51.5168, 
    51.55271, 51.58839, 51.62384, 51.65907, 51.69406, 51.72883, 51.76337, 
    51.79769, 51.83177, 51.86562, 51.89925, 51.93264, 51.9658, 51.99872, 
    52.03141, 52.06387, 52.09609, 52.12808, 52.15983, 52.19135, 52.22263, 
    52.25366, 52.28447, 52.31503, 52.34535, 52.37543, 52.40527, 52.43487, 
    52.46423, 52.49335, 52.52222, 52.55085, 52.57923, 52.60737, 52.63527, 
    52.66291, 52.69031, 52.71747, 52.74437, 52.77103, 52.79744, 52.8236, 
    52.84951, 52.87517, 52.90058, 52.92573, 52.95064, 52.97529, 52.99969, 
    53.02383, 53.04773, 53.07136, 53.09475, 53.11787, 53.14074, 53.16335, 
    53.18571, 53.20781, 53.22965, 53.25123, 53.27256, 53.29362, 53.31442, 
    53.33496, 53.35525, 53.37527, 53.39503, 53.41453, 53.43376, 53.45274, 
    53.47144, 53.48989, 53.50807, 53.52599, 53.54364, 53.56102, 53.57814, 
    53.59499, 53.61158, 53.6279, 53.64395, 53.65974, 53.67525, 53.6905, 
    53.70548, 53.72019, 53.73463, 53.74881, 53.76271, 53.77634, 53.7897, 
    53.80279, 53.81561, 53.82815, 53.84042, 53.85243, 53.86415, 53.87561, 
    53.8868, 53.89771, 53.90834, 53.91871, 53.9288, 53.93861, 53.94815, 
    53.95742, 53.96641, 53.97512, 53.98357, 53.99173, 53.99962, 54.00723, 
    54.01457, 54.02163, 54.02842, 54.03492, 54.04116, 54.04711, 54.05279, 
    54.05819, 54.06331, 54.06816, 54.07272, 54.07701, 54.08103, 54.08476, 
    54.08822, 54.0914, 54.0943, 54.09692, 54.09927, 54.10133, 54.10312, 
    54.10463, 54.10586, 54.10681, 54.10749, 54.10788, 54.108, 54.10784, 
    54.1074, 54.10668, 54.10568, 54.10441, 54.10286, 54.10102, 54.09891, 
    54.09652, 54.09386, 54.09091, 54.08769, 54.08419, 54.08041, 54.07635, 
    54.07202, 54.06741, 54.06252, 54.05735, 54.05191, 54.04619, 54.04019, 
    54.03391, 54.02736, 54.02053, 54.01343, 54.00605, 53.99839, 53.99046, 
    53.98225, 53.97377, 53.96501, 53.95597, 53.94666, 53.93708, 53.92722, 
    53.91709, 53.90668, 53.896, 53.88505, 53.87382, 53.86232, 53.85055, 
    53.8385, 53.82618, 53.81359, 53.80074, 53.7876, 53.7742, 53.76052, 
    53.74658, 53.73237, 53.71788, 53.70313, 53.68811, 53.67282, 53.65726, 
    53.64143, 53.62534, 53.60897, 53.59235, 53.57545, 53.55829, 53.54086, 
    53.52317, 53.50521, 53.48699, 53.4685, 53.44975, 53.43074, 53.41146, 
    53.39192, 53.37212, 53.35206, 53.33173, 53.31115, 53.29031, 53.2692, 
    53.24784, 53.22621, 53.20433, 53.18219, 53.15979, 53.13714, 53.11423, 
    53.09106, 53.06764, 53.04396, 53.02003, 52.99585, 52.97141, 52.94672, 
    52.92177, 52.89658, 52.87113, 52.84543, 52.81948, 52.79328, 52.76683, 
    52.74013, 52.71319, 52.68599, 52.65855, 52.63087, 52.60294, 52.57476, 
    52.54633, 52.51767, 52.48876, 52.4596, 52.43021, 52.40057, 52.37069, 
    52.34057, 52.31021, 52.27961, 52.24877, 52.21769, 52.18638, 52.15482, 
    52.12304, 52.09101, 52.05875, 52.02626, 51.99353, 51.96057, 51.92737, 
    51.89394, 51.86029, 51.8264, 51.79227, 51.75793, 51.72335, 51.68854, 
    51.65351, 51.61824, 51.58276, 51.54704, 51.5111, 51.47494, 51.43855, 
    51.40194, 51.36511, 51.32805, 51.29078, 51.25328, 51.21556, 51.17763, 
    51.13947, 51.1011, 51.06251, 51.0237, 50.98468, 50.94545, 50.90599, 
    50.86633, 50.82645, 50.78636, 50.74606, 50.70554, 50.66481, 50.62388, 
    50.58273, 50.54138, 50.49982, 50.45805, 50.41608, 50.3739, 50.33152, 
    50.28893, 50.24613,
  45.5717, 45.63057, 45.6893, 45.74789, 45.80634, 45.86464, 45.92279, 
    45.9808, 46.03866, 46.09638, 46.15395, 46.21136, 46.26864, 46.32576, 
    46.38273, 46.43955, 46.49622, 46.55274, 46.60911, 46.66532, 46.72138, 
    46.77729, 46.83303, 46.88863, 46.94407, 46.99935, 47.05447, 47.10944, 
    47.16424, 47.21889, 47.27338, 47.3277, 47.38187, 47.43587, 47.48971, 
    47.54338, 47.59689, 47.65024, 47.70342, 47.75644, 47.80929, 47.86197, 
    47.91449, 47.96683, 48.019, 48.07101, 48.12285, 48.17451, 48.226, 
    48.27732, 48.32847, 48.37944, 48.43024, 48.48086, 48.5313, 48.58157, 
    48.63167, 48.68158, 48.73132, 48.78087, 48.83025, 48.87944, 48.92846, 
    48.97729, 49.02594, 49.0744, 49.12268, 49.17078, 49.21869, 49.26641, 
    49.31395, 49.3613, 49.40847, 49.45544, 49.50222, 49.54881, 49.59522, 
    49.64143, 49.68745, 49.73327, 49.7789, 49.82434, 49.86958, 49.91463, 
    49.95948, 50.00413, 50.04858, 50.09284, 50.1369, 50.18076, 50.22441, 
    50.26787, 50.31112, 50.35417, 50.39702, 50.43966, 50.4821, 50.52433, 
    50.56636, 50.60818, 50.64979, 50.6912, 50.73239, 50.77338, 50.81416, 
    50.85472, 50.89507, 50.93521, 50.97514, 51.01486, 51.05436, 51.09365, 
    51.13272, 51.17157, 51.21021, 51.24863, 51.28683, 51.32481, 51.36257, 
    51.40012, 51.43744, 51.47454, 51.51141, 51.54807, 51.5845, 51.6207, 
    51.65668, 51.69244, 51.72797, 51.76328, 51.79835, 51.8332, 51.86782, 
    51.90221, 51.93636, 51.97029, 52.00399, 52.03745, 52.07069, 52.10368, 
    52.13645, 52.16898, 52.20127, 52.23333, 52.26516, 52.29675, 52.32809, 
    52.3592, 52.39007, 52.4207, 52.4511, 52.48125, 52.51116, 52.54082, 
    52.57025, 52.59943, 52.62837, 52.65707, 52.68552, 52.71372, 52.74168, 
    52.76939, 52.79686, 52.82407, 52.85104, 52.87776, 52.90424, 52.93045, 
    52.95642, 52.98215, 53.00761, 53.03283, 53.05779, 53.0825, 53.10696, 
    53.13116, 53.15511, 53.17881, 53.20224, 53.22543, 53.24835, 53.27102, 
    53.29343, 53.31558, 53.33747, 53.35911, 53.38048, 53.4016, 53.42245, 
    53.44304, 53.46338, 53.48344, 53.50325, 53.5228, 53.54208, 53.5611, 
    53.57985, 53.59834, 53.61657, 53.63453, 53.65222, 53.66965, 53.68681, 
    53.70371, 53.72034, 53.73669, 53.75279, 53.76861, 53.78417, 53.79945, 
    53.81447, 53.82922, 53.84369, 53.8579, 53.87184, 53.8855, 53.8989, 
    53.91202, 53.92487, 53.93744, 53.94975, 53.96178, 53.97354, 53.98503, 
    53.99624, 54.00718, 54.01784, 54.02823, 54.03835, 54.04818, 54.05775, 
    54.06704, 54.07605, 54.08479, 54.09325, 54.10144, 54.10934, 54.11698, 
    54.12433, 54.13141, 54.13821, 54.14474, 54.15099, 54.15696, 54.16265, 
    54.16806, 54.1732, 54.17805, 54.18264, 54.18694, 54.19096, 54.1947, 
    54.19817, 54.20135, 54.20426, 54.20689, 54.20924, 54.21132, 54.21311, 
    54.21462, 54.21585, 54.21681, 54.21748, 54.21788, 54.218, 54.21784, 
    54.2174, 54.21667, 54.21568, 54.2144, 54.21284, 54.21101, 54.20889, 
    54.2065, 54.20382, 54.20087, 54.19764, 54.19413, 54.19034, 54.18628, 
    54.18193, 54.1773, 54.17241, 54.16722, 54.16177, 54.15603, 54.15002, 
    54.14373, 54.13716, 54.13031, 54.12319, 54.11579, 54.10811, 54.10016, 
    54.09193, 54.08342, 54.07464, 54.06559, 54.05626, 54.04665, 54.03676, 
    54.0266, 54.01617, 54.00546, 53.99448, 53.98323, 53.9717, 53.9599, 
    53.94782, 53.93547, 53.92285, 53.90996, 53.89679, 53.88336, 53.86965, 
    53.85567, 53.84142, 53.8269, 53.81211, 53.79705, 53.78172, 53.76612, 
    53.75026, 53.73413, 53.71772, 53.70105, 53.68412, 53.66691, 53.64944, 
    53.63171, 53.6137, 53.59544, 53.5769, 53.55811, 53.53905, 53.51973, 
    53.50014, 53.48029, 53.46018, 53.4398, 53.41917, 53.39827, 53.37712, 
    53.3557, 53.33403, 53.31209, 53.2899, 53.26745, 53.24474, 53.22178, 
    53.19855, 53.17508, 53.15134, 53.12735, 53.10311, 53.07861, 53.05386, 
    53.02886, 53.0036, 52.97809, 52.95234, 52.92632, 52.90006, 52.87355, 
    52.84679, 52.81979, 52.79253, 52.76503, 52.73727, 52.70927, 52.68103, 
    52.65254, 52.62381, 52.59483, 52.56561, 52.53615, 52.50644, 52.47649, 
    52.4463, 52.41587, 52.3852, 52.3543, 52.32315, 52.29176, 52.26014, 
    52.22828, 52.19618, 52.16385, 52.13128, 52.09848, 52.06544, 52.03218, 
    51.99867, 51.96494, 51.93098, 51.89678, 51.86235, 51.8277, 51.79282, 
    51.75771, 51.72237, 51.6868, 51.65101, 51.61499, 51.57875, 51.54229, 
    51.5056, 51.46868, 51.43155, 51.39419, 51.35661, 51.31882, 51.2808, 
    51.24257, 51.20411, 51.16544, 51.12655, 51.08744, 51.04813, 51.00859, 
    50.96884, 50.92888, 50.88871, 50.84832, 50.80772, 50.76691, 50.72589, 
    50.68466, 50.64322, 50.60158, 50.55973, 50.51767, 50.4754, 50.43293, 
    50.39025, 50.34737,
  45.66447, 45.72343, 45.78226, 45.84093, 45.89947, 45.95786, 46.01611, 
    46.07421, 46.13216, 46.18997, 46.24763, 46.30514, 46.3625, 46.41972, 
    46.47678, 46.5337, 46.59046, 46.64707, 46.70353, 46.75983, 46.81598, 
    46.87197, 46.92782, 46.98351, 47.03903, 47.09441, 47.14962, 47.20468, 
    47.25957, 47.31432, 47.36889, 47.42331, 47.47757, 47.53166, 47.58559, 
    47.63936, 47.69297, 47.7464, 47.79968, 47.85279, 47.90573, 47.9585, 
    48.01111, 48.06355, 48.11581, 48.16791, 48.21984, 48.27159, 48.32318, 
    48.37459, 48.42582, 48.47689, 48.52778, 48.57849, 48.62903, 48.67939, 
    48.72957, 48.77958, 48.8294, 48.87905, 48.92852, 48.97781, 49.02691, 
    49.07583, 49.12457, 49.17313, 49.2215, 49.26969, 49.31769, 49.3655, 
    49.41313, 49.46057, 49.50782, 49.55489, 49.60176, 49.64844, 49.69493, 
    49.74123, 49.78734, 49.83326, 49.87897, 49.9245, 49.96983, 50.01497, 
    50.05991, 50.10464, 50.14919, 50.19353, 50.23768, 50.28162, 50.32537, 
    50.36891, 50.41225, 50.45539, 50.49832, 50.54105, 50.58358, 50.62589, 
    50.66801, 50.70991, 50.75161, 50.7931, 50.83438, 50.87545, 50.91631, 
    50.95696, 50.9974, 51.03762, 51.07764, 51.11744, 51.15702, 51.19639, 
    51.23554, 51.27448, 51.3132, 51.3517, 51.38998, 51.42804, 51.46589, 
    51.50351, 51.54091, 51.57809, 51.61505, 51.65178, 51.68829, 51.72458, 
    51.76064, 51.79647, 51.83208, 51.86746, 51.90261, 51.93753, 51.97223, 
    52.00669, 52.04093, 52.07493, 52.1087, 52.14225, 52.17555, 52.20863, 
    52.24146, 52.27407, 52.30643, 52.33857, 52.37046, 52.40212, 52.43354, 
    52.46472, 52.49566, 52.52636, 52.55682, 52.58704, 52.61702, 52.64676, 
    52.67625, 52.7055, 52.7345, 52.76327, 52.79178, 52.82005, 52.84808, 
    52.87585, 52.90338, 52.93066, 52.9577, 52.98448, 53.01101, 53.0373, 
    53.06333, 53.08911, 53.11464, 53.13991, 53.16494, 53.1897, 53.21422, 
    53.23848, 53.26249, 53.28624, 53.30973, 53.33297, 53.35595, 53.37867, 
    53.40113, 53.42334, 53.44529, 53.46697, 53.4884, 53.50956, 53.53047, 
    53.55111, 53.5715, 53.59161, 53.61147, 53.63106, 53.65039, 53.66946, 
    53.68826, 53.70679, 53.72506, 53.74306, 53.7608, 53.77827, 53.79548, 
    53.81242, 53.82908, 53.84549, 53.86162, 53.87748, 53.89307, 53.9084, 
    53.92345, 53.93824, 53.95275, 53.96699, 53.98096, 53.99466, 54.00809, 
    54.02124, 54.03413, 54.04673, 54.05907, 54.07113, 54.08292, 54.09444, 
    54.10567, 54.11664, 54.12733, 54.13775, 54.14789, 54.15775, 54.16734, 
    54.17665, 54.18569, 54.19445, 54.20293, 54.21114, 54.21907, 54.22672, 
    54.2341, 54.24119, 54.24801, 54.25455, 54.26081, 54.2668, 54.27251, 
    54.27794, 54.28308, 54.28795, 54.29255, 54.29686, 54.30089, 54.30464, 
    54.30812, 54.31131, 54.31423, 54.31686, 54.31922, 54.3213, 54.32309, 
    54.32461, 54.32585, 54.32681, 54.32748, 54.32788, 54.328, 54.32784, 
    54.3274, 54.32667, 54.32567, 54.32439, 54.32283, 54.32099, 54.31887, 
    54.31647, 54.31379, 54.31083, 54.30759, 54.30407, 54.30027, 54.29619, 
    54.29184, 54.2872, 54.28229, 54.2771, 54.27162, 54.26587, 54.25984, 
    54.25354, 54.24695, 54.24009, 54.23295, 54.22553, 54.21783, 54.20986, 
    54.20161, 54.19308, 54.18428, 54.1752, 54.16584, 54.15621, 54.1463, 
    54.13612, 54.12566, 54.11493, 54.10392, 54.09263, 54.08107, 54.06924, 
    54.05714, 54.04476, 54.0321, 54.01918, 54.00598, 53.99251, 53.97877, 
    53.96476, 53.95047, 53.93592, 53.92109, 53.90599, 53.89062, 53.87499, 
    53.85908, 53.84291, 53.82647, 53.80975, 53.79277, 53.77553, 53.75801, 
    53.74023, 53.72219, 53.70388, 53.6853, 53.66646, 53.64735, 53.62798, 
    53.60835, 53.58845, 53.56829, 53.54786, 53.52718, 53.50623, 53.48503, 
    53.46356, 53.44183, 53.41984, 53.3976, 53.37509, 53.35233, 53.32931, 
    53.30603, 53.2825, 53.25871, 53.23466, 53.21036, 53.1858, 53.161, 
    53.13593, 53.11061, 53.08504, 53.05923, 53.03315, 53.00683, 52.98026, 
    52.95344, 52.92636, 52.89904, 52.87148, 52.84366, 52.8156, 52.78729, 
    52.75874, 52.72993, 52.70089, 52.6716, 52.64207, 52.6123, 52.58228, 
    52.55202, 52.52152, 52.49078, 52.4598, 52.42859, 52.39713, 52.36543, 
    52.3335, 52.30133, 52.26892, 52.23628, 52.20341, 52.1703, 52.13696, 
    52.10338, 52.06957, 52.03553, 52.00126, 51.96676, 51.93203, 51.89707, 
    51.86188, 51.82646, 51.79082, 51.75495, 51.71885, 51.68253, 51.64598, 
    51.60921, 51.57222, 51.53501, 51.49757, 51.45992, 51.42204, 51.38394, 
    51.34562, 51.30709, 51.26833, 51.22936, 51.19017, 51.15077, 51.11116, 
    51.07132, 51.03128, 50.99102, 50.95055, 50.90986, 50.86897, 50.82787, 
    50.78655, 50.74503, 50.7033, 50.66136, 50.61921, 50.57686, 50.53431, 
    50.49154, 50.44858,
  45.75718, 45.81623, 45.87515, 45.93392, 45.99255, 46.05103, 46.10936, 
    46.16756, 46.2256, 46.2835, 46.34125, 46.39885, 46.45631, 46.51361, 
    46.57077, 46.62778, 46.68463, 46.74133, 46.79788, 46.85428, 46.91052, 
    46.96661, 47.02254, 47.07832, 47.13394, 47.18941, 47.24471, 47.29986, 
    47.35485, 47.40968, 47.46436, 47.51886, 47.57321, 47.6274, 47.68142, 
    47.73528, 47.78898, 47.84251, 47.89588, 47.94908, 48.00211, 48.05498, 
    48.10767, 48.16021, 48.21257, 48.26476, 48.31677, 48.36862, 48.4203, 
    48.4718, 48.52313, 48.57429, 48.62527, 48.67607, 48.7267, 48.77715, 
    48.82743, 48.87753, 48.92744, 48.97718, 49.02674, 49.07612, 49.12531, 
    49.17433, 49.22316, 49.2718, 49.32027, 49.36855, 49.41664, 49.46454, 
    49.51226, 49.55979, 49.60714, 49.65429, 49.70125, 49.74802, 49.79461, 
    49.841, 49.88719, 49.9332, 49.97901, 50.02462, 50.07004, 50.11526, 
    50.16029, 50.20512, 50.24975, 50.29419, 50.33842, 50.38245, 50.42628, 
    50.46991, 50.51334, 50.55656, 50.59958, 50.6424, 50.68501, 50.72742, 
    50.76962, 50.81161, 50.85339, 50.89497, 50.93633, 50.97749, 51.01843, 
    51.05917, 51.09969, 51.14, 51.1801, 51.21998, 51.25964, 51.2991, 
    51.33833, 51.37735, 51.41615, 51.45473, 51.4931, 51.53125, 51.56917, 
    51.60687, 51.64436, 51.68161, 51.71865, 51.75547, 51.79206, 51.82842, 
    51.86456, 51.90047, 51.93616, 51.97161, 52.00684, 52.04185, 52.07662, 
    52.11116, 52.14547, 52.17955, 52.2134, 52.24701, 52.28039, 52.31354, 
    52.34645, 52.37913, 52.41157, 52.44378, 52.47574, 52.50747, 52.53896, 
    52.57021, 52.60123, 52.632, 52.66253, 52.69282, 52.72287, 52.75267, 
    52.78223, 52.81155, 52.84062, 52.86945, 52.89803, 52.92637, 52.95446, 
    52.9823, 53.00989, 53.03724, 53.06433, 53.09118, 53.11777, 53.14412, 
    53.17021, 53.19606, 53.22165, 53.24698, 53.27206, 53.29689, 53.32146, 
    53.34578, 53.36985, 53.39365, 53.4172, 53.4405, 53.46353, 53.48631, 
    53.50883, 53.53109, 53.55309, 53.57483, 53.5963, 53.61752, 53.63848, 
    53.65917, 53.6796, 53.69977, 53.71967, 53.73932, 53.75869, 53.7778, 
    53.79665, 53.81523, 53.83355, 53.85159, 53.86938, 53.88689, 53.90414, 
    53.92112, 53.93782, 53.95427, 53.97044, 53.98634, 54.00198, 54.01734, 
    54.03243, 54.04725, 54.0618, 54.07608, 54.09008, 54.10382, 54.11728, 
    54.13046, 54.14338, 54.15602, 54.16839, 54.18048, 54.1923, 54.20384, 
    54.21511, 54.2261, 54.23682, 54.24726, 54.25743, 54.26732, 54.27693, 
    54.28627, 54.29533, 54.30411, 54.31261, 54.32084, 54.32879, 54.33646, 
    54.34386, 54.35097, 54.35781, 54.36436, 54.37064, 54.37664, 54.38237, 
    54.38781, 54.39297, 54.39785, 54.40245, 54.40678, 54.41082, 54.41459, 
    54.41807, 54.42127, 54.42419, 54.42683, 54.4292, 54.43128, 54.43308, 
    54.4346, 54.43584, 54.4368, 54.43748, 54.43788, 54.438, 54.43784, 
    54.43739, 54.43667, 54.43567, 54.43438, 54.43282, 54.43097, 54.42884, 
    54.42644, 54.42375, 54.42078, 54.41753, 54.41401, 54.4102, 54.40611, 
    54.40174, 54.3971, 54.39217, 54.38696, 54.38148, 54.37571, 54.36967, 
    54.36335, 54.35674, 54.34986, 54.3427, 54.33527, 54.32755, 54.31956, 
    54.31129, 54.30274, 54.29391, 54.28481, 54.27543, 54.26577, 54.25584, 
    54.24563, 54.23515, 54.22438, 54.21334, 54.20203, 54.19044, 54.17859, 
    54.16645, 54.15404, 54.14135, 54.1284, 54.11517, 54.10166, 54.08789, 
    54.07384, 54.05952, 54.04492, 54.03006, 54.01493, 53.99952, 53.98384, 
    53.9679, 53.95168, 53.9352, 53.91845, 53.90143, 53.88414, 53.86658, 
    53.84876, 53.83067, 53.81231, 53.79369, 53.7748, 53.75564, 53.73623, 
    53.71654, 53.6966, 53.67639, 53.65591, 53.63518, 53.61418, 53.59292, 
    53.5714, 53.54962, 53.52758, 53.50528, 53.48272, 53.4599, 53.43683, 
    53.41349, 53.3899, 53.36606, 53.34195, 53.3176, 53.29298, 53.26811, 
    53.24299, 53.21761, 53.19198, 53.1661, 53.13997, 53.11358, 53.08695, 
    53.06006, 53.03293, 53.00554, 52.97791, 52.95003, 52.9219, 52.89353, 
    52.86491, 52.83604, 52.80693, 52.77757, 52.74797, 52.71813, 52.68804, 
    52.65771, 52.62714, 52.59634, 52.56528, 52.534, 52.50247, 52.4707, 
    52.43869, 52.40645, 52.37397, 52.34126, 52.30831, 52.27513, 52.24171, 
    52.20806, 52.17418, 52.14006, 52.10571, 52.07113, 52.03632, 52.00129, 
    51.96602, 51.93053, 51.89481, 51.85886, 51.82268, 51.78628, 51.74966, 
    51.71281, 51.67574, 51.63844, 51.60093, 51.56319, 51.52523, 51.48705, 
    51.44865, 51.41003, 51.37119, 51.33214, 51.29287, 51.25338, 51.21368, 
    51.17377, 51.13364, 51.0933, 51.05274, 51.01197, 50.97099, 50.9298, 
    50.8884, 50.84679, 50.80498, 50.76295, 50.72072, 50.67828, 50.63564, 
    50.59279, 50.54974,
  45.84983, 45.90897, 45.96798, 46.02684, 46.08556, 46.14413, 46.20256, 
    46.26084, 46.31898, 46.37697, 46.43481, 46.49251, 46.55005, 46.60745, 
    46.6647, 46.72179, 46.77874, 46.83554, 46.89218, 46.94867, 47.005, 
    47.06118, 47.11721, 47.17308, 47.22879, 47.28435, 47.33975, 47.39499, 
    47.45007, 47.505, 47.55976, 47.61436, 47.6688, 47.72308, 47.7772, 
    47.83115, 47.88494, 47.93856, 47.99202, 48.04531, 48.09844, 48.1514, 
    48.20419, 48.25681, 48.30927, 48.36155, 48.41366, 48.4656, 48.51736, 
    48.56896, 48.62038, 48.67163, 48.72271, 48.7736, 48.82432, 48.87487, 
    48.92524, 48.97542, 49.02543, 49.07526, 49.12491, 49.17438, 49.22367, 
    49.27277, 49.3217, 49.37043, 49.41899, 49.46736, 49.51554, 49.56354, 
    49.61135, 49.65897, 49.7064, 49.75364, 49.8007, 49.84756, 49.89423, 
    49.94071, 49.987, 50.03309, 50.07899, 50.1247, 50.17021, 50.21552, 
    50.26064, 50.30555, 50.35027, 50.39479, 50.43911, 50.48323, 50.52715, 
    50.57087, 50.61439, 50.6577, 50.70081, 50.74371, 50.78641, 50.8289, 
    50.87119, 50.91327, 50.95514, 50.9968, 51.03825, 51.07949, 51.12052, 
    51.16134, 51.20195, 51.24234, 51.28252, 51.32249, 51.36224, 51.40177, 
    51.44109, 51.48019, 51.51908, 51.55774, 51.59619, 51.63441, 51.67242, 
    51.71021, 51.74777, 51.78511, 51.82223, 51.85912, 51.89579, 51.93223, 
    51.96845, 52.00444, 52.04021, 52.07574, 52.11105, 52.14613, 52.18098, 
    52.2156, 52.24998, 52.28414, 52.31806, 52.35175, 52.38521, 52.41843, 
    52.45142, 52.48417, 52.51668, 52.54896, 52.581, 52.6128, 52.64436, 
    52.67569, 52.70677, 52.73761, 52.76821, 52.79857, 52.82869, 52.85856, 
    52.88819, 52.91758, 52.94672, 52.97561, 53.00426, 53.03266, 53.06082, 
    53.08873, 53.11638, 53.14379, 53.17095, 53.19786, 53.22452, 53.25093, 
    53.27708, 53.30299, 53.32864, 53.35403, 53.37917, 53.40406, 53.4287, 
    53.45307, 53.47719, 53.50106, 53.52467, 53.54801, 53.5711, 53.59394, 
    53.61651, 53.63882, 53.66087, 53.68267, 53.7042, 53.72547, 53.74648, 
    53.76722, 53.7877, 53.80791, 53.82787, 53.84756, 53.86698, 53.88614, 
    53.90504, 53.92366, 53.94202, 53.96011, 53.97794, 53.9955, 54.01279, 
    54.02981, 54.04656, 54.06304, 54.07925, 54.0952, 54.11087, 54.12627, 
    54.1414, 54.15626, 54.17085, 54.18516, 54.1992, 54.21297, 54.22646, 
    54.23968, 54.25263, 54.2653, 54.2777, 54.28982, 54.30167, 54.31324, 
    54.32454, 54.33556, 54.34631, 54.35678, 54.36697, 54.37688, 54.38652, 
    54.39588, 54.40496, 54.41377, 54.42229, 54.43054, 54.43851, 54.4462, 
    54.45361, 54.46075, 54.4676, 54.47417, 54.48047, 54.48648, 54.49222, 
    54.49768, 54.50285, 54.50775, 54.51236, 54.5167, 54.52075, 54.52452, 
    54.52802, 54.53123, 54.53416, 54.53681, 54.53918, 54.54126, 54.54307, 
    54.54459, 54.54584, 54.5468, 54.54748, 54.54788, 54.548, 54.54784, 
    54.54739, 54.54667, 54.54566, 54.54437, 54.5428, 54.54095, 54.53882, 
    54.53641, 54.53371, 54.53074, 54.52748, 54.52394, 54.52013, 54.51603, 
    54.51165, 54.50699, 54.50205, 54.49683, 54.49133, 54.48555, 54.47949, 
    54.47316, 54.46654, 54.45964, 54.45246, 54.445, 54.43727, 54.42926, 
    54.42096, 54.41239, 54.40355, 54.39442, 54.38501, 54.37533, 54.36538, 
    54.35514, 54.34463, 54.33384, 54.32277, 54.31143, 54.29982, 54.28793, 
    54.27576, 54.26332, 54.2506, 54.23761, 54.22435, 54.21081, 54.19699, 
    54.18291, 54.16856, 54.15393, 54.13903, 54.12385, 54.10841, 54.09269, 
    54.07671, 54.06046, 54.04393, 54.02713, 54.01007, 53.99274, 53.97514, 
    53.95727, 53.93914, 53.92073, 53.90207, 53.88313, 53.86393, 53.84446, 
    53.82473, 53.80474, 53.78448, 53.76395, 53.74317, 53.72212, 53.70081, 
    53.67924, 53.6574, 53.63531, 53.61296, 53.59034, 53.56747, 53.54434, 
    53.52095, 53.4973, 53.4734, 53.44923, 53.42482, 53.40014, 53.37521, 
    53.35003, 53.3246, 53.2989, 53.27296, 53.24677, 53.22032, 53.19362, 
    53.16667, 53.13947, 53.11203, 53.08433, 53.05638, 53.02819, 52.99974, 
    52.97106, 52.94212, 52.91294, 52.88352, 52.85385, 52.82394, 52.79379, 
    52.76339, 52.73275, 52.70187, 52.67075, 52.63939, 52.60778, 52.57595, 
    52.54387, 52.51155, 52.479, 52.44621, 52.41319, 52.37993, 52.34644, 
    52.31271, 52.27875, 52.24456, 52.21014, 52.17548, 52.14059, 52.10548, 
    52.07014, 52.03456, 51.99876, 51.96274, 51.92648, 51.89, 51.8533, 
    51.81637, 51.77922, 51.74184, 51.70424, 51.66642, 51.62838, 51.59012, 
    51.55164, 51.51294, 51.47402, 51.43489, 51.39553, 51.35596, 51.31618, 
    51.27618, 51.23597, 51.19554, 51.1549, 51.11404, 51.07298, 51.0317, 
    50.99022, 50.94852, 50.90662, 50.86451, 50.82219, 50.77967, 50.73694, 
    50.694, 50.65086,
  45.94241, 46.00165, 46.06075, 46.1197, 46.17851, 46.23717, 46.29569, 
    46.35407, 46.4123, 46.47038, 46.52831, 46.5861, 46.64374, 46.70123, 
    46.75857, 46.81576, 46.8728, 46.92968, 46.98642, 47.043, 47.09942, 
    47.1557, 47.21181, 47.26778, 47.32359, 47.37923, 47.43473, 47.49006, 
    47.54523, 47.60025, 47.65511, 47.7098, 47.76434, 47.81871, 47.87292, 
    47.92696, 47.98084, 48.03456, 48.08811, 48.1415, 48.19472, 48.24777, 
    48.30065, 48.35336, 48.40591, 48.45829, 48.51049, 48.56252, 48.61438, 
    48.66607, 48.71758, 48.76892, 48.82009, 48.87108, 48.92189, 48.97253, 
    49.02299, 49.07327, 49.12337, 49.17329, 49.22304, 49.2726, 49.32198, 
    49.37117, 49.42019, 49.46902, 49.51766, 49.56612, 49.6144, 49.66248, 
    49.71038, 49.7581, 49.80562, 49.85295, 49.9001, 49.94705, 49.99382, 
    50.04039, 50.08676, 50.13295, 50.17894, 50.22473, 50.27033, 50.31573, 
    50.36094, 50.40594, 50.45075, 50.49536, 50.53977, 50.58398, 50.62799, 
    50.67179, 50.7154, 50.7588, 50.80199, 50.84498, 50.88777, 50.93035, 
    50.97272, 51.01488, 51.05684, 51.09859, 51.14013, 51.18145, 51.22257, 
    51.26347, 51.30416, 51.34464, 51.38491, 51.42496, 51.46479, 51.50441, 
    51.54382, 51.583, 51.62197, 51.66072, 51.69925, 51.73755, 51.77564, 
    51.81351, 51.85115, 51.88857, 51.92577, 51.96275, 51.99949, 52.03602, 
    52.07232, 52.10839, 52.14423, 52.17984, 52.21523, 52.25039, 52.28531, 
    52.32001, 52.35447, 52.3887, 52.4227, 52.45647, 52.49, 52.52329, 
    52.55635, 52.58918, 52.62177, 52.65412, 52.68623, 52.71811, 52.74974, 
    52.78114, 52.81229, 52.8432, 52.87387, 52.9043, 52.93449, 52.96443, 
    52.99413, 53.02359, 53.0528, 53.08176, 53.11047, 53.13894, 53.16716, 
    53.19513, 53.22286, 53.25033, 53.27755, 53.30453, 53.33125, 53.35772, 
    53.38394, 53.4099, 53.43561, 53.46107, 53.48627, 53.51122, 53.53591, 
    53.56035, 53.58453, 53.60845, 53.63211, 53.65552, 53.67867, 53.70155, 
    53.72418, 53.74655, 53.76865, 53.7905, 53.81208, 53.8334, 53.85446, 
    53.87526, 53.89579, 53.91605, 53.93606, 53.9558, 53.97527, 53.99447, 
    54.01341, 54.03209, 54.05049, 54.06863, 54.0865, 54.1041, 54.12143, 
    54.1385, 54.15529, 54.17181, 54.18806, 54.20405, 54.21976, 54.2352, 
    54.25037, 54.26526, 54.27988, 54.29424, 54.30831, 54.32211, 54.33564, 
    54.3489, 54.36187, 54.37458, 54.38701, 54.39916, 54.41104, 54.42265, 
    54.43397, 54.44502, 54.45579, 54.46629, 54.47651, 54.48644, 54.49611, 
    54.50549, 54.5146, 54.52342, 54.53197, 54.54024, 54.54823, 54.55594, 
    54.56337, 54.57052, 54.5774, 54.58399, 54.5903, 54.59633, 54.60208, 
    54.60755, 54.61274, 54.61765, 54.62227, 54.62662, 54.63068, 54.63446, 
    54.63797, 54.64119, 54.64412, 54.64678, 54.64915, 54.65125, 54.65306, 
    54.65459, 54.65583, 54.6568, 54.65748, 54.65788, 54.658, 54.65784, 
    54.65739, 54.65666, 54.65565, 54.65436, 54.65279, 54.65093, 54.6488, 
    54.64638, 54.64368, 54.64069, 54.63743, 54.63388, 54.63005, 54.62595, 
    54.62156, 54.61689, 54.61193, 54.6067, 54.60119, 54.59539, 54.58932, 
    54.58296, 54.57633, 54.56941, 54.56221, 54.55474, 54.54699, 54.53895, 
    54.53064, 54.52205, 54.51317, 54.50402, 54.49459, 54.48489, 54.47491, 
    54.46465, 54.45411, 54.44329, 54.4322, 54.42083, 54.40918, 54.39726, 
    54.38506, 54.37259, 54.35984, 54.34682, 54.33352, 54.31995, 54.3061, 
    54.29198, 54.27759, 54.26292, 54.24799, 54.23278, 54.21729, 54.20154, 
    54.18551, 54.16922, 54.15265, 54.13581, 54.11871, 54.10133, 54.08369, 
    54.06578, 54.0476, 54.02915, 54.01043, 53.99145, 53.9722, 53.95269, 
    53.93291, 53.91286, 53.89256, 53.87198, 53.85115, 53.83005, 53.80869, 
    53.78706, 53.76517, 53.74303, 53.72062, 53.69795, 53.67502, 53.65183, 
    53.62838, 53.60468, 53.58072, 53.5565, 53.53202, 53.50729, 53.4823, 
    53.45706, 53.43156, 53.40581, 53.37981, 53.35355, 53.32704, 53.30028, 
    53.27327, 53.246, 53.21849, 53.19072, 53.16271, 53.13445, 53.10595, 
    53.07719, 53.04819, 53.01894, 52.98945, 52.95971, 52.92973, 52.89951, 
    52.86904, 52.83833, 52.80738, 52.77618, 52.74475, 52.71308, 52.68117, 
    52.64902, 52.61663, 52.584, 52.55114, 52.51804, 52.48471, 52.45114, 
    52.41734, 52.3833, 52.34903, 52.31453, 52.2798, 52.24484, 52.20965, 
    52.17422, 52.13857, 52.1027, 52.06659, 52.03025, 51.9937, 51.95691, 
    51.9199, 51.88267, 51.84521, 51.80753, 51.76963, 51.73151, 51.69316, 
    51.6546, 51.61582, 51.57682, 51.5376, 51.49816, 51.45851, 51.41864, 
    51.37856, 51.33826, 51.29774, 51.25702, 51.21608, 51.17493, 51.13357, 
    51.092, 51.05022, 51.00823, 50.96603, 50.92363, 50.88102, 50.8382, 
    50.79517, 50.75195,
  46.03493, 46.09426, 46.15345, 46.21249, 46.2714, 46.33015, 46.38876, 
    46.44723, 46.50555, 46.56372, 46.62175, 46.67963, 46.73736, 46.79494, 
    46.85238, 46.90966, 46.96679, 47.02377, 47.08059, 47.13726, 47.19378, 
    47.25015, 47.30636, 47.36242, 47.41832, 47.47406, 47.52964, 47.58507, 
    47.64034, 47.69545, 47.7504, 47.80518, 47.85981, 47.91428, 47.96858, 
    48.02272, 48.07669, 48.1305, 48.18415, 48.23763, 48.29094, 48.34408, 
    48.39706, 48.44986, 48.5025, 48.55497, 48.60727, 48.65939, 48.71135, 
    48.76313, 48.81473, 48.86617, 48.91742, 48.96851, 49.01941, 49.07014, 
    49.12069, 49.17107, 49.22126, 49.27127, 49.32111, 49.37076, 49.42023, 
    49.46952, 49.51863, 49.56755, 49.61629, 49.66484, 49.7132, 49.76138, 
    49.80938, 49.85718, 49.90479, 49.95222, 49.99945, 50.0465, 50.09335, 
    50.14001, 50.18648, 50.23275, 50.27884, 50.32472, 50.37041, 50.4159, 
    50.46119, 50.50629, 50.55119, 50.59589, 50.64038, 50.68468, 50.72878, 
    50.77267, 50.81636, 50.85985, 50.90314, 50.94622, 50.98909, 51.03175, 
    51.07421, 51.11647, 51.15851, 51.20034, 51.24197, 51.28338, 51.32458, 
    51.36557, 51.40635, 51.44691, 51.48726, 51.5274, 51.56732, 51.60702, 
    51.6465, 51.68578, 51.72482, 51.76366, 51.80227, 51.84066, 51.87883, 
    51.91678, 51.9545, 51.992, 52.02929, 52.06634, 52.10317, 52.13977, 
    52.17615, 52.2123, 52.24822, 52.28392, 52.31938, 52.35461, 52.38962, 
    52.42439, 52.45893, 52.49324, 52.52731, 52.56115, 52.59476, 52.62813, 
    52.66127, 52.69417, 52.72683, 52.75925, 52.79144, 52.82339, 52.85509, 
    52.88656, 52.91779, 52.94877, 52.97952, 53.01002, 53.04027, 53.07029, 
    53.10005, 53.12957, 53.15885, 53.18788, 53.21666, 53.2452, 53.27349, 
    53.30153, 53.32931, 53.35685, 53.38414, 53.41117, 53.43796, 53.4645, 
    53.49078, 53.5168, 53.54258, 53.56809, 53.59336, 53.61836, 53.64311, 
    53.66761, 53.69184, 53.71582, 53.73954, 53.76301, 53.78621, 53.80915, 
    53.83184, 53.85426, 53.87642, 53.89832, 53.91995, 53.94133, 53.96244, 
    53.98328, 54.00386, 54.02418, 54.04424, 54.06402, 54.08354, 54.10279, 
    54.12178, 54.1405, 54.15895, 54.17714, 54.19505, 54.2127, 54.23007, 
    54.24718, 54.26401, 54.28057, 54.29687, 54.31289, 54.32864, 54.34412, 
    54.35933, 54.37426, 54.38892, 54.40331, 54.41742, 54.43126, 54.44482, 
    54.4581, 54.47112, 54.48386, 54.49632, 54.5085, 54.52041, 54.53204, 
    54.5434, 54.55447, 54.56527, 54.57579, 54.58604, 54.596, 54.60569, 
    54.6151, 54.62423, 54.63308, 54.64165, 54.64994, 54.65795, 54.66568, 
    54.67313, 54.6803, 54.68719, 54.69379, 54.70012, 54.70617, 54.71193, 
    54.71742, 54.72262, 54.72754, 54.73218, 54.73653, 54.74061, 54.7444, 
    54.74791, 54.75114, 54.75409, 54.75675, 54.75913, 54.76123, 54.76304, 
    54.76458, 54.76583, 54.76679, 54.76748, 54.76788, 54.768, 54.76783, 
    54.76739, 54.76666, 54.76565, 54.76435, 54.76278, 54.76091, 54.75877, 
    54.75635, 54.75364, 54.75065, 54.74738, 54.74382, 54.73998, 54.73587, 
    54.73146, 54.72678, 54.72182, 54.71657, 54.71104, 54.70523, 54.69914, 
    54.69277, 54.68612, 54.67918, 54.67197, 54.66447, 54.6567, 54.64864, 
    54.64031, 54.63169, 54.6228, 54.61363, 54.60418, 54.59444, 54.58443, 
    54.57415, 54.56358, 54.55274, 54.54162, 54.53022, 54.51854, 54.50659, 
    54.49436, 54.48186, 54.46908, 54.45602, 54.44269, 54.42908, 54.4152, 
    54.40105, 54.38662, 54.37192, 54.35694, 54.34169, 54.32617, 54.31038, 
    54.29431, 54.27797, 54.26137, 54.24449, 54.22734, 54.20992, 54.19223, 
    54.17427, 54.15605, 54.13756, 54.11879, 54.09977, 54.08047, 54.06091, 
    54.04108, 54.02098, 54.00063, 53.98, 53.95911, 53.93796, 53.91655, 
    53.89487, 53.87293, 53.85073, 53.82827, 53.80554, 53.78256, 53.75932, 
    53.73581, 53.71205, 53.68803, 53.66375, 53.63922, 53.61443, 53.58937, 
    53.56407, 53.53851, 53.5127, 53.48663, 53.46032, 53.43374, 53.40692, 
    53.37984, 53.35251, 53.32493, 53.2971, 53.26903, 53.2407, 53.21213, 
    53.1833, 53.15424, 53.12492, 53.09536, 53.06555, 53.0355, 53.00521, 
    52.97467, 52.94389, 52.91286, 52.8816, 52.8501, 52.81835, 52.78637, 
    52.75414, 52.72168, 52.68898, 52.65604, 52.62287, 52.58946, 52.55582, 
    52.52194, 52.48783, 52.45348, 52.4189, 52.38409, 52.34906, 52.31379, 
    52.27828, 52.24255, 52.2066, 52.17041, 52.134, 52.09736, 52.06049, 
    52.0234, 51.98609, 51.94855, 51.91079, 51.87281, 51.8346, 51.79617, 
    51.75753, 51.71866, 51.67958, 51.64027, 51.60075, 51.56102, 51.52106, 
    51.48089, 51.44051, 51.39991, 51.3591, 51.31808, 51.27684, 51.2354, 
    51.19374, 51.15187, 51.10979, 51.06751, 51.02502, 50.98232, 50.93941, 
    50.89631, 50.85299,
  46.12739, 46.18681, 46.24609, 46.30523, 46.36422, 46.42307, 46.48177, 
    46.54033, 46.59874, 46.65701, 46.71513, 46.7731, 46.83092, 46.8886, 
    46.94612, 47.00349, 47.06071, 47.11779, 47.17471, 47.23147, 47.28809, 
    47.34454, 47.40085, 47.457, 47.51299, 47.56882, 47.6245, 47.68002, 
    47.73539, 47.79058, 47.84563, 47.90051, 47.95523, 48.00979, 48.06418, 
    48.11842, 48.17248, 48.22638, 48.28012, 48.33369, 48.3871, 48.44033, 
    48.4934, 48.54631, 48.59904, 48.6516, 48.70399, 48.75621, 48.80825, 
    48.86013, 48.91183, 48.96335, 49.01471, 49.06588, 49.11688, 49.1677, 
    49.21835, 49.26881, 49.3191, 49.36921, 49.41913, 49.46888, 49.51844, 
    49.56782, 49.61702, 49.66603, 49.71486, 49.76351, 49.81197, 49.86024, 
    49.90832, 49.95621, 50.00392, 50.05144, 50.09876, 50.1459, 50.19284, 
    50.23959, 50.28615, 50.33252, 50.37869, 50.42466, 50.47044, 50.51602, 
    50.56141, 50.60659, 50.65158, 50.69637, 50.74096, 50.78534, 50.82953, 
    50.87351, 50.91729, 50.96087, 51.00424, 51.04741, 51.09037, 51.13312, 
    51.17567, 51.21801, 51.26014, 51.30206, 51.34377, 51.38527, 51.42656, 
    51.46763, 51.5085, 51.54914, 51.58958, 51.6298, 51.6698, 51.70959, 
    51.74916, 51.78851, 51.82765, 51.86656, 51.90526, 51.94373, 51.98198, 
    52.02002, 52.05782, 52.09541, 52.13277, 52.1699, 52.20681, 52.2435, 
    52.27995, 52.31618, 52.35218, 52.38796, 52.4235, 52.45881, 52.4939, 
    52.52875, 52.56336, 52.59775, 52.6319, 52.66582, 52.6995, 52.73295, 
    52.76616, 52.79913, 52.83187, 52.86437, 52.89663, 52.92865, 52.96043, 
    52.99197, 53.02327, 53.05432, 53.08514, 53.1157, 53.14603, 53.17611, 
    53.20595, 53.23554, 53.26489, 53.29398, 53.32283, 53.35144, 53.37979, 
    53.4079, 53.43575, 53.46336, 53.49071, 53.51781, 53.54466, 53.57125, 
    53.5976, 53.62368, 53.64952, 53.6751, 53.70042, 53.72549, 53.7503, 
    53.77486, 53.79915, 53.82319, 53.84697, 53.87049, 53.89375, 53.91674, 
    53.93948, 53.96196, 53.98417, 54.00613, 54.02781, 54.04924, 54.0704, 
    54.0913, 54.11193, 54.1323, 54.1524, 54.17224, 54.19181, 54.21111, 
    54.23014, 54.24891, 54.2674, 54.28563, 54.30359, 54.32128, 54.3387, 
    54.35585, 54.37273, 54.38933, 54.40567, 54.42173, 54.43752, 54.45304, 
    54.46828, 54.48325, 54.49795, 54.51237, 54.52652, 54.54039, 54.55399, 
    54.56731, 54.58036, 54.59312, 54.60562, 54.61783, 54.62977, 54.64143, 
    54.65282, 54.66392, 54.67475, 54.6853, 54.69557, 54.70556, 54.71527, 
    54.7247, 54.73386, 54.74273, 54.75132, 54.75963, 54.76766, 54.77541, 
    54.78288, 54.79007, 54.79698, 54.8036, 54.80995, 54.81601, 54.82179, 
    54.82729, 54.8325, 54.83744, 54.84209, 54.84645, 54.85054, 54.85434, 
    54.85786, 54.8611, 54.86405, 54.86672, 54.86911, 54.87121, 54.87303, 
    54.87457, 54.87582, 54.87679, 54.87748, 54.87788, 54.878, 54.87783, 
    54.87739, 54.87666, 54.87564, 54.87434, 54.87276, 54.8709, 54.86875, 
    54.86632, 54.8636, 54.8606, 54.85732, 54.85376, 54.84991, 54.84578, 
    54.84137, 54.83667, 54.8317, 54.82644, 54.82089, 54.81507, 54.80896, 
    54.80257, 54.79591, 54.78895, 54.78172, 54.77421, 54.76641, 54.75834, 
    54.74998, 54.74134, 54.73243, 54.72323, 54.71375, 54.704, 54.69396, 
    54.68365, 54.67306, 54.66219, 54.65104, 54.63961, 54.6279, 54.61592, 
    54.60366, 54.59113, 54.57831, 54.56522, 54.55186, 54.53822, 54.5243, 
    54.51011, 54.49564, 54.4809, 54.46589, 54.4506, 54.43504, 54.41921, 
    54.4031, 54.38673, 54.37008, 54.35315, 54.33596, 54.3185, 54.30077, 
    54.28277, 54.2645, 54.24596, 54.22715, 54.20807, 54.18873, 54.16912, 
    54.14924, 54.1291, 54.10868, 54.08801, 54.06707, 54.04587, 54.0244, 
    54.00267, 53.98068, 53.95842, 53.9359, 53.91312, 53.89008, 53.86678, 
    53.84322, 53.8194, 53.79533, 53.77099, 53.7464, 53.72154, 53.69643, 
    53.67107, 53.64545, 53.61958, 53.59344, 53.56706, 53.54043, 53.51354, 
    53.4864, 53.459, 53.43136, 53.40347, 53.37532, 53.34693, 53.31829, 
    53.2894, 53.26026, 53.23088, 53.20125, 53.17137, 53.14125, 53.11089, 
    53.08028, 53.04942, 53.01833, 52.987, 52.95542, 52.9236, 52.89154, 
    52.85924, 52.82671, 52.79393, 52.76092, 52.72767, 52.69419, 52.66047, 
    52.62651, 52.59233, 52.5579, 52.52325, 52.48836, 52.45324, 52.41789, 
    52.38231, 52.3465, 52.31047, 52.2742, 52.23771, 52.20099, 52.16404, 
    52.12687, 52.08948, 52.05186, 52.01401, 51.97595, 51.93766, 51.89915, 
    51.86042, 51.82147, 51.7823, 51.74292, 51.70331, 51.66349, 51.62345, 
    51.5832, 51.54273, 51.50204, 51.46115, 51.42004, 51.37872, 51.33718, 
    51.29544, 51.25349, 51.21133, 51.16895, 51.12637, 51.08359, 51.04059, 
    50.99739, 50.95399,
  46.21978, 46.2793, 46.33867, 46.39789, 46.45698, 46.51592, 46.57471, 
    46.63337, 46.69187, 46.75023, 46.80844, 46.8665, 46.92442, 46.98219, 
    47.0398, 47.09727, 47.15459, 47.21175, 47.26876, 47.32562, 47.38233, 
    47.43888, 47.49528, 47.55152, 47.6076, 47.66353, 47.7193, 47.77492, 
    47.83037, 47.88567, 47.9408, 47.99578, 48.05059, 48.10524, 48.15973, 
    48.21405, 48.26822, 48.32221, 48.37604, 48.42971, 48.48321, 48.53654, 
    48.5897, 48.64269, 48.69552, 48.74817, 48.80066, 48.85297, 48.90511, 
    48.95707, 49.00887, 49.06049, 49.11193, 49.1632, 49.21429, 49.26521, 
    49.31594, 49.3665, 49.41689, 49.46708, 49.5171, 49.56694, 49.6166, 
    49.66607, 49.71536, 49.76447, 49.81339, 49.86213, 49.91068, 49.95904, 
    50.00721, 50.0552, 50.103, 50.15061, 50.19802, 50.24525, 50.29229, 
    50.33913, 50.38578, 50.43224, 50.4785, 50.52456, 50.57043, 50.6161, 
    50.66158, 50.70686, 50.75193, 50.79681, 50.84149, 50.88596, 50.93024, 
    50.97431, 51.01818, 51.06184, 51.1053, 51.14856, 51.19161, 51.23445, 
    51.27708, 51.31951, 51.36173, 51.40374, 51.44553, 51.48712, 51.5285, 
    51.56966, 51.61061, 51.65134, 51.69186, 51.73217, 51.77225, 51.81213, 
    51.85178, 51.89122, 51.93044, 51.96944, 52.00821, 52.04677, 52.08511, 
    52.12322, 52.16111, 52.19878, 52.23622, 52.27343, 52.31042, 52.34719, 
    52.38373, 52.42004, 52.45612, 52.49197, 52.52759, 52.56298, 52.59814, 
    52.63307, 52.66777, 52.70223, 52.73646, 52.77045, 52.80421, 52.83774, 
    52.87102, 52.90407, 52.93688, 52.96946, 53.00179, 53.03388, 53.06573, 
    53.09735, 53.12872, 53.15985, 53.19073, 53.22137, 53.25177, 53.28192, 
    53.31183, 53.34149, 53.3709, 53.40007, 53.42899, 53.45766, 53.48608, 
    53.51425, 53.54217, 53.56984, 53.59726, 53.62442, 53.65134, 53.678, 
    53.7044, 53.73055, 53.75645, 53.78209, 53.80748, 53.8326, 53.85748, 
    53.88209, 53.90644, 53.93054, 53.95437, 53.97795, 54.00127, 54.02432, 
    54.04712, 54.06965, 54.09192, 54.11392, 54.13567, 54.15714, 54.17836, 
    54.19931, 54.21999, 54.24041, 54.26056, 54.28045, 54.30006, 54.31941, 
    54.33849, 54.3573, 54.37585, 54.39412, 54.41212, 54.42986, 54.44732, 
    54.46452, 54.48143, 54.49809, 54.51446, 54.53056, 54.54639, 54.56195, 
    54.57723, 54.59224, 54.60697, 54.62143, 54.63562, 54.64952, 54.66315, 
    54.67651, 54.68959, 54.70239, 54.71492, 54.72717, 54.73913, 54.75082, 
    54.76224, 54.77337, 54.78423, 54.7948, 54.8051, 54.81511, 54.82485, 
    54.83431, 54.84348, 54.85238, 54.86099, 54.86933, 54.87738, 54.88515, 
    54.89264, 54.89985, 54.90677, 54.91341, 54.91977, 54.92585, 54.93164, 
    54.93716, 54.94238, 54.94733, 54.95199, 54.95637, 54.96047, 54.96428, 
    54.96781, 54.97105, 54.97401, 54.97669, 54.97908, 54.98119, 54.98302, 
    54.98456, 54.98582, 54.98679, 54.98748, 54.98788, 54.988, 54.98783, 
    54.98738, 54.98665, 54.98563, 54.98433, 54.98275, 54.98088, 54.97873, 
    54.97629, 54.97356, 54.97056, 54.96727, 54.9637, 54.95984, 54.9557, 
    54.95127, 54.94657, 54.94158, 54.9363, 54.93074, 54.92491, 54.91879, 
    54.91238, 54.90569, 54.89872, 54.89147, 54.88394, 54.87612, 54.86803, 
    54.85965, 54.85099, 54.84205, 54.83283, 54.82333, 54.81355, 54.80349, 
    54.79315, 54.78253, 54.77163, 54.76045, 54.74899, 54.73726, 54.72525, 
    54.71296, 54.70039, 54.68754, 54.67442, 54.66102, 54.64734, 54.63339, 
    54.61916, 54.60466, 54.58989, 54.57483, 54.55951, 54.54391, 54.52803, 
    54.51189, 54.49547, 54.47878, 54.46181, 54.44458, 54.42707, 54.4093, 
    54.39125, 54.37293, 54.35435, 54.33549, 54.31637, 54.29697, 54.27732, 
    54.25739, 54.23719, 54.21674, 54.19601, 54.17502, 54.15376, 54.13224, 
    54.11046, 54.08841, 54.0661, 54.04353, 54.02069, 53.9976, 53.97424, 
    53.95062, 53.92674, 53.90261, 53.87821, 53.85356, 53.82865, 53.80348, 
    53.77805, 53.75237, 53.72643, 53.70024, 53.6738, 53.64709, 53.62014, 
    53.59294, 53.56548, 53.53777, 53.50981, 53.4816, 53.45314, 53.42443, 
    53.39547, 53.36627, 53.33681, 53.30711, 53.27717, 53.24698, 53.21654, 
    53.18586, 53.15494, 53.12377, 53.09237, 53.06071, 53.02882, 52.99669, 
    52.96432, 52.93171, 52.89886, 52.86577, 52.83245, 52.79889, 52.76509, 
    52.73106, 52.6968, 52.6623, 52.62756, 52.5926, 52.5574, 52.52197, 
    52.48632, 52.45043, 52.41431, 52.37796, 52.34139, 52.30459, 52.26756, 
    52.23031, 52.19283, 52.15513, 52.11721, 52.07906, 52.04069, 52.00209, 
    51.96328, 51.92425, 51.88499, 51.84552, 51.80584, 51.76593, 51.7258, 
    51.68547, 51.64491, 51.60414, 51.56316, 51.52197, 51.48056, 51.43894, 
    51.39711, 51.35506, 51.31282, 51.27036, 51.22769, 51.18481, 51.14173, 
    51.09845, 51.05495,
  46.31211, 46.37172, 46.43118, 46.4905, 46.54967, 46.60871, 46.66759, 
    46.72634, 46.78493, 46.84339, 46.90169, 46.95985, 47.01786, 47.07571, 
    47.13342, 47.19098, 47.24839, 47.30565, 47.36275, 47.41971, 47.47651, 
    47.53315, 47.58964, 47.64598, 47.70216, 47.75818, 47.81404, 47.86975, 
    47.9253, 47.98069, 48.03592, 48.09098, 48.14589, 48.20063, 48.25522, 
    48.30964, 48.36389, 48.41798, 48.4719, 48.52567, 48.57926, 48.63268, 
    48.68594, 48.73903, 48.79194, 48.84469, 48.89727, 48.94967, 49.00191, 
    49.05397, 49.10585, 49.15757, 49.20911, 49.26047, 49.31165, 49.36266, 
    49.41349, 49.46415, 49.51462, 49.56491, 49.61502, 49.66496, 49.7147, 
    49.76427, 49.81365, 49.86285, 49.91187, 49.96069, 50.00934, 50.05779, 
    50.10606, 50.15414, 50.20203, 50.24973, 50.29724, 50.34456, 50.39169, 
    50.43862, 50.48536, 50.53191, 50.57826, 50.62442, 50.67038, 50.71614, 
    50.7617, 50.80707, 50.85224, 50.89721, 50.94197, 50.98654, 51.03091, 
    51.07507, 51.11903, 51.16278, 51.20633, 51.24967, 51.29281, 51.33574, 
    51.37846, 51.42097, 51.46328, 51.50537, 51.54726, 51.58894, 51.63039, 
    51.67165, 51.71268, 51.7535, 51.79411, 51.8345, 51.87467, 51.91463, 
    51.95437, 51.99389, 52.03319, 52.07227, 52.11114, 52.14978, 52.18819, 
    52.22639, 52.26437, 52.30211, 52.33964, 52.37694, 52.41401, 52.45086, 
    52.48747, 52.52386, 52.56002, 52.59595, 52.63166, 52.66713, 52.70237, 
    52.73737, 52.77215, 52.80669, 52.841, 52.87506, 52.9089, 52.9425, 
    52.97586, 53.00899, 53.04187, 53.07452, 53.10693, 53.1391, 53.17102, 
    53.20271, 53.23415, 53.26535, 53.29631, 53.32702, 53.35749, 53.38771, 
    53.41769, 53.44742, 53.4769, 53.50613, 53.53512, 53.56386, 53.59235, 
    53.62059, 53.64857, 53.67631, 53.70379, 53.73102, 53.758, 53.78472, 
    53.81119, 53.83741, 53.86337, 53.88906, 53.91451, 53.9397, 53.96463, 
    53.9893, 54.01372, 54.03787, 54.06177, 54.0854, 54.10878, 54.13189, 
    54.15474, 54.17732, 54.19965, 54.22171, 54.2435, 54.26503, 54.2863, 
    54.3073, 54.32804, 54.34851, 54.36871, 54.38864, 54.40831, 54.4277, 
    54.44683, 54.46569, 54.48428, 54.50261, 54.52065, 54.53843, 54.55594, 
    54.57317, 54.59014, 54.60683, 54.62325, 54.63939, 54.65526, 54.67085, 
    54.68618, 54.70122, 54.71599, 54.73049, 54.74471, 54.75865, 54.77232, 
    54.78571, 54.79882, 54.81165, 54.82421, 54.83649, 54.84849, 54.86021, 
    54.87165, 54.88282, 54.8937, 54.9043, 54.91462, 54.92467, 54.93443, 
    54.94391, 54.95311, 54.96203, 54.97066, 54.97902, 54.98709, 54.99488, 
    55.00239, 55.00962, 55.01656, 55.02322, 55.02959, 55.03569, 55.0415, 
    55.04702, 55.05227, 55.05722, 55.0619, 55.06629, 55.0704, 55.07422, 
    55.07775, 55.08101, 55.08398, 55.08666, 55.08906, 55.09118, 55.09301, 
    55.09455, 55.09581, 55.09678, 55.09747, 55.09788, 55.098, 55.09784, 
    55.09739, 55.09665, 55.09563, 55.09433, 55.09274, 55.09086, 55.0887, 
    55.08625, 55.08353, 55.08051, 55.07721, 55.07363, 55.06977, 55.06561, 
    55.06118, 55.05646, 55.05146, 55.04617, 55.0406, 55.03474, 55.0286, 
    55.02218, 55.01548, 55.00849, 55.00122, 54.99367, 54.98583, 54.97771, 
    54.96931, 54.96064, 54.95167, 54.94243, 54.9329, 54.9231, 54.91301, 
    54.90264, 54.89199, 54.88107, 54.86986, 54.85838, 54.84661, 54.83456, 
    54.82224, 54.80964, 54.79676, 54.78361, 54.77018, 54.75646, 54.74248, 
    54.72821, 54.71368, 54.69886, 54.68377, 54.6684, 54.65277, 54.63685, 
    54.62067, 54.60421, 54.58747, 54.57047, 54.55319, 54.53564, 54.51781, 
    54.49973, 54.48136, 54.46273, 54.44382, 54.42466, 54.40522, 54.38551, 
    54.36553, 54.34529, 54.32478, 54.304, 54.28296, 54.26165, 54.24007, 
    54.21824, 54.19613, 54.17377, 54.15114, 54.12825, 54.10509, 54.08168, 
    54.05801, 54.03407, 54.00988, 53.98542, 53.9607, 53.93573, 53.9105, 
    53.88502, 53.85928, 53.83327, 53.80702, 53.78051, 53.75375, 53.72673, 
    53.69946, 53.67194, 53.64416, 53.61613, 53.58786, 53.55933, 53.53055, 
    53.50153, 53.47225, 53.44273, 53.41296, 53.38295, 53.35268, 53.32218, 
    53.29143, 53.26043, 53.22919, 53.19771, 53.16599, 53.13402, 53.10182, 
    53.06937, 53.03669, 53.00376, 52.9706, 52.9372, 52.90356, 52.86969, 
    52.83558, 52.80124, 52.76666, 52.73185, 52.69681, 52.66153, 52.62603, 
    52.59029, 52.55432, 52.51812, 52.4817, 52.44504, 52.40816, 52.37105, 
    52.33372, 52.29616, 52.25837, 52.22036, 52.18213, 52.14368, 52.105, 
    52.06611, 52.02699, 51.98765, 51.9481, 51.90832, 51.86833, 51.82812, 
    51.7877, 51.74706, 51.7062, 51.66513, 51.62385, 51.58236, 51.54065, 
    51.49873, 51.4566, 51.41426, 51.37172, 51.32896, 51.286, 51.24283, 
    51.19945, 51.15587,
  46.40437, 46.46407, 46.52362, 46.58303, 46.6423, 46.70143, 46.76041, 
    46.81924, 46.87794, 46.93648, 46.99488, 47.05313, 47.11123, 47.16918, 
    47.22698, 47.28463, 47.34214, 47.39949, 47.45668, 47.51373, 47.57063, 
    47.62736, 47.68395, 47.74038, 47.79665, 47.85276, 47.90872, 47.96452, 
    48.02016, 48.07565, 48.13097, 48.18613, 48.24113, 48.29597, 48.35065, 
    48.40516, 48.45951, 48.51369, 48.56771, 48.62156, 48.67525, 48.72877, 
    48.78212, 48.8353, 48.88831, 48.94115, 48.99383, 49.04633, 49.09865, 
    49.15081, 49.20279, 49.25459, 49.30622, 49.35768, 49.40896, 49.46006, 
    49.51099, 49.56173, 49.6123, 49.66269, 49.71289, 49.76292, 49.81276, 
    49.86242, 49.9119, 49.96119, 50.01029, 50.05922, 50.10795, 50.1565, 
    50.20486, 50.25303, 50.30101, 50.3488, 50.39641, 50.44382, 50.49104, 
    50.53806, 50.5849, 50.63153, 50.67798, 50.72422, 50.77028, 50.81613, 
    50.86179, 50.90725, 50.9525, 50.99756, 51.04242, 51.08707, 51.13153, 
    51.17578, 51.21983, 51.26367, 51.30731, 51.35074, 51.39397, 51.43699, 
    51.4798, 51.5224, 51.56479, 51.60698, 51.64895, 51.69071, 51.73226, 
    51.77359, 51.81472, 51.85562, 51.89632, 51.93679, 51.97705, 52.01709, 
    52.05692, 52.09653, 52.13591, 52.17508, 52.21402, 52.25275, 52.29125, 
    52.32953, 52.36759, 52.40542, 52.44302, 52.4804, 52.51756, 52.55449, 
    52.59119, 52.62766, 52.6639, 52.69991, 52.73569, 52.77124, 52.80656, 
    52.84164, 52.8765, 52.91112, 52.9455, 52.97965, 53.01356, 53.04724, 
    53.08067, 53.11388, 53.14684, 53.17956, 53.21204, 53.24428, 53.27628, 
    53.30804, 53.33956, 53.37083, 53.40186, 53.43264, 53.46318, 53.49348, 
    53.52353, 53.55332, 53.58287, 53.61218, 53.64124, 53.67004, 53.6986, 
    53.7269, 53.75496, 53.78276, 53.8103, 53.8376, 53.86464, 53.89143, 
    53.91796, 53.94424, 53.97026, 53.99603, 54.02153, 54.04678, 54.07178, 
    54.09651, 54.12098, 54.1452, 54.16915, 54.19284, 54.21627, 54.23944, 
    54.26234, 54.28499, 54.30737, 54.32948, 54.35133, 54.37292, 54.39423, 
    54.41529, 54.43607, 54.45659, 54.47684, 54.49683, 54.51654, 54.53599, 
    54.55517, 54.57407, 54.59271, 54.61108, 54.62917, 54.647, 54.66455, 
    54.68182, 54.69883, 54.71556, 54.73202, 54.74821, 54.76412, 54.77975, 
    54.79511, 54.8102, 54.82501, 54.83954, 54.85379, 54.86777, 54.88148, 
    54.8949, 54.90805, 54.92091, 54.9335, 54.94581, 54.95784, 54.96959, 
    54.98106, 54.99226, 55.00317, 55.0138, 55.02415, 55.03422, 55.044, 
    55.05351, 55.06273, 55.07167, 55.08033, 55.08871, 55.0968, 55.10461, 
    55.11214, 55.11938, 55.12635, 55.13302, 55.13942, 55.14552, 55.15135, 
    55.15689, 55.16215, 55.16712, 55.17181, 55.17621, 55.18032, 55.18415, 
    55.1877, 55.19096, 55.19394, 55.19663, 55.19904, 55.20116, 55.20299, 
    55.20454, 55.2058, 55.20678, 55.20747, 55.20788, 55.208, 55.20783, 
    55.20738, 55.20665, 55.20562, 55.20432, 55.20272, 55.20084, 55.19868, 
    55.19622, 55.19349, 55.19047, 55.18716, 55.18357, 55.17969, 55.17553, 
    55.17108, 55.16635, 55.16133, 55.15603, 55.15045, 55.14458, 55.13842, 
    55.13198, 55.12526, 55.11826, 55.11097, 55.1034, 55.09554, 55.0874, 
    55.07898, 55.07028, 55.06129, 55.05202, 55.04247, 55.03264, 55.02253, 
    55.01213, 55.00146, 54.99051, 54.97927, 54.96775, 54.95596, 54.94388, 
    54.93153, 54.9189, 54.90598, 54.8928, 54.87933, 54.86558, 54.85156, 
    54.83726, 54.82268, 54.80783, 54.7927, 54.7773, 54.76162, 54.74567, 
    54.72944, 54.71294, 54.69616, 54.67911, 54.66179, 54.6442, 54.62633, 
    54.60819, 54.58978, 54.5711, 54.55215, 54.53293, 54.51344, 54.49369, 
    54.47366, 54.45337, 54.4328, 54.41198, 54.39088, 54.36952, 54.34789, 
    54.326, 54.30384, 54.28142, 54.25874, 54.23579, 54.21258, 54.18911, 
    54.16538, 54.14138, 54.11713, 54.09261, 54.06784, 54.04281, 54.01752, 
    53.99197, 53.96616, 53.9401, 53.91378, 53.88721, 53.86038, 53.8333, 
    53.80597, 53.77837, 53.75053, 53.72244, 53.6941, 53.6655, 53.63665, 
    53.60756, 53.57822, 53.54863, 53.51879, 53.4887, 53.45837, 53.42779, 
    53.39697, 53.3659, 53.33459, 53.30304, 53.27124, 53.2392, 53.20692, 
    53.1744, 53.14164, 53.10864, 53.0754, 53.04193, 53.00821, 52.97426, 
    52.94008, 52.90565, 52.871, 52.83611, 52.80099, 52.76563, 52.73005, 
    52.69423, 52.65818, 52.6219, 52.5854, 52.54866, 52.5117, 52.47451, 
    52.43709, 52.39945, 52.36158, 52.32349, 52.28518, 52.24664, 52.20788, 
    52.1689, 52.1297, 52.09027, 52.05064, 52.01078, 51.9707, 51.9304, 
    51.88989, 51.84917, 51.80822, 51.76707, 51.7257, 51.68412, 51.64232, 
    51.60032, 51.5581, 51.51567, 51.47304, 51.4302, 51.38715, 51.34389, 
    51.30042, 51.25675,
  46.49657, 46.55636, 46.616, 46.67551, 46.73487, 46.79409, 46.85316, 
    46.91209, 46.97087, 47.02951, 47.088, 47.14634, 47.20454, 47.26258, 
    47.32048, 47.37822, 47.43582, 47.49326, 47.55056, 47.60769, 47.66468, 
    47.72151, 47.77819, 47.83471, 47.89108, 47.94729, 48.00334, 48.05923, 
    48.11497, 48.17055, 48.22596, 48.28122, 48.33632, 48.39125, 48.44602, 
    48.50063, 48.55507, 48.60935, 48.66346, 48.71741, 48.77119, 48.8248, 
    48.87824, 48.93152, 48.98463, 49.03756, 49.09033, 49.14292, 49.19534, 
    49.24759, 49.29967, 49.35157, 49.40329, 49.45484, 49.50621, 49.55741, 
    49.60843, 49.65927, 49.70993, 49.76041, 49.81071, 49.86083, 49.91076, 
    49.96051, 50.01009, 50.05947, 50.10867, 50.15768, 50.20651, 50.25515, 
    50.30361, 50.35187, 50.39995, 50.44783, 50.49553, 50.54303, 50.59034, 
    50.63746, 50.68438, 50.73111, 50.77765, 50.82399, 50.87013, 50.91608, 
    50.96182, 51.00737, 51.05272, 51.09787, 51.14282, 51.18756, 51.23211, 
    51.27645, 51.32059, 51.36452, 51.40825, 51.45177, 51.49509, 51.5382, 
    51.5811, 51.62379, 51.66627, 51.70854, 51.7506, 51.79245, 51.83408, 
    51.87551, 51.91671, 51.95771, 51.99849, 52.03905, 52.0794, 52.11953, 
    52.15944, 52.19913, 52.2386, 52.27785, 52.31688, 52.35569, 52.39428, 
    52.43264, 52.47078, 52.50869, 52.54638, 52.58384, 52.62108, 52.65809, 
    52.69487, 52.73142, 52.76775, 52.80384, 52.8397, 52.87533, 52.91072, 
    52.94589, 52.98082, 53.01552, 53.04998, 53.08421, 53.11819, 53.15195, 
    53.18546, 53.21874, 53.25178, 53.28457, 53.31713, 53.34945, 53.38152, 
    53.41335, 53.44494, 53.47629, 53.50739, 53.53825, 53.56886, 53.59922, 
    53.62934, 53.65921, 53.68883, 53.7182, 53.74733, 53.7762, 53.80482, 
    53.8332, 53.86132, 53.88919, 53.9168, 53.94416, 53.97127, 53.99812, 
    54.02472, 54.05106, 54.07714, 54.10297, 54.12854, 54.15385, 54.17891, 
    54.2037, 54.22823, 54.2525, 54.27652, 54.30027, 54.32375, 54.34698, 
    54.36994, 54.39264, 54.41507, 54.43724, 54.45914, 54.48079, 54.50216, 
    54.52326, 54.5441, 54.56467, 54.58497, 54.60501, 54.62477, 54.64427, 
    54.66349, 54.68245, 54.70113, 54.71954, 54.73768, 54.75555, 54.77315, 
    54.79047, 54.80752, 54.82429, 54.84079, 54.85702, 54.87297, 54.88865, 
    54.90405, 54.91917, 54.93402, 54.94859, 54.96288, 54.97689, 54.99063, 
    55.00409, 55.01727, 55.03017, 55.04279, 55.05513, 55.06719, 55.07898, 
    55.09048, 55.1017, 55.11264, 55.12329, 55.13367, 55.14376, 55.15358, 
    55.16311, 55.17235, 55.18132, 55.19, 55.1984, 55.20651, 55.21434, 
    55.22189, 55.22915, 55.23613, 55.24282, 55.24924, 55.25536, 55.2612, 
    55.26676, 55.27203, 55.27701, 55.28171, 55.28613, 55.29025, 55.29409, 
    55.29765, 55.30092, 55.30391, 55.3066, 55.30901, 55.31114, 55.31298, 
    55.31453, 55.3158, 55.31678, 55.31747, 55.31788, 55.318, 55.31783, 
    55.31738, 55.31664, 55.31562, 55.3143, 55.31271, 55.31082, 55.30865, 
    55.30619, 55.30345, 55.30042, 55.29711, 55.29351, 55.28962, 55.28545, 
    55.28099, 55.27624, 55.27121, 55.2659, 55.2603, 55.25441, 55.24824, 
    55.24179, 55.23505, 55.22802, 55.22071, 55.21312, 55.20525, 55.19709, 
    55.18864, 55.17992, 55.17091, 55.16162, 55.15204, 55.14219, 55.13205, 
    55.12162, 55.11092, 55.09994, 55.08868, 55.07713, 55.0653, 55.0532, 
    55.04081, 55.02814, 55.0152, 55.00198, 54.98848, 54.97469, 54.96064, 
    54.9463, 54.93169, 54.91679, 54.90163, 54.88618, 54.87046, 54.85447, 
    54.8382, 54.82166, 54.80484, 54.78775, 54.77038, 54.75274, 54.73483, 
    54.71665, 54.69819, 54.67947, 54.66047, 54.6412, 54.62166, 54.60186, 
    54.58178, 54.56144, 54.54082, 54.51994, 54.49879, 54.47738, 54.4557, 
    54.43375, 54.41154, 54.38906, 54.36633, 54.34332, 54.32005, 54.29652, 
    54.27274, 54.24868, 54.22437, 54.19979, 54.17496, 54.14986, 54.12451, 
    54.0989, 54.07304, 54.04691, 54.02053, 53.99389, 53.967, 53.93985, 
    53.91245, 53.8848, 53.85689, 53.82873, 53.80032, 53.77165, 53.74274, 
    53.71357, 53.68416, 53.6545, 53.62459, 53.59443, 53.56403, 53.53338, 
    53.50249, 53.47135, 53.43996, 53.40833, 53.37646, 53.34435, 53.312, 
    53.2794, 53.24657, 53.21349, 53.18018, 53.14663, 53.11283, 53.07881, 
    53.04454, 53.01004, 52.97531, 52.94034, 52.90514, 52.86971, 52.83404, 
    52.79814, 52.76201, 52.72565, 52.68907, 52.65225, 52.6152, 52.57793, 
    52.54043, 52.50271, 52.46476, 52.42659, 52.38819, 52.34956, 52.31072, 
    52.27166, 52.23237, 52.19286, 52.15314, 52.11319, 52.07303, 52.03265, 
    51.99205, 51.95124, 51.91021, 51.86897, 51.82751, 51.78584, 51.74396, 
    51.70187, 51.65956, 51.61705, 51.57432, 51.53139, 51.48825, 51.4449, 
    51.40135, 51.35759,
  46.5887, 46.64858, 46.70832, 46.76791, 46.82737, 46.88668, 46.94585, 
    47.00487, 47.06374, 47.12247, 47.18106, 47.23949, 47.29778, 47.35592, 
    47.41391, 47.47175, 47.52944, 47.58698, 47.64436, 47.7016, 47.75867, 
    47.8156, 47.87237, 47.92899, 47.98545, 48.04175, 48.0979, 48.15389, 
    48.20972, 48.26539, 48.3209, 48.37625, 48.43144, 48.48647, 48.54133, 
    48.59603, 48.65057, 48.70494, 48.75915, 48.81319, 48.86707, 48.92077, 
    48.97431, 49.02768, 49.08088, 49.13391, 49.18678, 49.23946, 49.29198, 
    49.34432, 49.39649, 49.44848, 49.50031, 49.55195, 49.60342, 49.65471, 
    49.70582, 49.75675, 49.80751, 49.85808, 49.90847, 49.95868, 50.00871, 
    50.05856, 50.10822, 50.1577, 50.207, 50.2561, 50.30503, 50.35376, 
    50.40231, 50.45066, 50.49883, 50.54681, 50.5946, 50.64219, 50.6896, 
    50.73681, 50.78382, 50.83065, 50.87727, 50.92371, 50.96994, 51.01598, 
    51.06182, 51.10746, 51.1529, 51.19814, 51.24318, 51.28801, 51.33265, 
    51.37708, 51.42131, 51.46533, 51.50915, 51.55276, 51.59616, 51.63936, 
    51.68235, 51.72513, 51.7677, 51.81006, 51.85221, 51.89415, 51.93587, 
    51.97738, 52.01868, 52.05976, 52.10062, 52.14127, 52.18171, 52.22192, 
    52.26191, 52.30169, 52.34125, 52.38058, 52.4197, 52.4586, 52.49726, 
    52.53571, 52.57393, 52.61193, 52.6497, 52.68725, 52.72457, 52.76166, 
    52.79852, 52.83516, 52.87156, 52.90773, 52.94367, 52.97939, 53.01486, 
    53.05011, 53.08511, 53.11989, 53.15443, 53.18874, 53.2228, 53.25663, 
    53.29022, 53.32357, 53.35669, 53.38956, 53.4222, 53.45459, 53.48674, 
    53.51864, 53.5503, 53.58172, 53.6129, 53.64383, 53.67451, 53.70494, 
    53.73513, 53.76507, 53.79477, 53.82421, 53.8534, 53.88234, 53.91104, 
    53.93948, 53.96766, 53.9956, 54.02328, 54.0507, 54.07788, 54.1048, 
    54.13146, 54.15786, 54.18401, 54.2099, 54.23553, 54.2609, 54.28602, 
    54.31087, 54.33546, 54.3598, 54.38387, 54.40768, 54.43122, 54.45451, 
    54.47752, 54.50028, 54.52277, 54.54499, 54.56695, 54.58864, 54.61007, 
    54.63123, 54.65212, 54.67274, 54.69309, 54.71318, 54.73299, 54.75253, 
    54.77181, 54.79081, 54.80954, 54.828, 54.84619, 54.8641, 54.88174, 
    54.89911, 54.9162, 54.93302, 54.94956, 54.96582, 54.98182, 54.99753, 
    55.01297, 55.02813, 55.04302, 55.05762, 55.07195, 55.08601, 55.09978, 
    55.11327, 55.12648, 55.13942, 55.15207, 55.16444, 55.17654, 55.18835, 
    55.19988, 55.21113, 55.2221, 55.23278, 55.24319, 55.25331, 55.26315, 
    55.2727, 55.28197, 55.29096, 55.29966, 55.30808, 55.31622, 55.32407, 
    55.33164, 55.33892, 55.34592, 55.35263, 55.35905, 55.3652, 55.37105, 
    55.37662, 55.3819, 55.3869, 55.39161, 55.39604, 55.40018, 55.40403, 
    55.4076, 55.41087, 55.41387, 55.41657, 55.41899, 55.42112, 55.42297, 
    55.42452, 55.42579, 55.42677, 55.42747, 55.42788, 55.428, 55.42783, 
    55.42738, 55.42664, 55.42561, 55.42429, 55.42269, 55.4208, 55.41863, 
    55.41616, 55.41341, 55.41037, 55.40705, 55.40344, 55.39954, 55.39536, 
    55.39089, 55.38613, 55.38109, 55.37576, 55.37014, 55.36425, 55.35806, 
    55.35159, 55.34483, 55.33779, 55.33046, 55.32285, 55.31495, 55.30677, 
    55.29831, 55.28956, 55.28053, 55.27121, 55.26161, 55.25172, 55.24156, 
    55.23111, 55.22038, 55.20937, 55.19808, 55.1865, 55.17464, 55.16251, 
    55.15009, 55.13739, 55.12441, 55.11116, 55.09762, 55.0838, 55.06971, 
    55.05533, 55.04068, 55.02575, 55.01055, 54.99506, 54.97931, 54.96327, 
    54.94696, 54.93037, 54.91351, 54.89638, 54.87897, 54.86129, 54.84333, 
    54.8251, 54.80659, 54.78782, 54.76878, 54.74946, 54.72987, 54.71002, 
    54.68989, 54.66949, 54.64883, 54.6279, 54.6067, 54.58523, 54.5635, 
    54.54149, 54.51923, 54.4967, 54.4739, 54.45084, 54.42751, 54.40393, 
    54.38008, 54.35596, 54.33159, 54.30696, 54.28206, 54.25691, 54.23149, 
    54.20582, 54.17989, 54.1537, 54.12726, 54.10056, 54.0736, 54.04639, 
    54.01892, 53.9912, 53.96322, 53.93499, 53.90651, 53.87778, 53.8488, 
    53.81957, 53.79008, 53.76035, 53.73037, 53.70015, 53.66967, 53.63895, 
    53.60798, 53.57677, 53.54531, 53.51361, 53.48167, 53.44948, 53.41705, 
    53.38438, 53.35147, 53.31832, 53.28492, 53.2513, 53.21743, 53.18332, 
    53.14898, 53.11441, 53.07959, 53.04454, 53.00927, 52.97375, 52.938, 
    52.90203, 52.86581, 52.82938, 52.79271, 52.75581, 52.71868, 52.68132, 
    52.64375, 52.60593, 52.5679, 52.52964, 52.49116, 52.45246, 52.41353, 
    52.37438, 52.33501, 52.29541, 52.2556, 52.21557, 52.17532, 52.13486, 
    52.09417, 52.05327, 52.01216, 51.97083, 51.92928, 51.88753, 51.84555, 
    51.80338, 51.76098, 51.71838, 51.67556, 51.63254, 51.58931, 51.54588, 
    51.50223, 51.45838,
  46.68076, 46.74073, 46.80057, 46.86026, 46.9198, 46.97921, 47.03847, 
    47.09758, 47.15655, 47.21537, 47.27405, 47.33258, 47.39096, 47.44919, 
    47.50727, 47.56521, 47.62299, 47.68062, 47.7381, 47.79543, 47.8526, 
    47.90963, 47.96649, 48.0232, 48.07975, 48.13615, 48.19239, 48.24848, 
    48.3044, 48.36017, 48.41578, 48.47122, 48.5265, 48.58162, 48.63659, 
    48.69138, 48.74601, 48.80048, 48.85478, 48.90892, 48.96289, 49.01669, 
    49.07032, 49.12379, 49.17708, 49.23021, 49.28316, 49.33595, 49.38855, 
    49.44099, 49.49326, 49.54535, 49.59726, 49.649, 49.70056, 49.75195, 
    49.80315, 49.85418, 49.90503, 49.9557, 50.00618, 50.05649, 50.10661, 
    50.15656, 50.20631, 50.25589, 50.30527, 50.35447, 50.40349, 50.45232, 
    50.50096, 50.54941, 50.59767, 50.64574, 50.69362, 50.74131, 50.78881, 
    50.83611, 50.88322, 50.93013, 50.97685, 51.02338, 51.0697, 51.11583, 
    51.16176, 51.20749, 51.25303, 51.29836, 51.34349, 51.38842, 51.43314, 
    51.47766, 51.52198, 51.5661, 51.61, 51.65371, 51.6972, 51.74049, 
    51.78357, 51.82644, 51.86909, 51.91154, 51.95378, 51.9958, 52.03762, 
    52.07921, 52.1206, 52.16177, 52.20272, 52.24345, 52.28397, 52.32428, 
    52.36436, 52.40422, 52.44386, 52.48329, 52.52249, 52.56146, 52.60022, 
    52.63875, 52.67706, 52.71514, 52.75299, 52.79062, 52.82803, 52.8652, 
    52.90214, 52.93886, 52.97534, 53.0116, 53.04762, 53.08341, 53.11897, 
    53.15429, 53.18938, 53.22424, 53.25885, 53.29324, 53.32738, 53.36129, 
    53.39496, 53.42839, 53.46158, 53.49453, 53.52723, 53.5597, 53.59192, 
    53.62391, 53.65564, 53.68713, 53.71838, 53.74938, 53.78014, 53.81065, 
    53.8409, 53.87092, 53.90068, 53.93019, 53.95945, 53.98847, 54.01723, 
    54.04573, 54.07399, 54.10199, 54.12974, 54.15723, 54.18447, 54.21145, 
    54.23818, 54.26465, 54.29086, 54.31681, 54.34251, 54.36794, 54.39312, 
    54.41803, 54.44268, 54.46708, 54.49121, 54.51507, 54.53868, 54.56202, 
    54.58509, 54.6079, 54.63045, 54.65273, 54.67474, 54.69649, 54.71797, 
    54.73918, 54.76012, 54.7808, 54.8012, 54.82133, 54.8412, 54.86079, 
    54.88012, 54.89917, 54.91794, 54.93645, 54.95468, 54.97264, 54.99033, 
    55.00774, 55.02487, 55.04173, 55.05832, 55.07463, 55.09066, 55.10641, 
    55.12189, 55.13709, 55.15202, 55.16666, 55.18103, 55.19511, 55.20892, 
    55.22245, 55.2357, 55.24866, 55.26135, 55.27376, 55.28588, 55.29773, 
    55.30928, 55.32056, 55.33156, 55.34227, 55.3527, 55.36285, 55.37271, 
    55.38229, 55.39159, 55.4006, 55.40933, 55.41777, 55.42593, 55.4338, 
    55.44138, 55.44868, 55.4557, 55.46243, 55.46888, 55.47503, 55.4809, 
    55.48649, 55.49178, 55.4968, 55.50152, 55.50595, 55.51011, 55.51397, 
    55.51754, 55.52083, 55.52383, 55.52654, 55.52896, 55.53111, 55.53295, 
    55.53451, 55.53579, 55.53677, 55.53747, 55.53788, 55.538, 55.53783, 
    55.53738, 55.53664, 55.5356, 55.53429, 55.53268, 55.53078, 55.5286, 
    55.52613, 55.52337, 55.52033, 55.51699, 55.51337, 55.50947, 55.50527, 
    55.50079, 55.49602, 55.49097, 55.48562, 55.47999, 55.47408, 55.46787, 
    55.46138, 55.45461, 55.44755, 55.4402, 55.43257, 55.42466, 55.41645, 
    55.40797, 55.39919, 55.39014, 55.3808, 55.37117, 55.36126, 55.35107, 
    55.3406, 55.32984, 55.3188, 55.30748, 55.29587, 55.28398, 55.27181, 
    55.25936, 55.24663, 55.23362, 55.22033, 55.20676, 55.19291, 55.17877, 
    55.16436, 55.14967, 55.13471, 55.11946, 55.10394, 55.08814, 55.07206, 
    55.05571, 55.03908, 55.02218, 55.005, 54.98755, 54.96982, 54.95182, 
    54.93354, 54.91499, 54.89617, 54.87708, 54.85771, 54.83807, 54.81817, 
    54.79799, 54.77754, 54.75683, 54.73584, 54.71459, 54.69307, 54.67128, 
    54.64922, 54.6269, 54.60431, 54.58146, 54.55834, 54.53496, 54.51131, 
    54.48741, 54.46323, 54.4388, 54.41411, 54.38915, 54.36393, 54.33846, 
    54.31273, 54.28673, 54.26048, 54.23397, 54.2072, 54.18018, 54.1529, 
    54.12537, 54.09758, 54.06954, 54.04124, 54.0127, 53.98389, 53.95484, 
    53.92554, 53.89599, 53.86618, 53.83614, 53.80584, 53.77529, 53.7445, 
    53.71346, 53.68217, 53.65064, 53.61886, 53.58684, 53.55458, 53.52208, 
    53.48933, 53.45634, 53.42311, 53.38965, 53.35594, 53.32199, 53.28782, 
    53.2534, 53.21874, 53.18385, 53.14872, 53.11336, 53.07776, 53.04194, 
    53.00588, 52.96959, 52.93307, 52.89631, 52.85933, 52.82212, 52.78469, 
    52.74702, 52.70913, 52.67101, 52.63267, 52.5941, 52.55531, 52.5163, 
    52.47707, 52.43761, 52.39793, 52.35803, 52.31792, 52.27758, 52.23703, 
    52.19625, 52.15527, 52.11407, 52.07265, 52.03102, 51.98917, 51.94711, 
    51.90484, 51.86236, 51.81967, 51.77676, 51.73365, 51.69033, 51.64681, 
    51.60307, 51.55913,
  46.77275, 46.83282, 46.89275, 46.95253, 47.01217, 47.07167, 47.13102, 
    47.19023, 47.24929, 47.30821, 47.36698, 47.4256, 47.48407, 47.5424, 
    47.60058, 47.6586, 47.71648, 47.77421, 47.83178, 47.8892, 47.94647, 
    48.00359, 48.06055, 48.11735, 48.174, 48.23049, 48.28683, 48.34301, 
    48.39902, 48.45489, 48.51059, 48.56613, 48.62151, 48.67672, 48.73178, 
    48.78667, 48.84139, 48.89595, 48.95035, 49.00459, 49.05865, 49.11255, 
    49.16628, 49.21983, 49.27322, 49.32644, 49.37949, 49.43237, 49.48508, 
    49.53761, 49.58997, 49.64215, 49.69416, 49.74599, 49.79765, 49.84913, 
    49.90043, 49.95155, 50.0025, 50.05326, 50.10384, 50.15424, 50.20446, 
    50.2545, 50.30435, 50.35402, 50.4035, 50.45279, 50.5019, 50.55082, 
    50.59956, 50.6481, 50.69646, 50.74462, 50.79259, 50.84038, 50.88797, 
    50.93536, 50.98256, 51.02957, 51.07639, 51.123, 51.16942, 51.21564, 
    51.26166, 51.30749, 51.35311, 51.39853, 51.44376, 51.48878, 51.53359, 
    51.57821, 51.62262, 51.66682, 51.71082, 51.75461, 51.79819, 51.84157, 
    51.88474, 51.9277, 51.97045, 52.01299, 52.05531, 52.09742, 52.13932, 
    52.18101, 52.22248, 52.26374, 52.30478, 52.3456, 52.38621, 52.4266, 
    52.46677, 52.50671, 52.54644, 52.58595, 52.62524, 52.6643, 52.70314, 
    52.74176, 52.78015, 52.81831, 52.85625, 52.89396, 52.93145, 52.9687, 
    53.00573, 53.04253, 53.0791, 53.11543, 53.15154, 53.18741, 53.22305, 
    53.25845, 53.29362, 53.32855, 53.36325, 53.39771, 53.43193, 53.46592, 
    53.49966, 53.53317, 53.56644, 53.59946, 53.63225, 53.66479, 53.69709, 
    53.72915, 53.76096, 53.79252, 53.82384, 53.85492, 53.88574, 53.91632, 
    53.94666, 53.97674, 54.00657, 54.03616, 54.06549, 54.09457, 54.1234, 
    54.15197, 54.1803, 54.20837, 54.23618, 54.26374, 54.29105, 54.31809, 
    54.34488, 54.37141, 54.39769, 54.42371, 54.44946, 54.47496, 54.5002, 
    54.52517, 54.54989, 54.57434, 54.59853, 54.62246, 54.64612, 54.66952, 
    54.69265, 54.71552, 54.73812, 54.76046, 54.78252, 54.80433, 54.82586, 
    54.84712, 54.86812, 54.88884, 54.9093, 54.92949, 54.9494, 54.96904, 
    54.98841, 55.00751, 55.02634, 55.04489, 55.06317, 55.08117, 55.0989, 
    55.11636, 55.13354, 55.15044, 55.16707, 55.18342, 55.19949, 55.21529, 
    55.23081, 55.24605, 55.26101, 55.27569, 55.29009, 55.30422, 55.31806, 
    55.33162, 55.34491, 55.35791, 55.37062, 55.38306, 55.39522, 55.40709, 
    55.41869, 55.42999, 55.44102, 55.45176, 55.46222, 55.47239, 55.48228, 
    55.49188, 55.5012, 55.51024, 55.51899, 55.52745, 55.53563, 55.54352, 
    55.55113, 55.55845, 55.56548, 55.57223, 55.57869, 55.58487, 55.59075, 
    55.59635, 55.60166, 55.60669, 55.61142, 55.61587, 55.62003, 55.62391, 
    55.62749, 55.63078, 55.63379, 55.63651, 55.63894, 55.64109, 55.64294, 
    55.6445, 55.64578, 55.64677, 55.64747, 55.64788, 55.648, 55.64783, 
    55.64738, 55.64663, 55.6456, 55.64428, 55.64267, 55.64077, 55.63858, 
    55.6361, 55.63334, 55.63028, 55.62694, 55.62331, 55.61939, 55.61518, 
    55.61069, 55.60591, 55.60084, 55.59549, 55.58984, 55.58391, 55.57769, 
    55.57118, 55.56439, 55.55731, 55.54995, 55.54229, 55.53436, 55.52613, 
    55.51762, 55.50883, 55.49975, 55.49038, 55.48073, 55.4708, 55.46058, 
    55.45008, 55.43929, 55.42822, 55.41687, 55.40524, 55.39331, 55.38111, 
    55.36863, 55.35587, 55.34282, 55.3295, 55.31589, 55.302, 55.28783, 
    55.27339, 55.25866, 55.24366, 55.22837, 55.21281, 55.19697, 55.18085, 
    55.16446, 55.14779, 55.13084, 55.11361, 55.09612, 55.07834, 55.0603, 
    55.04197, 55.02338, 55.00451, 54.98537, 54.96595, 54.94627, 54.92631, 
    54.90608, 54.88558, 54.86481, 54.84378, 54.82247, 54.80089, 54.77905, 
    54.75694, 54.73456, 54.71192, 54.68901, 54.66583, 54.6424, 54.61869, 
    54.59472, 54.57049, 54.546, 54.52124, 54.49622, 54.47095, 54.44541, 
    54.41961, 54.39355, 54.36724, 54.34066, 54.31383, 54.28674, 54.2594, 
    54.2318, 54.20394, 54.17583, 54.14747, 54.11885, 54.08998, 54.06086, 
    54.03149, 54.00187, 53.972, 53.94188, 53.9115, 53.88088, 53.85002, 
    53.8189, 53.78754, 53.75594, 53.72409, 53.692, 53.65966, 53.62708, 
    53.59426, 53.56119, 53.52789, 53.49434, 53.46056, 53.42654, 53.39228, 
    53.35778, 53.32304, 53.28807, 53.25286, 53.21742, 53.18175, 53.14584, 
    53.1097, 53.07333, 53.03672, 52.99989, 52.96283, 52.92553, 52.88801, 
    52.85027, 52.81229, 52.77409, 52.73566, 52.69701, 52.65813, 52.61904, 
    52.57972, 52.54017, 52.50041, 52.46043, 52.42022, 52.3798, 52.33916, 
    52.2983, 52.25723, 52.21593, 52.17443, 52.13271, 52.09077, 52.04863, 
    52.00627, 51.9637, 51.92092, 51.87793, 51.83472, 51.79131, 51.7477, 
    51.70387, 51.65984,
  46.86469, 46.92484, 46.98486, 47.04474, 47.10447, 47.16406, 47.22351, 
    47.28281, 47.34196, 47.40097, 47.45984, 47.51855, 47.57713, 47.63554, 
    47.69382, 47.75194, 47.80991, 47.86773, 47.9254, 47.98291, 48.04028, 
    48.09748, 48.15454, 48.21144, 48.26818, 48.32477, 48.3812, 48.43747, 
    48.49359, 48.54954, 48.60534, 48.66097, 48.71645, 48.77176, 48.82691, 
    48.88189, 48.93671, 48.99137, 49.04586, 49.10019, 49.15435, 49.20834, 
    49.26217, 49.31582, 49.36931, 49.42262, 49.47577, 49.52874, 49.58154, 
    49.63417, 49.68662, 49.7389, 49.791, 49.84293, 49.89469, 49.94626, 
    49.99766, 50.04887, 50.09991, 50.15077, 50.20145, 50.25194, 50.30225, 
    50.35239, 50.40233, 50.45209, 50.50167, 50.55106, 50.60026, 50.64928, 
    50.6981, 50.74674, 50.79519, 50.84345, 50.89152, 50.93939, 50.98708, 
    51.03456, 51.08186, 51.12896, 51.17587, 51.22258, 51.26909, 51.3154, 
    51.36152, 51.40743, 51.45315, 51.49866, 51.54398, 51.58909, 51.634, 
    51.6787, 51.72321, 51.7675, 51.81159, 51.85547, 51.89915, 51.94261, 
    51.98587, 52.02892, 52.07176, 52.11438, 52.1568, 52.199, 52.24099, 
    52.28277, 52.32433, 52.36567, 52.4068, 52.44771, 52.4884, 52.52888, 
    52.56914, 52.60917, 52.64899, 52.68858, 52.72795, 52.7671, 52.80603, 
    52.84473, 52.8832, 52.92145, 52.95948, 52.99727, 53.03484, 53.07218, 
    53.10929, 53.14617, 53.18282, 53.21923, 53.25542, 53.29137, 53.32709, 
    53.36258, 53.39783, 53.43284, 53.46762, 53.50216, 53.53646, 53.57052, 
    53.60435, 53.63793, 53.67128, 53.70438, 53.73724, 53.76986, 53.80223, 
    53.83436, 53.86625, 53.89788, 53.92928, 53.96043, 53.99133, 54.02198, 
    54.05238, 54.08254, 54.11244, 54.1421, 54.1715, 54.20065, 54.22955, 
    54.25819, 54.28658, 54.31472, 54.3426, 54.37023, 54.3976, 54.42471, 
    54.45157, 54.47817, 54.50451, 54.53059, 54.55641, 54.58197, 54.60727, 
    54.6323, 54.65708, 54.68159, 54.70584, 54.72982, 54.75355, 54.777, 
    54.80019, 54.82312, 54.84578, 54.86817, 54.89029, 54.91215, 54.93373, 
    54.95505, 54.9761, 54.99688, 55.01739, 55.03762, 55.05759, 55.07728, 
    55.0967, 55.11585, 55.13472, 55.15332, 55.17165, 55.1897, 55.20747, 
    55.22497, 55.2422, 55.25914, 55.27581, 55.29221, 55.30832, 55.32416, 
    55.33971, 55.355, 55.37, 55.38472, 55.39915, 55.41331, 55.4272, 55.44079, 
    55.45411, 55.46714, 55.4799, 55.49237, 55.50455, 55.51646, 55.52808, 
    55.53942, 55.55047, 55.56124, 55.57173, 55.58193, 55.59184, 55.60147, 
    55.61082, 55.61987, 55.62865, 55.63713, 55.64533, 55.65325, 55.66087, 
    55.66821, 55.67527, 55.68203, 55.68851, 55.6947, 55.7006, 55.70621, 
    55.71154, 55.71658, 55.72132, 55.72578, 55.72996, 55.73384, 55.73743, 
    55.74074, 55.74376, 55.74648, 55.74892, 55.75107, 55.75293, 55.75449, 
    55.75578, 55.75676, 55.75747, 55.75788, 55.758, 55.75783, 55.75737, 
    55.75663, 55.75559, 55.75426, 55.75265, 55.75075, 55.74855, 55.74607, 
    55.7433, 55.74023, 55.73689, 55.73325, 55.72932, 55.7251, 55.72059, 
    55.7158, 55.71072, 55.70535, 55.69968, 55.69374, 55.6875, 55.68098, 
    55.67417, 55.66707, 55.65969, 55.65202, 55.64405, 55.63581, 55.62728, 
    55.61846, 55.60936, 55.59997, 55.59029, 55.58033, 55.57009, 55.55956, 
    55.54874, 55.53764, 55.52626, 55.5146, 55.50265, 55.49041, 55.4779, 
    55.4651, 55.45202, 55.43866, 55.42502, 55.41109, 55.39689, 55.3824, 
    55.36764, 55.3526, 55.33727, 55.32167, 55.30579, 55.28963, 55.27319, 
    55.25648, 55.23949, 55.22222, 55.20468, 55.18686, 55.16877, 55.1504, 
    55.13175, 55.11283, 55.09365, 55.07418, 55.05445, 55.03444, 55.01416, 
    54.99361, 54.97279, 54.9517, 54.93034, 54.90871, 54.88681, 54.86464, 
    54.84221, 54.81951, 54.79654, 54.77331, 54.74981, 54.72605, 54.70202, 
    54.67773, 54.65318, 54.62836, 54.60328, 54.57794, 54.55234, 54.52648, 
    54.50036, 54.47398, 54.44734, 54.42044, 54.39329, 54.36588, 54.33821, 
    54.31029, 54.28211, 54.25368, 54.22499, 54.19606, 54.16687, 54.13742, 
    54.10773, 54.07779, 54.04759, 54.01715, 53.98646, 53.95552, 53.92433, 
    53.8929, 53.86122, 53.82929, 53.79712, 53.76471, 53.73206, 53.69916, 
    53.66602, 53.63263, 53.59901, 53.56515, 53.53105, 53.49671, 53.46213, 
    53.42732, 53.39227, 53.35698, 53.32146, 53.2857, 53.24971, 53.21349, 
    53.17704, 53.14035, 53.10344, 53.06629, 53.02891, 52.99131, 52.95348, 
    52.91542, 52.87713, 52.83862, 52.79988, 52.76092, 52.72174, 52.68233, 
    52.6427, 52.60285, 52.56278, 52.52249, 52.48198, 52.44125, 52.40031, 
    52.35915, 52.31777, 52.27617, 52.23436, 52.19234, 52.1501, 52.10766, 
    52.06499, 52.02213, 51.97904, 51.93575, 51.89225, 51.84855, 51.80463, 
    51.76051,
  46.95654, 47.0168, 47.07691, 47.13688, 47.1967, 47.25639, 47.31593, 
    47.37532, 47.43457, 47.49368, 47.55264, 47.61145, 47.67011, 47.72862, 
    47.78699, 47.8452, 47.90327, 47.96119, 48.01895, 48.07656, 48.13401, 
    48.19132, 48.24847, 48.30546, 48.3623, 48.41898, 48.47551, 48.53188, 
    48.58809, 48.64414, 48.70003, 48.75576, 48.81133, 48.86673, 48.92198, 
    48.97706, 49.03198, 49.08673, 49.14132, 49.19574, 49.24999, 49.30408, 
    49.358, 49.41175, 49.46533, 49.51875, 49.57198, 49.62505, 49.67795, 
    49.73067, 49.78322, 49.83559, 49.88779, 49.93982, 49.99166, 50.04333, 
    50.09483, 50.14614, 50.19727, 50.24823, 50.299, 50.34959, 50.39999, 
    50.45022, 50.50026, 50.55012, 50.59979, 50.64927, 50.69857, 50.74768, 
    50.7966, 50.84534, 50.89388, 50.94223, 50.99039, 51.03836, 51.08614, 
    51.13372, 51.18111, 51.22831, 51.2753, 51.32211, 51.36871, 51.41512, 
    51.46133, 51.50734, 51.55314, 51.59875, 51.64416, 51.68936, 51.73436, 
    51.77916, 51.82375, 51.86814, 51.91232, 51.95629, 52.00006, 52.04361, 
    52.08696, 52.1301, 52.17303, 52.21574, 52.25825, 52.30054, 52.34262, 
    52.38448, 52.42613, 52.46757, 52.50878, 52.54978, 52.59056, 52.63113, 
    52.67147, 52.71159, 52.7515, 52.79118, 52.83063, 52.86987, 52.90888, 
    52.94766, 52.98623, 53.02456, 53.06267, 53.10055, 53.1382, 53.17562, 
    53.21281, 53.24978, 53.28651, 53.32301, 53.35928, 53.39531, 53.43111, 
    53.46667, 53.50201, 53.5371, 53.57196, 53.60658, 53.64096, 53.6751, 
    53.709, 53.74266, 53.77608, 53.80926, 53.8422, 53.87489, 53.90734, 
    53.93955, 53.97151, 54.00323, 54.03469, 54.06591, 54.09689, 54.12761, 
    54.15809, 54.18832, 54.21829, 54.24802, 54.27749, 54.30671, 54.33568, 
    54.36439, 54.39285, 54.42106, 54.44901, 54.4767, 54.50414, 54.53132, 
    54.55824, 54.5849, 54.61131, 54.63745, 54.66333, 54.68896, 54.71432, 
    54.73942, 54.76425, 54.78883, 54.81314, 54.83718, 54.86096, 54.88448, 
    54.90772, 54.93071, 54.95342, 54.97587, 54.99805, 55.01996, 55.0416, 
    55.06297, 55.08407, 55.1049, 55.12546, 55.14575, 55.16577, 55.18551, 
    55.20498, 55.22417, 55.2431, 55.26175, 55.28012, 55.29821, 55.31603, 
    55.33358, 55.35085, 55.36784, 55.38455, 55.40099, 55.41714, 55.43302, 
    55.44862, 55.46394, 55.47898, 55.49374, 55.50821, 55.52241, 55.53632, 
    55.54996, 55.56331, 55.57638, 55.58916, 55.60167, 55.61389, 55.62582, 
    55.63747, 55.64884, 55.65992, 55.67072, 55.68123, 55.69146, 55.7014, 
    55.71106, 55.72042, 55.72951, 55.7383, 55.74681, 55.75504, 55.76297, 
    55.77062, 55.77798, 55.78505, 55.79183, 55.79832, 55.80453, 55.81045, 
    55.81608, 55.82141, 55.82647, 55.83123, 55.8357, 55.83988, 55.84378, 
    55.84738, 55.85069, 55.85372, 55.85645, 55.85889, 55.86105, 55.86291, 
    55.86449, 55.86577, 55.86676, 55.86747, 55.86788, 55.868, 55.86783, 
    55.86737, 55.86662, 55.86559, 55.86425, 55.86264, 55.86073, 55.85853, 
    55.85604, 55.85326, 55.85019, 55.84683, 55.84318, 55.83924, 55.83501, 
    55.83049, 55.82569, 55.82059, 55.8152, 55.80953, 55.80357, 55.79732, 
    55.79078, 55.78395, 55.77683, 55.76942, 55.76173, 55.75375, 55.74549, 
    55.73693, 55.72809, 55.71896, 55.70955, 55.69985, 55.68986, 55.67959, 
    55.66903, 55.65819, 55.64706, 55.63565, 55.62395, 55.61197, 55.59971, 
    55.58716, 55.57433, 55.56121, 55.54782, 55.53414, 55.52018, 55.50594, 
    55.49142, 55.47662, 55.46153, 55.44617, 55.43053, 55.4146, 55.3984, 
    55.38192, 55.36517, 55.34813, 55.33082, 55.31323, 55.29537, 55.27723, 
    55.25881, 55.24012, 55.22116, 55.20192, 55.1824, 55.16262, 55.14256, 
    55.12223, 55.10163, 55.08075, 55.05961, 55.03819, 55.01651, 54.99456, 
    54.97234, 54.94984, 54.92709, 54.90406, 54.88078, 54.85722, 54.83339, 
    54.80931, 54.78496, 54.76034, 54.73546, 54.71032, 54.68492, 54.65926, 
    54.63333, 54.60715, 54.5807, 54.554, 54.52703, 54.49981, 54.47234, 
    54.4446, 54.41661, 54.38837, 54.35987, 54.33111, 54.3021, 54.27285, 
    54.24333, 54.21357, 54.18355, 54.15329, 54.12277, 54.09201, 54.06099, 
    54.02973, 53.99823, 53.96647, 53.93447, 53.90223, 53.86974, 53.83701, 
    53.80403, 53.77081, 53.73735, 53.70366, 53.66971, 53.63553, 53.60112, 
    53.56646, 53.53156, 53.49643, 53.46107, 53.42546, 53.38963, 53.35355, 
    53.31725, 53.28072, 53.24395, 53.20695, 53.16972, 53.13226, 53.09457, 
    53.05665, 53.01851, 52.98014, 52.94154, 52.90272, 52.86367, 52.82441, 
    52.78491, 52.7452, 52.70526, 52.6651, 52.62473, 52.58413, 52.54331, 
    52.50228, 52.46103, 52.41956, 52.37788, 52.33598, 52.29387, 52.25154, 
    52.209, 52.16625, 52.12329, 52.08012, 52.03674, 51.99314, 51.94935, 
    51.90534, 51.86113,
  47.04834, 47.10868, 47.16888, 47.22895, 47.28887, 47.34864, 47.40828, 
    47.46777, 47.52711, 47.58631, 47.64536, 47.70427, 47.76302, 47.82163, 
    47.88009, 47.9384, 47.99656, 48.05457, 48.11243, 48.17014, 48.22769, 
    48.28509, 48.34233, 48.39942, 48.45636, 48.51313, 48.56976, 48.62622, 
    48.68252, 48.73867, 48.79465, 48.85048, 48.90614, 48.96165, 49.01699, 
    49.07216, 49.12718, 49.18203, 49.23671, 49.29123, 49.34558, 49.39976, 
    49.45378, 49.50762, 49.5613, 49.61481, 49.66814, 49.72131, 49.7743, 
    49.82712, 49.87976, 49.93223, 49.98453, 50.03665, 50.08859, 50.14035, 
    50.19194, 50.24335, 50.29458, 50.34563, 50.39649, 50.44718, 50.49768, 
    50.548, 50.59814, 50.64809, 50.69785, 50.74743, 50.79683, 50.84603, 
    50.89505, 50.94387, 50.99252, 51.04096, 51.08922, 51.13728, 51.18515, 
    51.23283, 51.28031, 51.3276, 51.37469, 51.42159, 51.46828, 51.51479, 
    51.56108, 51.60719, 51.65309, 51.69879, 51.74429, 51.78959, 51.83468, 
    51.87957, 51.92425, 51.96873, 52.013, 52.05706, 52.10092, 52.14457, 
    52.18801, 52.23124, 52.27426, 52.31707, 52.35966, 52.40204, 52.44421, 
    52.48616, 52.5279, 52.56942, 52.61073, 52.65181, 52.69268, 52.73333, 
    52.77377, 52.81398, 52.85397, 52.89373, 52.93328, 52.9726, 53.01169, 
    53.05056, 53.08921, 53.12763, 53.16582, 53.20379, 53.24152, 53.27903, 
    53.31631, 53.35336, 53.39017, 53.42675, 53.4631, 53.49922, 53.5351, 
    53.57074, 53.60616, 53.64133, 53.67627, 53.71096, 53.74543, 53.77965, 
    53.81363, 53.84737, 53.88087, 53.91412, 53.94714, 53.97991, 54.01243, 
    54.04472, 54.07675, 54.10854, 54.14008, 54.17138, 54.20243, 54.23322, 
    54.26377, 54.29407, 54.32412, 54.35392, 54.38346, 54.41275, 54.44179, 
    54.47057, 54.4991, 54.52737, 54.55539, 54.58315, 54.61066, 54.6379, 
    54.66489, 54.69162, 54.71809, 54.7443, 54.77024, 54.79593, 54.82135, 
    54.84652, 54.87141, 54.89605, 54.92042, 54.94452, 54.96836, 54.99194, 
    55.01524, 55.03828, 55.06105, 55.08356, 55.10579, 55.12776, 55.14945, 
    55.17088, 55.19204, 55.21292, 55.23353, 55.25387, 55.27393, 55.29373, 
    55.31325, 55.33249, 55.35146, 55.37016, 55.38858, 55.40672, 55.42459, 
    55.44218, 55.45949, 55.47652, 55.49328, 55.50976, 55.52596, 55.54187, 
    55.55751, 55.57287, 55.58795, 55.60275, 55.61726, 55.6315, 55.64545, 
    55.65912, 55.6725, 55.68561, 55.69843, 55.71096, 55.72321, 55.73518, 
    55.74686, 55.75826, 55.76937, 55.7802, 55.79074, 55.80099, 55.81096, 
    55.82064, 55.83004, 55.83914, 55.84796, 55.85649, 55.86473, 55.87269, 
    55.88036, 55.88774, 55.89482, 55.90163, 55.90814, 55.91436, 55.9203, 
    55.92594, 55.93129, 55.93636, 55.94113, 55.94561, 55.94981, 55.95371, 
    55.95732, 55.96065, 55.96368, 55.96642, 55.96887, 55.97103, 55.9729, 
    55.97448, 55.97576, 55.97676, 55.97746, 55.97787, 55.978, 55.97783, 
    55.97737, 55.97662, 55.97558, 55.97425, 55.97262, 55.97071, 55.9685, 
    55.96601, 55.96322, 55.96014, 55.95677, 55.95311, 55.94917, 55.94492, 
    55.9404, 55.93557, 55.93047, 55.92506, 55.91938, 55.91339, 55.90713, 
    55.90057, 55.89372, 55.88659, 55.87917, 55.87145, 55.86345, 55.85516, 
    55.84658, 55.83772, 55.82857, 55.81913, 55.8094, 55.79939, 55.78909, 
    55.7785, 55.76764, 55.75648, 55.74503, 55.73331, 55.72129, 55.709, 
    55.69642, 55.68356, 55.67041, 55.65697, 55.64326, 55.62926, 55.61499, 
    55.60043, 55.58559, 55.57046, 55.55506, 55.53938, 55.52341, 55.50717, 
    55.49065, 55.47385, 55.45677, 55.43941, 55.42178, 55.40387, 55.38568, 
    55.36722, 55.34848, 55.32947, 55.31018, 55.29062, 55.27078, 55.25067, 
    55.23029, 55.20963, 55.18871, 55.16751, 55.14604, 55.1243, 55.10229, 
    55.08001, 55.05747, 55.03465, 55.01157, 54.98822, 54.96461, 54.94073, 
    54.91658, 54.89217, 54.86749, 54.84255, 54.81735, 54.79188, 54.76616, 
    54.74017, 54.71392, 54.68741, 54.66064, 54.63361, 54.60632, 54.57878, 
    54.55098, 54.52292, 54.49461, 54.46604, 54.43721, 54.40813, 54.3788, 
    54.34922, 54.31938, 54.2893, 54.25896, 54.22837, 54.19753, 54.16645, 
    54.13511, 54.10353, 54.0717, 54.03963, 54.00731, 53.97474, 53.94193, 
    53.90888, 53.87558, 53.84204, 53.80827, 53.77425, 53.73999, 53.70549, 
    53.67075, 53.63578, 53.60057, 53.56512, 53.52944, 53.49352, 53.45737, 
    53.42098, 53.38436, 53.34751, 53.31043, 53.27311, 53.23557, 53.1978, 
    53.1598, 53.12157, 53.08311, 53.04443, 53.00552, 52.96639, 52.92704, 
    52.88745, 52.84765, 52.80763, 52.76738, 52.72692, 52.68623, 52.64533, 
    52.60421, 52.56287, 52.52131, 52.47954, 52.43755, 52.39535, 52.35294, 
    52.31031, 52.26747, 52.22441, 52.18115, 52.13768, 52.094, 52.05011, 
    52.00601, 51.9617,
  47.14006, 47.2005, 47.2608, 47.32095, 47.38097, 47.44084, 47.50056, 
    47.56015, 47.61959, 47.67888, 47.73803, 47.79702, 47.85588, 47.91458, 
    47.97313, 48.03154, 48.08979, 48.1479, 48.20585, 48.26365, 48.3213, 
    48.37879, 48.43613, 48.49332, 48.55035, 48.60722, 48.66394, 48.7205, 
    48.7769, 48.83314, 48.88922, 48.94514, 49.0009, 49.0565, 49.11193, 
    49.16721, 49.22232, 49.27726, 49.33204, 49.38665, 49.4411, 49.49538, 
    49.54949, 49.60343, 49.65721, 49.71081, 49.76424, 49.8175, 49.87059, 
    49.9235, 49.97625, 50.02881, 50.0812, 50.13342, 50.18546, 50.23732, 
    50.289, 50.3405, 50.39183, 50.44297, 50.49393, 50.54472, 50.59531, 
    50.64573, 50.69596, 50.74601, 50.79587, 50.84554, 50.89503, 50.94433, 
    50.99344, 51.04237, 51.0911, 51.13964, 51.18799, 51.23615, 51.28411, 
    51.33189, 51.37946, 51.42685, 51.47403, 51.52102, 51.56781, 51.61441, 
    51.6608, 51.70699, 51.75299, 51.79878, 51.84438, 51.88976, 51.93495, 
    51.97993, 52.0247, 52.06927, 52.11364, 52.15779, 52.20174, 52.24548, 
    52.28902, 52.33234, 52.37545, 52.41834, 52.46103, 52.5035, 52.54576, 
    52.5878, 52.62963, 52.67124, 52.71263, 52.75381, 52.79477, 52.83551, 
    52.87602, 52.91632, 52.9564, 52.99625, 53.03588, 53.07529, 53.11448, 
    53.15343, 53.19217, 53.23067, 53.26895, 53.307, 53.34482, 53.38241, 
    53.41977, 53.4569, 53.4938, 53.53046, 53.56689, 53.60309, 53.63905, 
    53.67478, 53.71027, 53.74553, 53.78055, 53.81533, 53.84986, 53.88417, 
    53.91822, 53.95205, 53.98562, 54.01896, 54.05205, 54.0849, 54.1175, 
    54.14986, 54.18197, 54.21383, 54.24545, 54.27682, 54.30794, 54.33881, 
    54.36943, 54.39981, 54.42992, 54.45979, 54.48941, 54.51877, 54.54788, 
    54.57673, 54.60533, 54.63367, 54.66176, 54.68959, 54.71716, 54.74447, 
    54.77152, 54.79832, 54.82485, 54.85112, 54.87714, 54.90289, 54.92837, 
    54.95359, 54.97856, 55.00325, 55.02768, 55.05185, 55.07575, 55.09938, 
    55.12275, 55.14584, 55.16867, 55.19123, 55.21352, 55.23555, 55.2573, 
    55.27877, 55.29998, 55.32092, 55.34159, 55.36198, 55.3821, 55.40194, 
    55.42151, 55.4408, 55.45982, 55.47857, 55.49703, 55.51522, 55.53313, 
    55.55077, 55.56813, 55.58521, 55.60201, 55.61852, 55.63477, 55.65073, 
    55.6664, 55.6818, 55.69692, 55.71176, 55.72631, 55.74058, 55.75457, 
    55.76827, 55.7817, 55.79483, 55.80769, 55.82026, 55.83254, 55.84454, 
    55.85625, 55.86768, 55.87882, 55.88967, 55.90024, 55.91052, 55.92052, 
    55.93022, 55.93964, 55.94877, 55.95761, 55.96617, 55.97443, 55.98241, 
    55.9901, 55.99749, 56.0046, 56.01143, 56.01795, 56.02419, 56.03014, 
    56.0358, 56.04117, 56.04625, 56.05103, 56.05553, 56.05973, 56.06365, 
    56.06727, 56.0706, 56.07364, 56.07639, 56.07885, 56.08101, 56.08289, 
    56.08447, 56.08576, 56.08675, 56.08746, 56.08788, 56.088, 56.08783, 
    56.08737, 56.08662, 56.08557, 56.08424, 56.08261, 56.08069, 56.07848, 
    56.07597, 56.07318, 56.07009, 56.06672, 56.06305, 56.05909, 56.05484, 
    56.05029, 56.04546, 56.04034, 56.03492, 56.02922, 56.02322, 56.01694, 
    56.01036, 56.0035, 55.99635, 55.9889, 55.98117, 55.97314, 55.96483, 
    55.95623, 55.94735, 55.93817, 55.92871, 55.91895, 55.90892, 55.89859, 
    55.88797, 55.87708, 55.86589, 55.85442, 55.84266, 55.83062, 55.81829, 
    55.80567, 55.79277, 55.77959, 55.76612, 55.75238, 55.73834, 55.72403, 
    55.70943, 55.69455, 55.67939, 55.66394, 55.64822, 55.63221, 55.61593, 
    55.59937, 55.58252, 55.5654, 55.548, 55.53032, 55.51236, 55.49413, 
    55.47562, 55.45683, 55.43777, 55.41843, 55.39882, 55.37893, 55.35877, 
    55.33833, 55.31763, 55.29665, 55.2754, 55.25387, 55.23208, 55.21001, 
    55.18768, 55.16508, 55.14221, 55.11907, 55.09566, 55.07198, 55.04804, 
    55.02383, 54.99936, 54.97462, 54.94962, 54.92436, 54.89883, 54.87304, 
    54.84698, 54.82067, 54.7941, 54.76726, 54.74017, 54.71281, 54.6852, 
    54.65733, 54.6292, 54.60082, 54.57219, 54.54329, 54.51414, 54.48474, 
    54.45509, 54.42518, 54.39502, 54.36461, 54.33395, 54.30304, 54.27187, 
    54.24047, 54.20881, 54.1769, 54.14475, 54.11236, 54.07972, 54.04683, 
    54.0137, 53.98033, 53.94671, 53.91285, 53.87876, 53.84442, 53.80984, 
    53.77502, 53.73997, 53.70468, 53.66915, 53.63338, 53.59738, 53.56115, 
    53.52468, 53.48798, 53.45104, 53.41388, 53.37648, 53.33885, 53.30099, 
    53.26291, 53.22459, 53.18605, 53.14729, 53.10829, 53.06907, 53.02963, 
    52.98996, 52.95007, 52.90996, 52.86963, 52.82907, 52.7883, 52.74731, 
    52.7061, 52.66467, 52.62302, 52.58117, 52.53909, 52.4968, 52.45429, 
    52.41157, 52.36864, 52.3255, 52.28214, 52.23858, 52.19481, 52.15083, 
    52.10664, 52.06224,
  47.23171, 47.29224, 47.35263, 47.41289, 47.473, 47.53296, 47.59278, 
    47.65246, 47.71199, 47.77138, 47.83062, 47.88971, 47.94866, 48.00746, 
    48.06611, 48.12461, 48.18296, 48.24116, 48.29921, 48.3571, 48.41484, 
    48.47243, 48.52987, 48.58715, 48.64427, 48.70124, 48.75805, 48.81471, 
    48.8712, 48.92754, 48.98372, 49.03974, 49.09559, 49.15129, 49.20682, 
    49.26219, 49.31739, 49.37244, 49.42731, 49.48202, 49.53656, 49.59094, 
    49.64515, 49.69918, 49.75305, 49.80675, 49.86028, 49.91364, 49.96682, 
    50.01983, 50.07267, 50.12533, 50.17782, 50.23013, 50.28226, 50.33422, 
    50.386, 50.4376, 50.48902, 50.54026, 50.59132, 50.6422, 50.69289, 
    50.7434, 50.79373, 50.84387, 50.89383, 50.9436, 50.99318, 51.04258, 
    51.09179, 51.1408, 51.18963, 51.23827, 51.28671, 51.33496, 51.38303, 
    51.43089, 51.47857, 51.52604, 51.57332, 51.6204, 51.66729, 51.71398, 
    51.76046, 51.80676, 51.85284, 51.89873, 51.94441, 51.98989, 52.03518, 
    52.08025, 52.12511, 52.16978, 52.21423, 52.25848, 52.30252, 52.34636, 
    52.38998, 52.43339, 52.47659, 52.51958, 52.56236, 52.60492, 52.64726, 
    52.6894, 52.73132, 52.77301, 52.8145, 52.85576, 52.89681, 52.93764, 
    52.97824, 53.01863, 53.0588, 53.09874, 53.13845, 53.17795, 53.21722, 
    53.25626, 53.29508, 53.33367, 53.37204, 53.41017, 53.44807, 53.48575, 
    53.5232, 53.56041, 53.59739, 53.63414, 53.67065, 53.70694, 53.74298, 
    53.77879, 53.81437, 53.8497, 53.8848, 53.91966, 53.95428, 53.98866, 
    54.0228, 54.05669, 54.09035, 54.12376, 54.15693, 54.18986, 54.22254, 
    54.25497, 54.28716, 54.3191, 54.35079, 54.38224, 54.41343, 54.44438, 
    54.47507, 54.50552, 54.53571, 54.56565, 54.59534, 54.62477, 54.65395, 
    54.68287, 54.71154, 54.73995, 54.7681, 54.796, 54.82364, 54.85102, 
    54.87814, 54.905, 54.9316, 54.95794, 54.98401, 55.00983, 55.03538, 
    55.06066, 55.08569, 55.11044, 55.13493, 55.15916, 55.18312, 55.20681, 
    55.23024, 55.25339, 55.27628, 55.2989, 55.32124, 55.34332, 55.36513, 
    55.38666, 55.40792, 55.42891, 55.44963, 55.47007, 55.49024, 55.51014, 
    55.52976, 55.5491, 55.56817, 55.58696, 55.60548, 55.62371, 55.64167, 
    55.65935, 55.67675, 55.69388, 55.71072, 55.72728, 55.74357, 55.75957, 
    55.77529, 55.79073, 55.80589, 55.82076, 55.83535, 55.84966, 55.86369, 
    55.87743, 55.89088, 55.90405, 55.91694, 55.92954, 55.94186, 55.95389, 
    55.96563, 55.97709, 55.98826, 55.99915, 56.00974, 56.02005, 56.03007, 
    56.0398, 56.04924, 56.0584, 56.06726, 56.07584, 56.08413, 56.09213, 
    56.09983, 56.10725, 56.11438, 56.12122, 56.12777, 56.13402, 56.13998, 
    56.14566, 56.15104, 56.15613, 56.16093, 56.16544, 56.16966, 56.17358, 
    56.17721, 56.18055, 56.1836, 56.18636, 56.18882, 56.19099, 56.19287, 
    56.19446, 56.19575, 56.19675, 56.19746, 56.19788, 56.198, 56.19783, 
    56.19737, 56.19661, 56.19556, 56.19423, 56.19259, 56.19067, 56.18845, 
    56.18594, 56.18314, 56.18005, 56.17666, 56.17298, 56.16901, 56.16475, 
    56.16019, 56.15535, 56.15021, 56.14478, 56.13906, 56.13305, 56.12675, 
    56.12016, 56.11327, 56.1061, 56.09864, 56.09088, 56.08284, 56.0745, 
    56.06588, 56.05697, 56.04777, 56.03828, 56.0285, 56.01844, 56.00808, 
    55.99744, 55.98651, 55.9753, 55.96379, 55.952, 55.93993, 55.92757, 
    55.91492, 55.90199, 55.88877, 55.87527, 55.86148, 55.84742, 55.83306, 
    55.81842, 55.8035, 55.7883, 55.77282, 55.75706, 55.74101, 55.72468, 
    55.70808, 55.69119, 55.67402, 55.65657, 55.63885, 55.62085, 55.60257, 
    55.58401, 55.56517, 55.54606, 55.52667, 55.50701, 55.48707, 55.46686, 
    55.44637, 55.42561, 55.40458, 55.38327, 55.36169, 55.33985, 55.31773, 
    55.29534, 55.27267, 55.24974, 55.22655, 55.20308, 55.17935, 55.15535, 
    55.13108, 55.10654, 55.08175, 55.05668, 55.03135, 55.00576, 54.9799, 
    54.95379, 54.92741, 54.90077, 54.87387, 54.84671, 54.81928, 54.7916, 
    54.76367, 54.73547, 54.70702, 54.67831, 54.64935, 54.62013, 54.59066, 
    54.56093, 54.53095, 54.50072, 54.47023, 54.4395, 54.40851, 54.37728, 
    54.34579, 54.31406, 54.28208, 54.24986, 54.21738, 54.18467, 54.1517, 
    54.1185, 54.08504, 54.05135, 54.01741, 53.98323, 53.94882, 53.91416, 
    53.87926, 53.84413, 53.80875, 53.77314, 53.73729, 53.70121, 53.66489, 
    53.62834, 53.59156, 53.55454, 53.51729, 53.4798, 53.44209, 53.40415, 
    53.36598, 53.32758, 53.28896, 53.2501, 53.21102, 53.17171, 53.13219, 
    53.09243, 53.05246, 53.01226, 52.97184, 52.93119, 52.89033, 52.84925, 
    52.80795, 52.76643, 52.7247, 52.68275, 52.64058, 52.5982, 52.5556, 
    52.51279, 52.46977, 52.42654, 52.38309, 52.33944, 52.29557, 52.2515, 
    52.20722, 52.16273,
  47.3233, 47.38392, 47.4444, 47.50475, 47.56495, 47.62501, 47.68493, 
    47.7447, 47.80433, 47.86381, 47.92315, 47.98233, 48.04137, 48.10027, 
    48.15901, 48.21761, 48.27605, 48.33435, 48.39249, 48.45048, 48.50832, 
    48.56601, 48.62354, 48.68091, 48.73814, 48.7952, 48.85211, 48.90886, 
    48.96545, 49.02188, 49.07816, 49.13427, 49.19022, 49.24601, 49.30164, 
    49.35711, 49.41241, 49.46755, 49.52252, 49.57732, 49.63197, 49.68644, 
    49.74074, 49.79488, 49.84884, 49.90264, 49.95626, 50.00971, 50.063, 
    50.1161, 50.16904, 50.22179, 50.27438, 50.32679, 50.37902, 50.43107, 
    50.48294, 50.53464, 50.58616, 50.6375, 50.68865, 50.73962, 50.79041, 
    50.84102, 50.89145, 50.94168, 50.99174, 51.0416, 51.09128, 51.14077, 
    51.19007, 51.23919, 51.28811, 51.33684, 51.38538, 51.43373, 51.48189, 
    51.52985, 51.57761, 51.62519, 51.67256, 51.71974, 51.76672, 51.8135, 
    51.86008, 51.90647, 51.95265, 51.99863, 52.04441, 52.08998, 52.13535, 
    52.18052, 52.22548, 52.27024, 52.31479, 52.35913, 52.40326, 52.44718, 
    52.4909, 52.5344, 52.57769, 52.62077, 52.66364, 52.70629, 52.74873, 
    52.79095, 52.83296, 52.87475, 52.91632, 52.95768, 52.99881, 53.03973, 
    53.08043, 53.1209, 53.16115, 53.20118, 53.24099, 53.28057, 53.31993, 
    53.35906, 53.39796, 53.43664, 53.47509, 53.51331, 53.5513, 53.58906, 
    53.62659, 53.66389, 53.70095, 53.73779, 53.77438, 53.81075, 53.84687, 
    53.88277, 53.91842, 53.95384, 53.98902, 54.02396, 54.05866, 54.09312, 
    54.12734, 54.16132, 54.19505, 54.22854, 54.26179, 54.29479, 54.32755, 
    54.36006, 54.39233, 54.42434, 54.45611, 54.48763, 54.5189, 54.54992, 
    54.58069, 54.61121, 54.64147, 54.67148, 54.70124, 54.73074, 54.75999, 
    54.78899, 54.81773, 54.84621, 54.87443, 54.9024, 54.9301, 54.95755, 
    54.98474, 55.01166, 55.03833, 55.06473, 55.09087, 55.11675, 55.14236, 
    55.16771, 55.1928, 55.21762, 55.24217, 55.26646, 55.29048, 55.31423, 
    55.33771, 55.36093, 55.38387, 55.40655, 55.42895, 55.45108, 55.47295, 
    55.49453, 55.51585, 55.5369, 55.55767, 55.57816, 55.59838, 55.61833, 
    55.638, 55.65739, 55.67651, 55.69535, 55.71391, 55.7322, 55.7502, 
    55.76793, 55.78537, 55.80254, 55.81943, 55.83604, 55.85236, 55.8684, 
    55.88417, 55.89965, 55.91484, 55.92976, 55.94439, 55.95873, 55.97279, 
    55.98657, 56.00006, 56.01327, 56.02619, 56.03883, 56.05117, 56.06324, 
    56.07501, 56.0865, 56.0977, 56.10861, 56.11924, 56.12957, 56.13962, 
    56.14938, 56.15885, 56.16803, 56.17691, 56.18552, 56.19382, 56.20184, 
    56.20957, 56.21701, 56.22416, 56.23101, 56.23758, 56.24385, 56.24983, 
    56.25552, 56.26091, 56.26602, 56.27083, 56.27535, 56.27958, 56.28352, 
    56.28716, 56.29051, 56.29356, 56.29633, 56.2988, 56.30097, 56.30286, 
    56.30445, 56.30574, 56.30675, 56.30746, 56.30788, 56.308, 56.30783, 
    56.30737, 56.30661, 56.30556, 56.30421, 56.30258, 56.30065, 56.29842, 
    56.29591, 56.2931, 56.29, 56.2866, 56.28291, 56.27893, 56.27466, 
    56.27009, 56.26523, 56.26008, 56.25464, 56.2489, 56.24287, 56.23656, 
    56.22995, 56.22305, 56.21585, 56.20837, 56.2006, 56.19253, 56.18417, 
    56.17553, 56.16659, 56.15737, 56.14785, 56.13805, 56.12796, 56.11758, 
    56.10691, 56.09595, 56.0847, 56.07317, 56.06135, 56.04924, 56.03685, 
    56.02417, 56.0112, 55.99795, 55.98441, 55.97059, 55.95648, 55.94209, 
    55.92742, 55.91246, 55.89722, 55.88169, 55.86589, 55.8498, 55.83343, 
    55.81678, 55.79985, 55.78263, 55.76514, 55.74737, 55.72932, 55.71099, 
    55.69239, 55.6735, 55.65434, 55.6349, 55.61519, 55.5952, 55.57494, 
    55.5544, 55.53358, 55.5125, 55.49114, 55.46951, 55.4476, 55.42542, 
    55.40298, 55.38026, 55.35727, 55.33401, 55.31049, 55.28669, 55.26263, 
    55.2383, 55.21371, 55.18885, 55.16372, 55.13833, 55.11267, 55.08675, 
    55.06057, 55.03413, 55.00742, 54.98045, 54.95322, 54.92574, 54.89799, 
    54.86998, 54.84172, 54.8132, 54.78442, 54.75539, 54.72609, 54.69655, 
    54.66675, 54.6367, 54.6064, 54.57584, 54.54503, 54.51397, 54.48266, 
    54.4511, 54.41929, 54.38724, 54.35493, 54.32238, 54.28959, 54.25655, 
    54.22326, 54.18973, 54.15596, 54.12194, 54.08768, 54.05319, 54.01845, 
    53.98347, 53.94825, 53.9128, 53.87711, 53.84118, 53.80501, 53.76861, 
    53.73198, 53.69511, 53.658, 53.62067, 53.5831, 53.54531, 53.50728, 
    53.46902, 53.43054, 53.39182, 53.35288, 53.31372, 53.27432, 53.23471, 
    53.19487, 53.1548, 53.11451, 53.07401, 53.03327, 52.99232, 52.95115, 
    52.90976, 52.86816, 52.82633, 52.78429, 52.74203, 52.69956, 52.65687, 
    52.61397, 52.57086, 52.52753, 52.484, 52.44025, 52.39629, 52.35213, 
    52.30775, 52.26317,
  47.41481, 47.47553, 47.53611, 47.59655, 47.65684, 47.717, 47.77701, 
    47.83687, 47.8966, 47.95617, 48.0156, 48.07489, 48.13402, 48.19301, 
    48.25185, 48.31054, 48.36908, 48.42747, 48.48571, 48.5438, 48.60173, 
    48.65952, 48.71714, 48.77461, 48.83193, 48.88909, 48.94609, 49.00294, 
    49.05963, 49.11616, 49.17253, 49.22874, 49.28479, 49.34068, 49.3964, 
    49.45197, 49.50736, 49.5626, 49.61766, 49.67257, 49.7273, 49.78187, 
    49.83627, 49.8905, 49.94457, 49.99846, 50.05218, 50.10573, 50.15911, 
    50.21231, 50.26534, 50.3182, 50.37088, 50.42339, 50.47571, 50.52786, 
    50.57983, 50.63163, 50.68324, 50.73467, 50.78593, 50.83699, 50.88788, 
    50.93859, 50.98911, 51.03944, 51.08959, 51.13955, 51.18933, 51.23891, 
    51.28831, 51.33752, 51.38654, 51.43537, 51.484, 51.53245, 51.5807, 
    51.62875, 51.67662, 51.72428, 51.77175, 51.81902, 51.8661, 51.91298, 
    51.95965, 52.00613, 52.05241, 52.09848, 52.14435, 52.19002, 52.23549, 
    52.28075, 52.3258, 52.37065, 52.41529, 52.45972, 52.50395, 52.54797, 
    52.59177, 52.63537, 52.67875, 52.72192, 52.76488, 52.80762, 52.85015, 
    52.89247, 52.93457, 52.97645, 53.01811, 53.05956, 53.10078, 53.14178, 
    53.18257, 53.22313, 53.26347, 53.30359, 53.34349, 53.38316, 53.4226, 
    53.46182, 53.50081, 53.53957, 53.57811, 53.61641, 53.65449, 53.69234, 
    53.72995, 53.76733, 53.80449, 53.8414, 53.87808, 53.91453, 53.95074, 
    53.98671, 54.02245, 54.05795, 54.09321, 54.12823, 54.16302, 54.19756, 
    54.23185, 54.26591, 54.29972, 54.33329, 54.36662, 54.3997, 54.43254, 
    54.46512, 54.49746, 54.52956, 54.5614, 54.593, 54.62434, 54.65544, 
    54.68628, 54.71687, 54.74721, 54.77729, 54.80713, 54.8367, 54.86602, 
    54.89508, 54.92389, 54.95245, 54.98074, 55.00877, 55.03654, 55.06406, 
    55.09132, 55.11831, 55.14504, 55.17151, 55.19771, 55.22366, 55.24933, 
    55.27475, 55.2999, 55.32478, 55.34939, 55.37374, 55.39782, 55.42163, 
    55.44518, 55.46845, 55.49145, 55.51418, 55.53664, 55.55883, 55.58075, 
    55.6024, 55.62377, 55.64487, 55.66569, 55.68624, 55.70651, 55.72651, 
    55.74623, 55.76567, 55.78484, 55.80373, 55.82234, 55.84067, 55.85872, 
    55.8765, 55.89399, 55.9112, 55.92813, 55.94478, 55.96115, 55.97723, 
    55.99304, 56.00856, 56.0238, 56.03875, 56.05342, 56.0678, 56.0819, 
    56.09571, 56.10924, 56.12248, 56.13544, 56.14811, 56.16049, 56.17258, 
    56.18439, 56.19591, 56.20713, 56.21808, 56.22873, 56.23909, 56.24917, 
    56.25895, 56.26844, 56.27765, 56.28656, 56.29519, 56.30352, 56.31156, 
    56.31931, 56.32676, 56.33393, 56.34081, 56.34739, 56.35368, 56.35967, 
    56.36538, 56.37079, 56.37591, 56.38073, 56.38527, 56.3895, 56.39345, 
    56.3971, 56.40046, 56.40352, 56.4063, 56.40877, 56.41095, 56.41284, 
    56.41444, 56.41574, 56.41674, 56.41746, 56.41787, 56.418, 56.41783, 
    56.41737, 56.41661, 56.41555, 56.4142, 56.41256, 56.41063, 56.4084, 
    56.40588, 56.40306, 56.39995, 56.39654, 56.39285, 56.38885, 56.38457, 
    56.37999, 56.37512, 56.36995, 56.36449, 56.35875, 56.3527, 56.34636, 
    56.33974, 56.33282, 56.3256, 56.3181, 56.31031, 56.30222, 56.29384, 
    56.28517, 56.27621, 56.26696, 56.25742, 56.24759, 56.23747, 56.22706, 
    56.21637, 56.20538, 56.1941, 56.18254, 56.17069, 56.15855, 56.14612, 
    56.13341, 56.12041, 56.10712, 56.09355, 56.07969, 56.06554, 56.05111, 
    56.0364, 56.0214, 56.00612, 55.99056, 55.97471, 55.95858, 55.94217, 
    55.92547, 55.9085, 55.89124, 55.8737, 55.85588, 55.83779, 55.81941, 
    55.80076, 55.78183, 55.76262, 55.74313, 55.72336, 55.70332, 55.68301, 
    55.66241, 55.64154, 55.62041, 55.59899, 55.5773, 55.55534, 55.53311, 
    55.5106, 55.48783, 55.46478, 55.44147, 55.41788, 55.39403, 55.36991, 
    55.34552, 55.32086, 55.29593, 55.27074, 55.24529, 55.21957, 55.19358, 
    55.16734, 55.14083, 55.11406, 55.08702, 55.05973, 55.03217, 55.00435, 
    54.97628, 54.94794, 54.91935, 54.89051, 54.8614, 54.83204, 54.80242, 
    54.77255, 54.74243, 54.71205, 54.68142, 54.65054, 54.6194, 54.58802, 
    54.55638, 54.5245, 54.49237, 54.45998, 54.42736, 54.39449, 54.36137, 
    54.328, 54.29439, 54.26054, 54.22644, 54.19211, 54.15753, 54.12271, 
    54.08765, 54.05235, 54.01682, 53.98104, 53.94503, 53.90878, 53.8723, 
    53.83558, 53.79862, 53.76144, 53.72402, 53.68637, 53.64848, 53.61037, 
    53.57203, 53.53345, 53.49466, 53.45563, 53.41637, 53.3769, 53.33719, 
    53.29726, 53.25711, 53.21673, 53.17613, 53.13531, 53.09427, 53.05301, 
    53.01154, 52.96984, 52.92792, 52.88579, 52.84344, 52.80088, 52.7581, 
    52.71511, 52.6719, 52.62849, 52.58486, 52.54102, 52.49697, 52.45271, 
    52.40825, 52.36357,
  47.50625, 47.56706, 47.62774, 47.68827, 47.74866, 47.80891, 47.86901, 
    47.92897, 47.98879, 48.04847, 48.10799, 48.16737, 48.2266, 48.28569, 
    48.34462, 48.40341, 48.46204, 48.52053, 48.57887, 48.63705, 48.69508, 
    48.75296, 48.81068, 48.86825, 48.92566, 48.98292, 49.04002, 49.09696, 
    49.15375, 49.21037, 49.26684, 49.32315, 49.37929, 49.43528, 49.4911, 
    49.54676, 49.60225, 49.65758, 49.71275, 49.76775, 49.82258, 49.87725, 
    49.93174, 49.98607, 50.04023, 50.09422, 50.14804, 50.20169, 50.25516, 
    50.30846, 50.36159, 50.41454, 50.46732, 50.51992, 50.57235, 50.6246, 
    50.67666, 50.72855, 50.78027, 50.83179, 50.88314, 50.93431, 50.98529, 
    51.03609, 51.08671, 51.13714, 51.18739, 51.23745, 51.28732, 51.337, 
    51.38649, 51.4358, 51.48491, 51.53384, 51.58257, 51.63111, 51.67945, 
    51.72761, 51.77557, 51.82333, 51.87089, 51.91826, 51.96543, 52.0124, 
    52.05917, 52.10574, 52.15211, 52.19828, 52.24425, 52.29001, 52.33557, 
    52.38093, 52.42607, 52.47102, 52.51575, 52.56028, 52.6046, 52.6487, 
    52.6926, 52.73629, 52.77977, 52.82303, 52.86608, 52.90892, 52.95154, 
    52.99394, 53.03613, 53.0781, 53.11985, 53.16139, 53.20271, 53.2438, 
    53.28468, 53.32533, 53.36576, 53.40596, 53.44595, 53.4857, 53.52523, 
    53.56454, 53.60362, 53.64247, 53.68109, 53.71949, 53.75765, 53.79558, 
    53.83328, 53.87075, 53.90798, 53.94498, 53.98175, 54.01828, 54.05457, 
    54.09063, 54.12645, 54.16203, 54.19738, 54.23248, 54.26734, 54.30196, 
    54.33634, 54.37048, 54.40437, 54.43802, 54.47142, 54.50459, 54.53749, 
    54.57016, 54.60258, 54.63475, 54.66667, 54.69834, 54.72976, 54.76093, 
    54.79185, 54.82251, 54.85292, 54.88308, 54.91299, 54.94263, 54.97203, 
    55.00116, 55.03004, 55.05866, 55.08702, 55.11513, 55.14297, 55.17055, 
    55.19788, 55.22493, 55.25173, 55.27827, 55.30454, 55.33055, 55.35629, 
    55.38176, 55.40697, 55.43192, 55.4566, 55.48101, 55.50515, 55.52902, 
    55.55262, 55.57595, 55.59902, 55.62181, 55.64433, 55.66657, 55.68855, 
    55.71025, 55.73167, 55.75282, 55.7737, 55.7943, 55.81463, 55.83467, 
    55.85445, 55.87394, 55.89316, 55.9121, 55.93076, 55.94913, 55.96724, 
    55.98505, 56.00259, 56.01985, 56.03683, 56.05352, 56.06993, 56.08606, 
    56.1019, 56.11747, 56.13274, 56.14773, 56.16244, 56.17686, 56.191, 
    56.20485, 56.21841, 56.23169, 56.24468, 56.25738, 56.26979, 56.28192, 
    56.29376, 56.30531, 56.31657, 56.32754, 56.33822, 56.34861, 56.35871, 
    56.36852, 56.37804, 56.38727, 56.39621, 56.40485, 56.41321, 56.42127, 
    56.42904, 56.43652, 56.4437, 56.4506, 56.4572, 56.4635, 56.46952, 
    56.47523, 56.48066, 56.48579, 56.49063, 56.49518, 56.49943, 56.50338, 
    56.50705, 56.51041, 56.51348, 56.51626, 56.51875, 56.52094, 56.52283, 
    56.52443, 56.52573, 56.52674, 56.52745, 56.52787, 56.528, 56.52783, 
    56.52736, 56.5266, 56.52555, 56.5242, 56.52255, 56.52061, 56.51837, 
    56.51584, 56.51302, 56.5099, 56.50648, 56.50278, 56.49878, 56.49448, 
    56.48989, 56.485, 56.47982, 56.47435, 56.46858, 56.46252, 56.45617, 
    56.44952, 56.44258, 56.43536, 56.42783, 56.42001, 56.41191, 56.40351, 
    56.39481, 56.38583, 56.37656, 56.36699, 56.35713, 56.34699, 56.33655, 
    56.32582, 56.31481, 56.3035, 56.2919, 56.28002, 56.26785, 56.25539, 
    56.24264, 56.22961, 56.21629, 56.20267, 56.18878, 56.1746, 56.16013, 
    56.14538, 56.13034, 56.11502, 56.09941, 56.08353, 56.06735, 56.0509, 
    56.03416, 56.01714, 55.99984, 55.98225, 55.96439, 55.94625, 55.92782, 
    55.90912, 55.89014, 55.87088, 55.85134, 55.83152, 55.81143, 55.79106, 
    55.77042, 55.7495, 55.7283, 55.70683, 55.68509, 55.66307, 55.64078, 
    55.61822, 55.59539, 55.57228, 55.54891, 55.52526, 55.50135, 55.47717, 
    55.45271, 55.42799, 55.40301, 55.37775, 55.35223, 55.32645, 55.3004, 
    55.27409, 55.24751, 55.22067, 55.19357, 55.16621, 55.13858, 55.1107, 
    55.08255, 55.05415, 55.02549, 54.99657, 54.9674, 54.93796, 54.90827, 
    54.87833, 54.84813, 54.81768, 54.78698, 54.75602, 54.72481, 54.69335, 
    54.66164, 54.62968, 54.59747, 54.56501, 54.53231, 54.49936, 54.46616, 
    54.43271, 54.39902, 54.36509, 54.33092, 54.2965, 54.26184, 54.22694, 
    54.1918, 54.15642, 54.1208, 54.08494, 54.04885, 54.01252, 53.97595, 
    53.93914, 53.90211, 53.86483, 53.82733, 53.78959, 53.75163, 53.71343, 
    53.675, 53.63634, 53.59745, 53.55834, 53.519, 53.47943, 53.43964, 
    53.39962, 53.35938, 53.31891, 53.27822, 53.23732, 53.19619, 53.15483, 
    53.11327, 53.07148, 53.02947, 52.98725, 52.94481, 52.90215, 52.85928, 
    52.8162, 52.7729, 52.72939, 52.68567, 52.64174, 52.5976, 52.55325, 
    52.50869, 52.46392,
  47.59762, 47.65853, 47.7193, 47.77992, 47.84041, 47.90075, 47.96095, 
    48.02101, 48.08092, 48.14069, 48.20031, 48.25978, 48.31911, 48.37829, 
    48.43732, 48.4962, 48.55494, 48.61352, 48.67195, 48.73023, 48.78836, 
    48.84633, 48.90415, 48.96181, 49.01932, 49.07668, 49.13387, 49.19091, 
    49.2478, 49.30452, 49.36108, 49.41748, 49.47373, 49.52981, 49.58573, 
    49.64148, 49.69708, 49.75251, 49.80777, 49.86287, 49.91779, 49.97256, 
    50.02715, 50.08158, 50.13584, 50.18992, 50.24384, 50.29758, 50.35115, 
    50.40455, 50.45778, 50.51083, 50.56371, 50.6164, 50.66893, 50.72127, 
    50.77344, 50.82542, 50.87723, 50.92886, 50.9803, 51.03157, 51.08265, 
    51.13354, 51.18426, 51.23479, 51.28513, 51.33529, 51.38525, 51.43503, 
    51.48462, 51.53403, 51.58324, 51.63226, 51.68108, 51.72972, 51.77816, 
    51.82641, 51.87446, 51.92232, 51.96998, 52.01744, 52.06471, 52.11178, 
    52.15865, 52.20531, 52.25178, 52.29804, 52.3441, 52.38996, 52.43561, 
    52.48106, 52.5263, 52.57134, 52.61617, 52.66079, 52.7052, 52.7494, 
    52.79339, 52.83717, 52.88074, 52.9241, 52.96724, 53.01016, 53.05288, 
    53.09537, 53.13765, 53.17971, 53.22156, 53.26318, 53.30459, 53.34578, 
    53.38674, 53.42748, 53.468, 53.5083, 53.54837, 53.58821, 53.62783, 
    53.66722, 53.70639, 53.74533, 53.78404, 53.82252, 53.86077, 53.89878, 
    53.93657, 53.97412, 54.01144, 54.04853, 54.08538, 54.12199, 54.15837, 
    54.19452, 54.23042, 54.26608, 54.30151, 54.33669, 54.37164, 54.40634, 
    54.4408, 54.47502, 54.50899, 54.54272, 54.5762, 54.60944, 54.64243, 
    54.67517, 54.70767, 54.73991, 54.77191, 54.80366, 54.83516, 54.8664, 
    54.89739, 54.92813, 54.95862, 54.98885, 55.01883, 55.04855, 55.07801, 
    55.10722, 55.13617, 55.16486, 55.19329, 55.22146, 55.24937, 55.27703, 
    55.30442, 55.33154, 55.35841, 55.38501, 55.41135, 55.43742, 55.46323, 
    55.48877, 55.51404, 55.53905, 55.56379, 55.58826, 55.61246, 55.63639, 
    55.66006, 55.68345, 55.70657, 55.72942, 55.752, 55.7743, 55.79633, 
    55.81808, 55.83957, 55.86077, 55.8817, 55.90236, 55.92273, 55.94284, 
    55.96266, 55.9822, 56.00147, 56.02046, 56.03917, 56.05759, 56.07574, 
    56.09361, 56.11119, 56.12849, 56.14551, 56.16225, 56.1787, 56.19487, 
    56.21076, 56.22636, 56.24168, 56.25671, 56.27146, 56.28592, 56.30009, 
    56.31398, 56.32758, 56.34089, 56.35392, 56.36665, 56.3791, 56.39126, 
    56.40313, 56.41471, 56.426, 56.437, 56.44771, 56.45813, 56.46825, 
    56.47809, 56.48764, 56.49689, 56.50585, 56.51452, 56.5229, 56.53098, 
    56.53877, 56.54627, 56.55347, 56.56039, 56.56701, 56.57333, 56.57936, 
    56.58509, 56.59053, 56.59568, 56.60053, 56.60509, 56.60935, 56.61332, 
    56.61699, 56.62037, 56.62344, 56.62623, 56.62872, 56.63092, 56.63282, 
    56.63442, 56.63573, 56.63674, 56.63745, 56.63787, 56.638, 56.63783, 
    56.63736, 56.6366, 56.63554, 56.63419, 56.63253, 56.63059, 56.62835, 
    56.62581, 56.62298, 56.61985, 56.61643, 56.61271, 56.6087, 56.60439, 
    56.59978, 56.59488, 56.58969, 56.58421, 56.57842, 56.57235, 56.56598, 
    56.55931, 56.55236, 56.5451, 56.53756, 56.52972, 56.52159, 56.51317, 
    56.50445, 56.49545, 56.48615, 56.47655, 56.46667, 56.4565, 56.44603, 
    56.43528, 56.42423, 56.4129, 56.40127, 56.38935, 56.37715, 56.36466, 
    56.35188, 56.33881, 56.32545, 56.3118, 56.29787, 56.28365, 56.26915, 
    56.25435, 56.23928, 56.22392, 56.20827, 56.19234, 56.17612, 56.15962, 
    56.14284, 56.12577, 56.10843, 56.0908, 56.07289, 56.0547, 56.03622, 
    56.01747, 55.99844, 55.97913, 55.95954, 55.93967, 55.91953, 55.89911, 
    55.87841, 55.85744, 55.83619, 55.81466, 55.79286, 55.77079, 55.74844, 
    55.72582, 55.70293, 55.67977, 55.65633, 55.63263, 55.60865, 55.58441, 
    55.55989, 55.53511, 55.51006, 55.48475, 55.45916, 55.43331, 55.4072, 
    55.38082, 55.35418, 55.32727, 55.3001, 55.27267, 55.24498, 55.21702, 
    55.18881, 55.16034, 55.1316, 55.10262, 55.07337, 55.04386, 55.0141, 
    54.98409, 54.95381, 54.92329, 54.89251, 54.86147, 54.83019, 54.79866, 
    54.76687, 54.73483, 54.70255, 54.67001, 54.63723, 54.6042, 54.57092, 
    54.5374, 54.50363, 54.46962, 54.43536, 54.40086, 54.36612, 54.33114, 
    54.29592, 54.26046, 54.22475, 54.18881, 54.15263, 54.11622, 54.07957, 
    54.04268, 54.00556, 53.9682, 53.93061, 53.89279, 53.85473, 53.81645, 
    53.77793, 53.73919, 53.70021, 53.66101, 53.62158, 53.58192, 53.54204, 
    53.50194, 53.46161, 53.42105, 53.38028, 53.33928, 53.29806, 53.25661, 
    53.21495, 53.17308, 53.13098, 53.08867, 53.04613, 53.00339, 52.96043, 
    52.91725, 52.87386, 52.83026, 52.78645, 52.74242, 52.69818, 52.65374, 
    52.60909, 52.56423,
  47.68892, 47.74992, 47.81078, 47.87151, 47.93209, 47.99252, 48.05282, 
    48.11297, 48.17298, 48.23284, 48.29256, 48.35213, 48.41155, 48.47083, 
    48.52995, 48.58893, 48.64776, 48.70644, 48.76497, 48.82334, 48.88157, 
    48.93964, 48.99755, 49.05531, 49.11292, 49.17037, 49.22766, 49.2848, 
    49.34178, 49.3986, 49.45526, 49.51176, 49.5681, 49.62428, 49.68029, 
    49.73615, 49.79184, 49.84736, 49.90273, 49.95792, 50.01295, 50.06781, 
    50.1225, 50.17702, 50.23138, 50.28556, 50.33958, 50.39342, 50.44709, 
    50.50058, 50.55391, 50.60706, 50.66003, 50.71282, 50.76544, 50.81789, 
    50.87015, 50.92223, 50.97414, 51.02586, 51.07741, 51.12877, 51.17995, 
    51.23094, 51.28175, 51.33237, 51.38282, 51.43307, 51.48314, 51.53301, 
    51.5827, 51.6322, 51.68151, 51.73062, 51.77955, 51.82828, 51.87682, 
    51.92516, 51.97331, 52.02126, 52.06902, 52.11658, 52.16394, 52.21111, 
    52.25806, 52.30483, 52.35139, 52.39775, 52.4439, 52.48986, 52.5356, 
    52.58115, 52.62648, 52.67161, 52.71653, 52.76125, 52.80575, 52.85005, 
    52.89413, 52.93801, 52.98167, 53.02512, 53.06835, 53.11137, 53.15417, 
    53.19676, 53.23914, 53.28129, 53.32322, 53.36494, 53.40644, 53.44771, 
    53.48877, 53.5296, 53.57021, 53.61059, 53.65075, 53.69069, 53.73039, 
    53.76987, 53.80913, 53.84816, 53.88695, 53.92552, 53.96386, 54.00196, 
    54.03983, 54.07747, 54.11488, 54.15205, 54.18898, 54.22568, 54.26214, 
    54.29837, 54.33435, 54.3701, 54.40561, 54.44088, 54.4759, 54.51068, 
    54.54523, 54.57952, 54.61358, 54.64739, 54.68095, 54.71427, 54.74734, 
    54.78016, 54.81273, 54.84505, 54.87713, 54.90895, 54.94053, 54.97185, 
    55.00291, 55.03373, 55.06429, 55.09459, 55.12464, 55.15443, 55.18397, 
    55.21325, 55.24227, 55.27103, 55.29954, 55.32778, 55.35576, 55.38348, 
    55.41094, 55.43813, 55.46507, 55.49173, 55.51814, 55.54427, 55.57014, 
    55.59575, 55.62109, 55.64616, 55.67096, 55.6955, 55.71976, 55.74375, 
    55.76748, 55.79093, 55.81411, 55.83701, 55.85965, 55.88201, 55.9041, 
    55.92591, 55.94744, 55.96871, 55.98969, 56.0104, 56.03083, 56.05098, 
    56.07086, 56.09045, 56.10977, 56.12881, 56.14756, 56.16604, 56.18423, 
    56.20215, 56.21978, 56.23713, 56.25419, 56.27097, 56.28747, 56.30368, 
    56.31961, 56.33526, 56.35062, 56.36569, 56.38047, 56.39497, 56.40918, 
    56.42311, 56.43674, 56.45009, 56.46315, 56.47592, 56.4884, 56.50059, 
    56.51249, 56.52411, 56.53542, 56.54646, 56.55719, 56.56764, 56.57779, 
    56.58766, 56.59723, 56.60651, 56.61549, 56.62418, 56.63258, 56.64069, 
    56.6485, 56.65602, 56.66325, 56.67017, 56.67681, 56.68315, 56.6892, 
    56.69495, 56.70041, 56.70556, 56.71043, 56.715, 56.71927, 56.72325, 
    56.72693, 56.73032, 56.73341, 56.7362, 56.7387, 56.7409, 56.7428, 
    56.74441, 56.74572, 56.74673, 56.74745, 56.74788, 56.748, 56.74783, 
    56.74736, 56.74659, 56.74553, 56.74417, 56.74252, 56.74057, 56.73832, 
    56.73578, 56.73294, 56.7298, 56.72637, 56.72264, 56.71862, 56.71429, 
    56.70968, 56.70477, 56.69956, 56.69406, 56.68826, 56.68217, 56.67578, 
    56.6691, 56.66212, 56.65485, 56.64729, 56.63943, 56.63128, 56.62283, 
    56.61409, 56.60506, 56.59573, 56.58612, 56.57621, 56.56601, 56.55551, 
    56.54473, 56.53365, 56.52229, 56.51063, 56.49868, 56.48645, 56.47392, 
    56.4611, 56.448, 56.4346, 56.42092, 56.40695, 56.3927, 56.37815, 
    56.36332, 56.34821, 56.3328, 56.31711, 56.30114, 56.28488, 56.26834, 
    56.25151, 56.2344, 56.21701, 56.19933, 56.18138, 56.16314, 56.14462, 
    56.12582, 56.10674, 56.08738, 56.06773, 56.04781, 56.02762, 56.00714, 
    55.98639, 55.96536, 55.94406, 55.92248, 55.90062, 55.87849, 55.85609, 
    55.83341, 55.81046, 55.78724, 55.76374, 55.73997, 55.71594, 55.69163, 
    55.66706, 55.64221, 55.6171, 55.59172, 55.56607, 55.54016, 55.51398, 
    55.48753, 55.46082, 55.43385, 55.40661, 55.37911, 55.35135, 55.32333, 
    55.29504, 55.2665, 55.2377, 55.20864, 55.17932, 55.14974, 55.11991, 
    55.08982, 55.05947, 55.02887, 54.99802, 54.96691, 54.93555, 54.90393, 
    54.87207, 54.83996, 54.80759, 54.77498, 54.74212, 54.70901, 54.67566, 
    54.64206, 54.60821, 54.57412, 54.53978, 54.5052, 54.47038, 54.43531, 
    54.40001, 54.36446, 54.32868, 54.29265, 54.25639, 54.21989, 54.18316, 
    54.14618, 54.10897, 54.07153, 54.03386, 53.99594, 53.95781, 53.91943, 
    53.88083, 53.842, 53.80294, 53.76365, 53.72413, 53.68438, 53.64441, 
    53.60422, 53.5638, 53.52315, 53.48228, 53.4412, 53.39989, 53.35836, 
    53.3166, 53.27464, 53.23244, 53.19004, 53.14742, 53.10458, 53.06152, 
    53.01826, 52.97478, 52.93108, 52.88717, 52.84306, 52.79873, 52.75419, 
    52.70944, 52.66449,
  47.78014, 47.84124, 47.9022, 47.96302, 48.02369, 48.08422, 48.14462, 
    48.20486, 48.26497, 48.32492, 48.38474, 48.4444, 48.50392, 48.56329, 
    48.62252, 48.68159, 48.74052, 48.79929, 48.85791, 48.91639, 48.9747, 
    49.03287, 49.09089, 49.14874, 49.20645, 49.264, 49.32138, 49.37862, 
    49.4357, 49.49261, 49.54937, 49.60597, 49.66241, 49.71869, 49.7748, 
    49.83075, 49.88654, 49.94216, 49.99762, 50.05291, 50.10804, 50.16299, 
    50.21778, 50.2724, 50.32686, 50.38114, 50.43525, 50.48919, 50.54296, 
    50.59655, 50.64997, 50.70322, 50.75629, 50.80919, 50.8619, 50.91444, 
    50.9668, 51.01899, 51.07099, 51.12281, 51.17445, 51.22591, 51.27719, 
    51.32828, 51.37919, 51.42991, 51.48045, 51.5308, 51.58096, 51.63093, 
    51.68072, 51.73032, 51.77972, 51.82893, 51.87796, 51.92678, 51.97542, 
    52.02386, 52.07211, 52.12016, 52.16801, 52.21566, 52.26312, 52.31038, 
    52.35744, 52.4043, 52.45095, 52.49741, 52.54366, 52.5897, 52.63555, 
    52.68118, 52.72662, 52.77184, 52.81686, 52.86166, 52.90627, 52.95065, 
    52.99483, 53.0388, 53.08255, 53.12609, 53.16942, 53.21253, 53.25543, 
    53.29811, 53.34057, 53.38282, 53.42485, 53.46665, 53.50824, 53.54961, 
    53.59075, 53.63167, 53.67237, 53.71284, 53.7531, 53.79312, 53.83292, 
    53.87249, 53.91183, 53.95094, 53.98983, 54.02848, 54.06691, 54.10509, 
    54.14305, 54.18078, 54.21827, 54.25553, 54.29255, 54.32933, 54.36588, 
    54.40219, 54.43826, 54.47409, 54.50968, 54.54503, 54.58014, 54.615, 
    54.64963, 54.68401, 54.71814, 54.75203, 54.78567, 54.81907, 54.85221, 
    54.88512, 54.91777, 54.95017, 54.98232, 55.01422, 55.04587, 55.07727, 
    55.10841, 55.1393, 55.16993, 55.20031, 55.23043, 55.2603, 55.28991, 
    55.31926, 55.34835, 55.37719, 55.40576, 55.43407, 55.46213, 55.48991, 
    55.51744, 55.5447, 55.5717, 55.59844, 55.62491, 55.65111, 55.67705, 
    55.70272, 55.72812, 55.75326, 55.77812, 55.80272, 55.82704, 55.8511, 
    55.87488, 55.89839, 55.92163, 55.9446, 55.96729, 55.98971, 56.01185, 
    56.03372, 56.05531, 56.07663, 56.09767, 56.11843, 56.13892, 56.15912, 
    56.17905, 56.1987, 56.21806, 56.23715, 56.25595, 56.27448, 56.29272, 
    56.31068, 56.32836, 56.34575, 56.36287, 56.37969, 56.39623, 56.41249, 
    56.42846, 56.44415, 56.45954, 56.47466, 56.48948, 56.50402, 56.51826, 
    56.53223, 56.5459, 56.55928, 56.57238, 56.58518, 56.5977, 56.60992, 
    56.62185, 56.6335, 56.64485, 56.65591, 56.66668, 56.67715, 56.68733, 
    56.69722, 56.70682, 56.71612, 56.72513, 56.73385, 56.74227, 56.7504, 
    56.75823, 56.76577, 56.77301, 56.77996, 56.78662, 56.79297, 56.79904, 
    56.8048, 56.81027, 56.81545, 56.82033, 56.82491, 56.82919, 56.83318, 
    56.83687, 56.84027, 56.84336, 56.84617, 56.84867, 56.85088, 56.85279, 
    56.8544, 56.85571, 56.85673, 56.85745, 56.85787, 56.858, 56.85783, 
    56.85736, 56.85659, 56.85553, 56.85416, 56.8525, 56.85055, 56.84829, 
    56.84575, 56.8429, 56.83975, 56.83631, 56.83257, 56.82853, 56.8242, 
    56.81957, 56.81465, 56.80943, 56.80391, 56.7981, 56.79199, 56.78558, 
    56.77888, 56.77189, 56.7646, 56.75701, 56.74913, 56.74096, 56.73249, 
    56.72373, 56.71467, 56.70532, 56.69568, 56.68574, 56.67551, 56.66499, 
    56.65417, 56.64307, 56.63168, 56.61999, 56.60801, 56.59574, 56.58318, 
    56.57032, 56.55719, 56.54376, 56.53004, 56.51603, 56.50174, 56.48715, 
    56.47228, 56.45713, 56.44168, 56.42595, 56.40993, 56.39363, 56.37705, 
    56.36018, 56.34302, 56.32558, 56.30786, 56.28986, 56.27157, 56.253, 
    56.23415, 56.21502, 56.19561, 56.17591, 56.15594, 56.1357, 56.11517, 
    56.09436, 56.07328, 56.05192, 56.03028, 56.00837, 55.98618, 55.96372, 
    55.94098, 55.91798, 55.89469, 55.87114, 55.84731, 55.82321, 55.79884, 
    55.77421, 55.7493, 55.72412, 55.69868, 55.67297, 55.64698, 55.62074, 
    55.59423, 55.56745, 55.54041, 55.5131, 55.48554, 55.45771, 55.42962, 
    55.40126, 55.37265, 55.34377, 55.31464, 55.28524, 55.2556, 55.22569, 
    55.19553, 55.1651, 55.13443, 55.1035, 55.07232, 55.04088, 55.00919, 
    54.97725, 54.94506, 54.91262, 54.87993, 54.84699, 54.8138, 54.78036, 
    54.74669, 54.71276, 54.67858, 54.64417, 54.6095, 54.5746, 54.53945, 
    54.50407, 54.46844, 54.43257, 54.39646, 54.36011, 54.32353, 54.28671, 
    54.24965, 54.21236, 54.17483, 54.13707, 54.09907, 54.06084, 54.02238, 
    53.98369, 53.94477, 53.90562, 53.86625, 53.82664, 53.7868, 53.74675, 
    53.70646, 53.66595, 53.62521, 53.58426, 53.54308, 53.50167, 53.46005, 
    53.41821, 53.37615, 53.33387, 53.29137, 53.24866, 53.20573, 53.16258, 
    53.11922, 53.07565, 53.03186, 52.98786, 52.94365, 52.89922, 52.85459, 
    52.80975, 52.7647,
  47.8713, 47.93249, 47.99354, 48.05445, 48.11523, 48.17585, 48.23634, 
    48.29668, 48.35688, 48.41693, 48.47684, 48.53661, 48.59622, 48.65569, 
    48.71501, 48.77418, 48.8332, 48.89207, 48.95079, 49.00936, 49.06778, 
    49.12604, 49.18415, 49.24211, 49.29991, 49.35755, 49.41504, 49.47237, 
    49.52954, 49.58656, 49.64342, 49.70011, 49.75665, 49.81302, 49.86923, 
    49.92528, 49.98117, 50.03689, 50.09245, 50.14783, 50.20306, 50.25811, 
    50.313, 50.36773, 50.42228, 50.47665, 50.53086, 50.5849, 50.63877, 
    50.69246, 50.74598, 50.79932, 50.85249, 50.90548, 50.9583, 51.01094, 
    51.0634, 51.11568, 51.16778, 51.2197, 51.27144, 51.32299, 51.37437, 
    51.42556, 51.47657, 51.52739, 51.57802, 51.62847, 51.67873, 51.7288, 
    51.77868, 51.82838, 51.87788, 51.92719, 51.97631, 52.02523, 52.07397, 
    52.12251, 52.17085, 52.21899, 52.26694, 52.3147, 52.36225, 52.4096, 
    52.45676, 52.50371, 52.55046, 52.59702, 52.64336, 52.6895, 52.73544, 
    52.78117, 52.8267, 52.87202, 52.91713, 52.96203, 53.00673, 53.05121, 
    53.09548, 53.13954, 53.18339, 53.22702, 53.27045, 53.31365, 53.35664, 
    53.39941, 53.44197, 53.48431, 53.52642, 53.56833, 53.61, 53.65146, 
    53.6927, 53.73371, 53.7745, 53.81506, 53.8554, 53.89552, 53.9354, 
    53.97506, 54.01449, 54.0537, 54.09267, 54.13141, 54.16992, 54.2082, 
    54.24624, 54.28405, 54.32163, 54.35897, 54.39608, 54.43295, 54.46958, 
    54.50597, 54.54213, 54.57804, 54.61372, 54.64915, 54.68434, 54.71929, 
    54.75399, 54.78846, 54.82267, 54.85664, 54.89037, 54.92384, 54.95707, 
    54.99005, 55.02278, 55.05526, 55.08749, 55.11946, 55.15119, 55.18266, 
    55.21388, 55.24485, 55.27555, 55.30601, 55.33621, 55.36615, 55.39583, 
    55.42525, 55.45442, 55.48332, 55.51197, 55.54035, 55.56847, 55.59633, 
    55.62392, 55.65126, 55.67833, 55.70513, 55.73166, 55.75793, 55.78394, 
    55.80967, 55.83514, 55.86034, 55.88527, 55.90992, 55.93431, 55.95843, 
    55.98227, 56.00584, 56.02914, 56.05217, 56.07492, 56.0974, 56.1196, 
    56.14152, 56.16317, 56.18454, 56.20564, 56.22646, 56.24699, 56.26725, 
    56.28723, 56.30693, 56.32635, 56.34548, 56.36434, 56.38291, 56.4012, 
    56.41921, 56.43694, 56.45437, 56.47153, 56.4884, 56.50499, 56.52129, 
    56.5373, 56.55302, 56.56847, 56.58362, 56.59848, 56.61306, 56.62735, 
    56.64134, 56.65505, 56.66847, 56.6816, 56.69444, 56.70699, 56.71925, 
    56.73121, 56.74289, 56.75427, 56.76536, 56.77615, 56.78666, 56.79687, 
    56.80678, 56.81641, 56.82573, 56.83477, 56.84351, 56.85196, 56.8601, 
    56.86796, 56.87552, 56.88278, 56.88975, 56.89642, 56.9028, 56.90887, 
    56.91466, 56.92014, 56.92533, 56.93022, 56.93482, 56.93911, 56.94311, 
    56.94682, 56.95022, 56.95333, 56.95613, 56.95864, 56.96086, 56.96277, 
    56.96439, 56.96571, 56.96673, 56.96745, 56.96787, 56.968, 56.96783, 
    56.96735, 56.96659, 56.96552, 56.96415, 56.96249, 56.96053, 56.95827, 
    56.95571, 56.95285, 56.9497, 56.94625, 56.9425, 56.93845, 56.93411, 
    56.92947, 56.92453, 56.9193, 56.91376, 56.90793, 56.90181, 56.89539, 
    56.88867, 56.88165, 56.87434, 56.86674, 56.85883, 56.85064, 56.84215, 
    56.83336, 56.82428, 56.8149, 56.80523, 56.79527, 56.78502, 56.77446, 
    56.76362, 56.75249, 56.74106, 56.72934, 56.71733, 56.70502, 56.69243, 
    56.67954, 56.66637, 56.6529, 56.63915, 56.6251, 56.61077, 56.59615, 
    56.58124, 56.56604, 56.55056, 56.53478, 56.51873, 56.50238, 56.48575, 
    56.46883, 56.45163, 56.43415, 56.41638, 56.39833, 56.37999, 56.36137, 
    56.34248, 56.32329, 56.30383, 56.28409, 56.26406, 56.24376, 56.22318, 
    56.20232, 56.18118, 56.15977, 56.13807, 56.1161, 56.09386, 56.07134, 
    56.04855, 56.02548, 56.00213, 55.97852, 55.95463, 55.93047, 55.90604, 
    55.88134, 55.85637, 55.83113, 55.80562, 55.77984, 55.7538, 55.72748, 
    55.7009, 55.67406, 55.64695, 55.61958, 55.59194, 55.56404, 55.53588, 
    55.50745, 55.47877, 55.44982, 55.42062, 55.39115, 55.36143, 55.33145, 
    55.30121, 55.27072, 55.23997, 55.20896, 55.1777, 55.14619, 55.11443, 
    55.08241, 55.05014, 55.01762, 54.98485, 54.95183, 54.91856, 54.88505, 
    54.85128, 54.81728, 54.78302, 54.74852, 54.71378, 54.67879, 54.64356, 
    54.60809, 54.57238, 54.53643, 54.50023, 54.4638, 54.42713, 54.39022, 
    54.35308, 54.3157, 54.27809, 54.24024, 54.20216, 54.16385, 54.1253, 
    54.08652, 54.04751, 54.00827, 53.9688, 53.92911, 53.88919, 53.84904, 
    53.80866, 53.76806, 53.72724, 53.68619, 53.64492, 53.60342, 53.56171, 
    53.51978, 53.47762, 53.43525, 53.39266, 53.34985, 53.30683, 53.26359, 
    53.22014, 53.17647, 53.13259, 53.08849, 53.04419, 52.99967, 52.95494, 
    52.91001, 52.86486,
  47.96238, 48.02367, 48.08481, 48.14582, 48.20669, 48.26741, 48.32799, 
    48.38843, 48.44873, 48.50888, 48.56888, 48.62874, 48.68845, 48.74801, 
    48.80743, 48.8667, 48.92582, 48.98478, 49.0436, 49.10227, 49.16078, 
    49.21914, 49.27735, 49.3354, 49.3933, 49.45104, 49.50863, 49.56606, 
    49.62333, 49.68044, 49.7374, 49.79419, 49.85082, 49.9073, 49.9636, 
    50.01975, 50.07573, 50.13155, 50.18721, 50.24269, 50.29802, 50.35317, 
    50.40816, 50.46298, 50.51763, 50.57211, 50.62642, 50.68055, 50.73452, 
    50.78831, 50.84192, 50.89537, 50.94863, 51.00172, 51.05464, 51.10738, 
    51.15993, 51.21231, 51.26451, 51.31653, 51.36837, 51.42002, 51.4715, 
    51.52279, 51.57389, 51.62481, 51.67554, 51.72609, 51.77644, 51.82661, 
    51.87659, 51.92638, 51.97598, 52.02539, 52.07461, 52.12363, 52.17246, 
    52.2211, 52.26954, 52.31778, 52.36583, 52.41368, 52.46133, 52.50878, 
    52.55603, 52.60308, 52.64993, 52.69657, 52.74302, 52.78925, 52.83529, 
    52.88111, 52.92674, 52.97215, 53.01736, 53.06236, 53.10714, 53.15172, 
    53.19609, 53.24024, 53.28418, 53.32791, 53.37143, 53.41473, 53.45781, 
    53.50068, 53.54332, 53.58575, 53.62796, 53.66996, 53.71173, 53.75327, 
    53.7946, 53.8357, 53.87658, 53.91724, 53.95767, 53.99787, 54.03785, 
    54.0776, 54.11712, 54.15641, 54.19547, 54.2343, 54.2729, 54.31126, 
    54.3494, 54.38729, 54.42496, 54.46239, 54.49958, 54.53653, 54.57325, 
    54.60973, 54.64597, 54.68197, 54.71773, 54.75324, 54.78852, 54.82355, 
    54.85833, 54.89288, 54.92717, 54.96122, 54.99503, 55.02858, 55.06189, 
    55.09495, 55.12776, 55.16032, 55.19263, 55.22468, 55.25648, 55.28804, 
    55.31933, 55.35037, 55.38116, 55.41168, 55.44196, 55.47197, 55.50172, 
    55.53122, 55.56046, 55.58944, 55.61815, 55.64661, 55.6748, 55.70272, 
    55.73039, 55.75779, 55.78493, 55.8118, 55.8384, 55.86473, 55.8908, 
    55.91661, 55.94214, 55.9674, 55.99239, 56.01711, 56.04156, 56.06574, 
    56.08965, 56.11328, 56.13664, 56.15973, 56.18254, 56.20507, 56.22733, 
    56.24931, 56.27102, 56.29245, 56.31359, 56.33447, 56.35506, 56.37537, 
    56.3954, 56.41515, 56.43462, 56.4538, 56.47271, 56.49133, 56.50967, 
    56.52773, 56.5455, 56.56298, 56.58018, 56.5971, 56.61373, 56.63007, 
    56.64613, 56.6619, 56.67738, 56.69257, 56.70748, 56.72209, 56.73642, 
    56.75045, 56.7642, 56.77766, 56.79082, 56.8037, 56.81628, 56.82857, 
    56.84056, 56.85227, 56.86368, 56.8748, 56.88563, 56.89616, 56.9064, 
    56.91634, 56.92599, 56.93534, 56.9444, 56.95317, 56.96164, 56.96981, 
    56.97768, 56.98526, 56.99255, 56.99953, 57.00623, 57.01262, 57.01871, 
    57.02451, 57.03001, 57.03521, 57.04012, 57.04473, 57.04903, 57.05304, 
    57.05676, 57.06017, 57.06329, 57.0661, 57.06862, 57.07084, 57.07276, 
    57.07438, 57.0757, 57.07673, 57.07745, 57.07787, 57.078, 57.07783, 
    57.07735, 57.07658, 57.07551, 57.07414, 57.07248, 57.07051, 57.06824, 
    57.06568, 57.06281, 57.05965, 57.05619, 57.05243, 57.04837, 57.04402, 
    57.03936, 57.03441, 57.02916, 57.02361, 57.01777, 57.01163, 57.00519, 
    56.99845, 56.99142, 56.98409, 56.97646, 56.96854, 56.96032, 56.9518, 
    56.94299, 56.93388, 56.92448, 56.91479, 56.9048, 56.89451, 56.88393, 
    56.87306, 56.8619, 56.85044, 56.83869, 56.82664, 56.8143, 56.80168, 
    56.78876, 56.77555, 56.76205, 56.74825, 56.73417, 56.7198, 56.70514, 
    56.69019, 56.67495, 56.65942, 56.64361, 56.62751, 56.61112, 56.59444, 
    56.57748, 56.56024, 56.54271, 56.52489, 56.50679, 56.48841, 56.46974, 
    56.45079, 56.43156, 56.41204, 56.39225, 56.37217, 56.35182, 56.33118, 
    56.31027, 56.28907, 56.2676, 56.24585, 56.22383, 56.20152, 56.17895, 
    56.15609, 56.13297, 56.10956, 56.08588, 56.06194, 56.03772, 56.01322, 
    55.98846, 55.96342, 55.93812, 55.91254, 55.8867, 55.86059, 55.83421, 
    55.80756, 55.78065, 55.75348, 55.72603, 55.69833, 55.67036, 55.64212, 
    55.61363, 55.58487, 55.55585, 55.52657, 55.49704, 55.46724, 55.43718, 
    55.40687, 55.3763, 55.34548, 55.3144, 55.28306, 55.25147, 55.21963, 
    55.18753, 55.15519, 55.12259, 55.08974, 55.05664, 55.02329, 54.9897, 
    54.95586, 54.92176, 54.88743, 54.85285, 54.81802, 54.78295, 54.74764, 
    54.71209, 54.67629, 54.64025, 54.60398, 54.56746, 54.5307, 54.49371, 
    54.45648, 54.41902, 54.38132, 54.34338, 54.30521, 54.26681, 54.22817, 
    54.18931, 54.15021, 54.11088, 54.07133, 54.03154, 53.99153, 53.95129, 
    53.91082, 53.87013, 53.82922, 53.78808, 53.74672, 53.70513, 53.66333, 
    53.6213, 53.57906, 53.53659, 53.49391, 53.45101, 53.40789, 53.36456, 
    53.32101, 53.27725, 53.23327, 53.18908, 53.14468, 53.10007, 53.05525, 
    53.01022, 52.96498,
  48.05338, 48.11477, 48.17601, 48.23711, 48.29808, 48.35889, 48.41957, 
    48.48011, 48.5405, 48.60074, 48.66084, 48.7208, 48.78061, 48.84027, 
    48.89978, 48.95914, 49.01836, 49.07743, 49.13634, 49.1951, 49.25372, 
    49.31217, 49.37048, 49.42863, 49.48662, 49.54446, 49.60215, 49.65968, 
    49.71704, 49.77425, 49.83131, 49.8882, 49.94493, 50.0015, 50.05791, 
    50.11415, 50.17023, 50.22615, 50.28191, 50.33749, 50.39291, 50.44817, 
    50.50325, 50.55817, 50.61292, 50.6675, 50.7219, 50.77613, 50.8302, 
    50.88409, 50.93781, 50.99134, 51.04471, 51.0979, 51.15092, 51.20375, 
    51.25641, 51.30889, 51.36118, 51.4133, 51.46524, 51.51699, 51.56856, 
    51.61995, 51.67115, 51.72217, 51.773, 51.82364, 51.8741, 51.92437, 
    51.97445, 52.02433, 52.07404, 52.12354, 52.17286, 52.22198, 52.2709, 
    52.31964, 52.36817, 52.41652, 52.46466, 52.5126, 52.56035, 52.6079, 
    52.65525, 52.70239, 52.74934, 52.79608, 52.84262, 52.88895, 52.93509, 
    52.98101, 53.02673, 53.07224, 53.11754, 53.16263, 53.20752, 53.25219, 
    53.29665, 53.3409, 53.38493, 53.42876, 53.47236, 53.51575, 53.55893, 
    53.60189, 53.64463, 53.68716, 53.72946, 53.77154, 53.8134, 53.85505, 
    53.89647, 53.93766, 53.97863, 54.01938, 54.0599, 54.10019, 54.14026, 
    54.1801, 54.21971, 54.25909, 54.29824, 54.33715, 54.37584, 54.4143, 
    54.45251, 54.4905, 54.52825, 54.56577, 54.60305, 54.64009, 54.67689, 
    54.71345, 54.74977, 54.78586, 54.8217, 54.8573, 54.89266, 54.92777, 
    54.96264, 54.99727, 55.03165, 55.06578, 55.09966, 55.1333, 55.16669, 
    55.19983, 55.23272, 55.26535, 55.29774, 55.32988, 55.36176, 55.39338, 
    55.42475, 55.45587, 55.48673, 55.51733, 55.54768, 55.57777, 55.6076, 
    55.63717, 55.66648, 55.69553, 55.72432, 55.75284, 55.7811, 55.8091, 
    55.83683, 55.8643, 55.89151, 55.91845, 55.94512, 55.97152, 55.99766, 
    56.02352, 56.04912, 56.07445, 56.0995, 56.12429, 56.1488, 56.17304, 
    56.19701, 56.2207, 56.24413, 56.26727, 56.29014, 56.31273, 56.33505, 
    56.35709, 56.37885, 56.40033, 56.42154, 56.44246, 56.46311, 56.48347, 
    56.50356, 56.52336, 56.54288, 56.56212, 56.58107, 56.59975, 56.61813, 
    56.63624, 56.65406, 56.67159, 56.68884, 56.7058, 56.72247, 56.73886, 
    56.75496, 56.77077, 56.78629, 56.80152, 56.81647, 56.83112, 56.84549, 
    56.85956, 56.87334, 56.88684, 56.90004, 56.91294, 56.92556, 56.93789, 
    56.94991, 56.96165, 56.97309, 56.98425, 56.9951, 57.00566, 57.01593, 
    57.0259, 57.03557, 57.04495, 57.05404, 57.06282, 57.07132, 57.07951, 
    57.08741, 57.09501, 57.10231, 57.10932, 57.11603, 57.12244, 57.12855, 
    57.13437, 57.13988, 57.1451, 57.15001, 57.15463, 57.15895, 57.16298, 
    57.1667, 57.17012, 57.17324, 57.17607, 57.17859, 57.18082, 57.18274, 
    57.18437, 57.1857, 57.18672, 57.18745, 57.18787, 57.188, 57.18782, 
    57.18735, 57.18658, 57.1855, 57.18413, 57.18246, 57.18048, 57.17822, 
    57.17564, 57.17277, 57.1696, 57.16613, 57.16236, 57.15829, 57.15392, 
    57.14926, 57.14429, 57.13903, 57.13346, 57.1276, 57.12144, 57.11499, 
    57.10823, 57.10118, 57.09383, 57.08618, 57.07824, 57.06999, 57.06145, 
    57.05262, 57.04349, 57.03406, 57.02434, 57.01432, 57.00401, 56.9934, 
    56.9825, 56.97131, 56.95982, 56.94803, 56.93596, 56.92358, 56.91092, 
    56.89797, 56.88472, 56.87118, 56.85735, 56.84324, 56.82882, 56.81412, 
    56.79913, 56.78385, 56.76828, 56.75243, 56.73628, 56.71985, 56.70313, 
    56.68613, 56.66883, 56.65126, 56.63339, 56.61524, 56.59681, 56.57809, 
    56.55909, 56.53981, 56.52024, 56.5004, 56.48027, 56.45986, 56.43917, 
    56.4182, 56.39695, 56.37543, 56.35362, 56.33154, 56.30918, 56.28654, 
    56.26363, 56.24044, 56.21698, 56.19324, 56.16923, 56.14494, 56.12039, 
    56.09556, 56.07046, 56.04509, 56.01945, 55.99354, 55.96736, 55.94092, 
    55.9142, 55.88722, 55.85998, 55.83247, 55.80469, 55.77665, 55.74834, 
    55.71978, 55.69095, 55.66186, 55.63251, 55.6029, 55.57303, 55.5429, 
    55.51251, 55.48186, 55.45097, 55.41981, 55.38839, 55.35673, 55.32481, 
    55.29263, 55.26021, 55.22753, 55.1946, 55.16143, 55.128, 55.09432, 
    55.0604, 55.02623, 54.99181, 54.95715, 54.92224, 54.88708, 54.85169, 
    54.81605, 54.78017, 54.74405, 54.70768, 54.67108, 54.63424, 54.59716, 
    54.55985, 54.5223, 54.48451, 54.44648, 54.40823, 54.36974, 54.33101, 
    54.29206, 54.25287, 54.21346, 54.17381, 54.13393, 54.09383, 54.0535, 
    54.01295, 53.97216, 53.93116, 53.88993, 53.84847, 53.8068, 53.7649, 
    53.72278, 53.68044, 53.63789, 53.59511, 53.55212, 53.50891, 53.46548, 
    53.42184, 53.37798, 53.33391, 53.28963, 53.24514, 53.20043, 53.15551, 
    53.11039, 53.06505,
  48.14432, 48.2058, 48.26714, 48.32833, 48.38939, 48.45031, 48.51108, 
    48.57171, 48.6322, 48.69254, 48.75274, 48.81279, 48.87269, 48.93245, 
    48.99206, 49.05152, 49.11083, 49.16999, 49.22901, 49.28787, 49.34658, 
    49.40513, 49.46354, 49.52178, 49.57988, 49.63782, 49.6956, 49.75322, 
    49.81069, 49.868, 49.92515, 49.98214, 50.03897, 50.09564, 50.15215, 
    50.20849, 50.26467, 50.32069, 50.37654, 50.43222, 50.48774, 50.54309, 
    50.59828, 50.65329, 50.70814, 50.76282, 50.81733, 50.87166, 50.92582, 
    50.97981, 51.03362, 51.08727, 51.14073, 51.19402, 51.24713, 51.30006, 
    51.35282, 51.4054, 51.45779, 51.51001, 51.56205, 51.6139, 51.66557, 
    51.71706, 51.76836, 51.81947, 51.8704, 51.92114, 51.9717, 52.02207, 
    52.07224, 52.12223, 52.17203, 52.22163, 52.27105, 52.32026, 52.36929, 
    52.41812, 52.46675, 52.51519, 52.56343, 52.61148, 52.65932, 52.70697, 
    52.75441, 52.80166, 52.8487, 52.89554, 52.94218, 52.98861, 53.03483, 
    53.08085, 53.12667, 53.17227, 53.21767, 53.26286, 53.30784, 53.3526, 
    53.39716, 53.44151, 53.48563, 53.52955, 53.57325, 53.61674, 53.66001, 
    53.70306, 53.7459, 53.78852, 53.83091, 53.87309, 53.91504, 53.95678, 
    53.99829, 54.03957, 54.08064, 54.12148, 54.16209, 54.20247, 54.24263, 
    54.28255, 54.32225, 54.36172, 54.40096, 54.43997, 54.47875, 54.51729, 
    54.5556, 54.59367, 54.63151, 54.66911, 54.70648, 54.7436, 54.78049, 
    54.81714, 54.85355, 54.88972, 54.92565, 54.96133, 54.99677, 55.03197, 
    55.06692, 55.10163, 55.13609, 55.1703, 55.20427, 55.23799, 55.27146, 
    55.30468, 55.33765, 55.37036, 55.40283, 55.43504, 55.467, 55.4987, 
    55.53015, 55.56134, 55.59228, 55.62296, 55.65338, 55.68354, 55.71345, 
    55.74309, 55.77248, 55.8016, 55.83046, 55.85905, 55.88739, 55.91545, 
    55.94326, 55.9708, 55.99807, 56.02508, 56.05182, 56.07829, 56.10449, 
    56.13042, 56.15609, 56.18148, 56.2066, 56.23145, 56.25602, 56.28033, 
    56.30436, 56.32811, 56.35159, 56.3748, 56.39773, 56.42038, 56.44275, 
    56.46485, 56.48667, 56.50821, 56.52947, 56.55045, 56.57115, 56.59157, 
    56.61171, 56.63156, 56.65113, 56.67042, 56.68943, 56.70815, 56.72659, 
    56.74474, 56.7626, 56.78018, 56.79747, 56.81448, 56.8312, 56.84763, 
    56.86377, 56.87963, 56.89519, 56.91047, 56.92545, 56.94015, 56.95455, 
    56.96866, 56.98248, 56.99601, 57.00925, 57.02219, 57.03484, 57.0472, 
    57.05926, 57.07103, 57.0825, 57.09369, 57.10457, 57.11516, 57.12545, 
    57.13545, 57.14515, 57.15456, 57.16367, 57.17248, 57.181, 57.18921, 
    57.19713, 57.20475, 57.21208, 57.2191, 57.22583, 57.23226, 57.23838, 
    57.24422, 57.24974, 57.25498, 57.25991, 57.26454, 57.26888, 57.27291, 
    57.27664, 57.28007, 57.2832, 57.28604, 57.28857, 57.2908, 57.29273, 
    57.29436, 57.29569, 57.29672, 57.29744, 57.29787, 57.298, 57.29782, 
    57.29735, 57.29657, 57.2955, 57.29412, 57.29244, 57.29047, 57.28819, 
    57.28561, 57.28273, 57.27955, 57.27607, 57.27229, 57.26821, 57.26383, 
    57.25915, 57.25417, 57.24889, 57.24331, 57.23743, 57.23126, 57.22478, 
    57.21801, 57.21094, 57.20357, 57.1959, 57.18793, 57.17967, 57.1711, 
    57.16225, 57.15309, 57.14364, 57.13389, 57.12384, 57.1135, 57.10287, 
    57.09193, 57.08071, 57.06919, 57.05737, 57.04526, 57.03286, 57.02016, 
    57.00717, 56.99389, 56.98032, 56.96645, 56.95229, 56.93784, 56.9231, 
    56.90807, 56.89275, 56.87714, 56.86124, 56.84505, 56.82858, 56.81181, 
    56.79476, 56.77742, 56.7598, 56.74189, 56.72369, 56.70521, 56.68644, 
    56.66739, 56.64806, 56.62844, 56.60854, 56.58836, 56.56789, 56.54715, 
    56.52613, 56.50482, 56.48324, 56.46137, 56.43923, 56.41681, 56.39412, 
    56.37114, 56.3479, 56.32437, 56.30058, 56.2765, 56.25216, 56.22754, 
    56.20264, 56.17748, 56.15204, 56.12634, 56.10036, 56.07412, 56.04761, 
    56.02082, 55.99378, 55.96646, 55.93888, 55.91103, 55.88292, 55.85455, 
    55.82591, 55.79701, 55.76785, 55.73842, 55.70874, 55.67879, 55.64859, 
    55.61813, 55.5874, 55.55643, 55.52519, 55.49371, 55.46196, 55.42996, 
    55.39771, 55.3652, 55.33245, 55.29944, 55.26618, 55.23267, 55.19891, 
    55.16491, 55.13066, 55.09616, 55.06141, 55.02642, 54.99118, 54.9557, 
    54.91998, 54.88401, 54.84781, 54.81136, 54.77467, 54.73775, 54.70058, 
    54.66318, 54.62554, 54.58767, 54.54955, 54.51121, 54.47263, 54.43382, 
    54.39477, 54.3555, 54.31599, 54.27626, 54.23629, 54.1961, 54.15568, 
    54.11503, 54.07416, 54.03306, 53.99174, 53.95019, 53.90842, 53.86643, 
    53.82422, 53.78179, 53.73914, 53.69627, 53.65318, 53.60988, 53.56636, 
    53.52262, 53.47867, 53.43451, 53.39013, 53.34554, 53.30074, 53.25573, 
    53.2105, 53.16507,
  48.23517, 48.29675, 48.35818, 48.41948, 48.48063, 48.54164, 48.60251, 
    48.66324, 48.72382, 48.78426, 48.84455, 48.9047, 48.96471, 49.02456, 
    49.08427, 49.14383, 49.20324, 49.2625, 49.32161, 49.38056, 49.43937, 
    49.49802, 49.55652, 49.61487, 49.67306, 49.7311, 49.78898, 49.8467, 
    49.90427, 49.96167, 50.01892, 50.07601, 50.13294, 50.18971, 50.24632, 
    50.30276, 50.35904, 50.41515, 50.4711, 50.52689, 50.5825, 50.63796, 
    50.69324, 50.74836, 50.8033, 50.85808, 50.91268, 50.96712, 51.02138, 
    51.07547, 51.12938, 51.18312, 51.23668, 51.29007, 51.34328, 51.39632, 
    51.44917, 51.50185, 51.55435, 51.60666, 51.65879, 51.71075, 51.76252, 
    51.8141, 51.8655, 51.91672, 51.96775, 52.01859, 52.06924, 52.11971, 
    52.16998, 52.22007, 52.26997, 52.31967, 52.36918, 52.4185, 52.46762, 
    52.51655, 52.56528, 52.61382, 52.66216, 52.7103, 52.75824, 52.80599, 
    52.85353, 52.90087, 52.94801, 52.99495, 53.04168, 53.08821, 53.13453, 
    53.18065, 53.22656, 53.27226, 53.31775, 53.36304, 53.40811, 53.45298, 
    53.49763, 53.54206, 53.58629, 53.6303, 53.6741, 53.71768, 53.76105, 
    53.80419, 53.84712, 53.88983, 53.93232, 53.97459, 54.01664, 54.05846, 
    54.10007, 54.14145, 54.1826, 54.22353, 54.26423, 54.30471, 54.34496, 
    54.38498, 54.42477, 54.46432, 54.50365, 54.54275, 54.58162, 54.62025, 
    54.65864, 54.6968, 54.73473, 54.77242, 54.80987, 54.84709, 54.88406, 
    54.9208, 54.95729, 54.99355, 55.02956, 55.06533, 55.10085, 55.13614, 
    55.17117, 55.20596, 55.24051, 55.2748, 55.30885, 55.34265, 55.3762, 
    55.4095, 55.44255, 55.47535, 55.50789, 55.54018, 55.57222, 55.604, 
    55.63552, 55.66679, 55.69781, 55.72856, 55.75906, 55.7893, 55.81927, 
    55.849, 55.87845, 55.90765, 55.93658, 55.96524, 55.99365, 56.02179, 
    56.04967, 56.07727, 56.10462, 56.13169, 56.1585, 56.18504, 56.21131, 
    56.2373, 56.26303, 56.28849, 56.31367, 56.33859, 56.36323, 56.3876, 
    56.41169, 56.4355, 56.45905, 56.48231, 56.5053, 56.52801, 56.55045, 
    56.5726, 56.59447, 56.61607, 56.63739, 56.65842, 56.67918, 56.69965, 
    56.71984, 56.73975, 56.75938, 56.77872, 56.79777, 56.81654, 56.83503, 
    56.85323, 56.87114, 56.88877, 56.90611, 56.92316, 56.93993, 56.9564, 
    56.97258, 56.98848, 57.00409, 57.01941, 57.03443, 57.04916, 57.06361, 
    57.07775, 57.09161, 57.10518, 57.11845, 57.13143, 57.14412, 57.15651, 
    57.1686, 57.1804, 57.19191, 57.20312, 57.21404, 57.22466, 57.23498, 
    57.245, 57.25473, 57.26416, 57.2733, 57.28213, 57.29067, 57.29891, 
    57.30685, 57.3145, 57.32184, 57.32888, 57.33563, 57.34208, 57.34822, 
    57.35406, 57.35961, 57.36486, 57.3698, 57.37445, 57.37879, 57.38284, 
    57.38658, 57.39002, 57.39316, 57.396, 57.39854, 57.40078, 57.40271, 
    57.40435, 57.40568, 57.40672, 57.40744, 57.40787, 57.408, 57.40783, 
    57.40735, 57.40657, 57.40549, 57.40411, 57.40243, 57.40044, 57.39816, 
    57.39557, 57.39268, 57.3895, 57.38601, 57.38222, 57.37812, 57.37373, 
    57.36904, 57.36405, 57.35875, 57.35316, 57.34727, 57.34108, 57.33458, 
    57.32779, 57.3207, 57.3133, 57.30561, 57.29763, 57.28934, 57.28075, 
    57.27187, 57.26269, 57.25321, 57.24343, 57.23336, 57.223, 57.21233, 
    57.20137, 57.19011, 57.17856, 57.16671, 57.15457, 57.14213, 57.1294, 
    57.11637, 57.10305, 57.08944, 57.07554, 57.06134, 57.04685, 57.03207, 
    57.017, 57.00164, 56.98598, 56.97004, 56.95381, 56.93729, 56.92048, 
    56.90339, 56.886, 56.86833, 56.85037, 56.83212, 56.81359, 56.79478, 
    56.77568, 56.75629, 56.73662, 56.71667, 56.69643, 56.67591, 56.65512, 
    56.63404, 56.61267, 56.59103, 56.56911, 56.54692, 56.52444, 56.50168, 
    56.47865, 56.45534, 56.43176, 56.40789, 56.38376, 56.35935, 56.33467, 
    56.30971, 56.28448, 56.25898, 56.23321, 56.20717, 56.18086, 56.15428, 
    56.12743, 56.10031, 56.07293, 56.04527, 56.01736, 55.98917, 55.96073, 
    55.93202, 55.90305, 55.87381, 55.84431, 55.81455, 55.78453, 55.75425, 
    55.72371, 55.69292, 55.66187, 55.63055, 55.59899, 55.56717, 55.53509, 
    55.50276, 55.47017, 55.43734, 55.40425, 55.37091, 55.33732, 55.30348, 
    55.26939, 55.23506, 55.20047, 55.16565, 55.13057, 55.09525, 55.05968, 
    55.02388, 54.98783, 54.95153, 54.915, 54.87823, 54.84122, 54.80396, 
    54.76648, 54.72875, 54.69078, 54.65258, 54.61415, 54.57549, 54.53658, 
    54.49745, 54.45808, 54.41849, 54.37866, 54.3386, 54.29832, 54.25781, 
    54.21707, 54.17611, 54.13492, 54.0935, 54.05186, 54.01, 53.96792, 
    53.92561, 53.88309, 53.84035, 53.79738, 53.7542, 53.7108, 53.66719, 
    53.62336, 53.57931, 53.53505, 53.49058, 53.44589, 53.401, 53.35589, 
    53.31057, 53.26505,
  48.32595, 48.38763, 48.44916, 48.51055, 48.5718, 48.6329, 48.69387, 
    48.7547, 48.81537, 48.87591, 48.9363, 48.99654, 49.05664, 49.1166, 
    49.1764, 49.23606, 49.29556, 49.35492, 49.41413, 49.47319, 49.53209, 
    49.59084, 49.64944, 49.70789, 49.76617, 49.82431, 49.88229, 49.94011, 
    49.99778, 50.05528, 50.11263, 50.16982, 50.22684, 50.28371, 50.34042, 
    50.39696, 50.45333, 50.50955, 50.5656, 50.62148, 50.6772, 50.73275, 
    50.78814, 50.84335, 50.8984, 50.95327, 51.00798, 51.06251, 51.11687, 
    51.17106, 51.22507, 51.27891, 51.33258, 51.38606, 51.43938, 51.49251, 
    51.54546, 51.59824, 51.65084, 51.70325, 51.75549, 51.80754, 51.85941, 
    51.91109, 51.96259, 52.0139, 52.06503, 52.11597, 52.16673, 52.21729, 
    52.26767, 52.31785, 52.36785, 52.41765, 52.46726, 52.51667, 52.5659, 
    52.61493, 52.66376, 52.71239, 52.76083, 52.80907, 52.85711, 52.90495, 
    52.95259, 53.00003, 53.04727, 53.0943, 53.14113, 53.18776, 53.23418, 
    53.28039, 53.3264, 53.3722, 53.41779, 53.46317, 53.50834, 53.5533, 
    53.59805, 53.64258, 53.6869, 53.73101, 53.7749, 53.81858, 53.86203, 
    53.90528, 53.9483, 53.9911, 54.03369, 54.07605, 54.11819, 54.16011, 
    54.20181, 54.24328, 54.28452, 54.32555, 54.36634, 54.40691, 54.44725, 
    54.48736, 54.52724, 54.56689, 54.60631, 54.64549, 54.68445, 54.72317, 
    54.76165, 54.7999, 54.83792, 54.87569, 54.91323, 54.95053, 54.9876, 
    55.02442, 55.061, 55.09734, 55.13344, 55.16929, 55.2049, 55.24027, 
    55.27539, 55.31026, 55.34489, 55.37927, 55.4134, 55.44728, 55.48091, 
    55.51429, 55.54742, 55.5803, 55.61292, 55.64529, 55.67741, 55.70927, 
    55.74087, 55.77222, 55.80331, 55.83414, 55.86471, 55.89503, 55.92508, 
    55.95487, 55.9844, 56.01367, 56.04268, 56.07141, 56.09989, 56.12811, 
    56.15605, 56.18373, 56.21114, 56.23829, 56.26516, 56.29177, 56.3181, 
    56.34417, 56.36996, 56.39549, 56.42074, 56.44572, 56.47042, 56.49485, 
    56.519, 56.54288, 56.56649, 56.58981, 56.61286, 56.63563, 56.65812, 
    56.68034, 56.70227, 56.72393, 56.7453, 56.76639, 56.7872, 56.80772, 
    56.82797, 56.84793, 56.86761, 56.887, 56.90611, 56.92493, 56.94346, 
    56.96171, 56.97968, 56.99735, 57.01473, 57.03183, 57.04864, 57.06516, 
    57.08139, 57.09733, 57.11298, 57.12833, 57.1434, 57.15818, 57.17266, 
    57.18685, 57.20074, 57.21434, 57.22765, 57.24067, 57.25339, 57.26581, 
    57.27794, 57.28978, 57.30131, 57.31255, 57.3235, 57.33415, 57.3445, 
    57.35455, 57.36431, 57.37376, 57.38292, 57.39178, 57.40034, 57.40861, 
    57.41657, 57.42424, 57.4316, 57.43866, 57.44543, 57.45189, 57.45805, 
    57.46392, 57.46948, 57.47474, 57.4797, 57.48436, 57.48871, 57.49277, 
    57.49652, 57.49997, 57.50312, 57.50597, 57.50851, 57.51076, 57.5127, 
    57.51434, 57.51567, 57.51671, 57.51744, 57.51787, 57.518, 57.51782, 
    57.51735, 57.51657, 57.51548, 57.5141, 57.51241, 57.51043, 57.50813, 
    57.50554, 57.50264, 57.49945, 57.49594, 57.49215, 57.48804, 57.48364, 
    57.47893, 57.47393, 57.46862, 57.46301, 57.4571, 57.45089, 57.44438, 
    57.43756, 57.43045, 57.42304, 57.41533, 57.40732, 57.39901, 57.3904, 
    57.38149, 57.37229, 57.36278, 57.35298, 57.34288, 57.33248, 57.32179, 
    57.31079, 57.29951, 57.28792, 57.27604, 57.26387, 57.2514, 57.23863, 
    57.22557, 57.21221, 57.19856, 57.18462, 57.17039, 57.15586, 57.14104, 
    57.12593, 57.11052, 57.09483, 57.07884, 57.06256, 57.046, 57.02915, 
    57.012, 56.99457, 56.97685, 56.95884, 56.94055, 56.92197, 56.9031, 
    56.88395, 56.86451, 56.84479, 56.82479, 56.8045, 56.78392, 56.76307, 
    56.74194, 56.72052, 56.69882, 56.67684, 56.65459, 56.63205, 56.60923, 
    56.58614, 56.56277, 56.53912, 56.5152, 56.491, 56.46653, 56.44178, 
    56.41676, 56.39147, 56.3659, 56.34007, 56.31396, 56.28758, 56.26093, 
    56.23401, 56.20683, 56.17937, 56.15165, 56.12366, 56.09541, 56.06689, 
    56.03811, 56.00906, 55.97975, 55.95018, 55.92034, 55.89025, 55.85989, 
    55.82928, 55.79841, 55.76728, 55.73589, 55.70424, 55.67234, 55.64019, 
    55.60778, 55.57512, 55.5422, 55.50903, 55.47561, 55.44194, 55.40802, 
    55.37384, 55.33943, 55.30476, 55.26985, 55.23469, 55.19929, 55.16364, 
    55.12774, 55.09161, 55.05523, 55.01861, 54.98175, 54.94465, 54.90731, 
    54.86974, 54.83192, 54.79387, 54.75558, 54.71706, 54.6783, 54.63931, 
    54.60009, 54.56063, 54.52095, 54.48103, 54.44088, 54.40051, 54.3599, 
    54.31907, 54.27802, 54.23673, 54.19522, 54.1535, 54.11154, 54.06936, 
    54.02697, 53.98435, 53.94151, 53.89845, 53.85518, 53.81168, 53.76797, 
    53.72404, 53.6799, 53.63555, 53.59098, 53.5462, 53.50121, 53.45601, 
    53.41059, 53.36497,
  48.41666, 48.47843, 48.54005, 48.60154, 48.66289, 48.72409, 48.78516, 
    48.84607, 48.90685, 48.96748, 49.02797, 49.08831, 49.14851, 49.20856, 
    49.26846, 49.32822, 49.38782, 49.44728, 49.50658, 49.56573, 49.62474, 
    49.68359, 49.74229, 49.80083, 49.85922, 49.91745, 49.97553, 50.03345, 
    50.09121, 50.14882, 50.20626, 50.26355, 50.32068, 50.37764, 50.43445, 
    50.49109, 50.54757, 50.60388, 50.66003, 50.71601, 50.77183, 50.82748, 
    50.88297, 50.93828, 50.99343, 51.0484, 51.10321, 51.15784, 51.2123, 
    51.26659, 51.3207, 51.37464, 51.42841, 51.48199, 51.5354, 51.58864, 
    51.64169, 51.69457, 51.74726, 51.79978, 51.85211, 51.90426, 51.95623, 
    52.00801, 52.05962, 52.11103, 52.16226, 52.2133, 52.26415, 52.31482, 
    52.36529, 52.41558, 52.46567, 52.51557, 52.56528, 52.6148, 52.66412, 
    52.71325, 52.76218, 52.81091, 52.85945, 52.90778, 52.95592, 53.00386, 
    53.0516, 53.09914, 53.14647, 53.1936, 53.24053, 53.28725, 53.33377, 
    53.38008, 53.42619, 53.47208, 53.51777, 53.56325, 53.60852, 53.65357, 
    53.69842, 53.74305, 53.78746, 53.83167, 53.87565, 53.91943, 53.96298, 
    54.00632, 54.04943, 54.09233, 54.13501, 54.17747, 54.2197, 54.26171, 
    54.3035, 54.34507, 54.38641, 54.42752, 54.46841, 54.50907, 54.5495, 
    54.5897, 54.62967, 54.66941, 54.70892, 54.7482, 54.78724, 54.82605, 
    54.86462, 54.90297, 54.94107, 54.97893, 55.01656, 55.05395, 55.0911, 
    55.12801, 55.16468, 55.2011, 55.23729, 55.27322, 55.30892, 55.34437, 
    55.37957, 55.41453, 55.44924, 55.4837, 55.51792, 55.55188, 55.58559, 
    55.61906, 55.65226, 55.68522, 55.71793, 55.75038, 55.78257, 55.81451, 
    55.84619, 55.87762, 55.90878, 55.93969, 55.97034, 56.00073, 56.03086, 
    56.06073, 56.09033, 56.11967, 56.14875, 56.17757, 56.20612, 56.2344, 
    56.26242, 56.29016, 56.31765, 56.34486, 56.3718, 56.39848, 56.42488, 
    56.45102, 56.47688, 56.50247, 56.52778, 56.55283, 56.57759, 56.60209, 
    56.6263, 56.65025, 56.67391, 56.6973, 56.72041, 56.74324, 56.76579, 
    56.78806, 56.81005, 56.83176, 56.8532, 56.87434, 56.89521, 56.91579, 
    56.93608, 56.9561, 56.97583, 56.99527, 57.01443, 57.0333, 57.05189, 
    57.07019, 57.0882, 57.10592, 57.12335, 57.1405, 57.15735, 57.17391, 
    57.19019, 57.20617, 57.22186, 57.23726, 57.25237, 57.26718, 57.2817, 
    57.29593, 57.30986, 57.32351, 57.33685, 57.3499, 57.36266, 57.37511, 
    57.38728, 57.39914, 57.41071, 57.42199, 57.43296, 57.44364, 57.45401, 
    57.4641, 57.47388, 57.48336, 57.49255, 57.50143, 57.51002, 57.5183, 
    57.52629, 57.53397, 57.54136, 57.54844, 57.55523, 57.56171, 57.56789, 
    57.57376, 57.57934, 57.58462, 57.58959, 57.59426, 57.59863, 57.6027, 
    57.60646, 57.60992, 57.61308, 57.61594, 57.61849, 57.62074, 57.62268, 
    57.62433, 57.62567, 57.62671, 57.62744, 57.62787, 57.628, 57.62782, 
    57.62735, 57.62656, 57.62548, 57.62409, 57.6224, 57.6204, 57.6181, 
    57.61551, 57.6126, 57.60939, 57.60588, 57.60207, 57.59796, 57.59354, 
    57.58883, 57.5838, 57.57848, 57.57286, 57.56693, 57.5607, 57.55417, 
    57.54734, 57.54021, 57.53278, 57.52504, 57.51701, 57.50868, 57.50005, 
    57.49112, 57.48188, 57.47235, 57.46252, 57.45239, 57.44197, 57.43124, 
    57.42022, 57.4089, 57.39729, 57.38537, 57.37316, 57.36066, 57.34785, 
    57.33476, 57.32137, 57.30768, 57.2937, 57.27943, 57.26486, 57.25, 
    57.23484, 57.2194, 57.20366, 57.18763, 57.17131, 57.1547, 57.1378, 
    57.12061, 57.10313, 57.08537, 57.06731, 57.04897, 57.03034, 57.01142, 
    56.99221, 56.97272, 56.95295, 56.93289, 56.91255, 56.89193, 56.87101, 
    56.84982, 56.82835, 56.80659, 56.78456, 56.76224, 56.73965, 56.71677, 
    56.69362, 56.67019, 56.64648, 56.62249, 56.59823, 56.57369, 56.54888, 
    56.5238, 56.49844, 56.47281, 56.4469, 56.42072, 56.39428, 56.36756, 
    56.34057, 56.31332, 56.28579, 56.258, 56.22994, 56.20162, 56.17303, 
    56.14417, 56.11505, 56.08567, 56.05602, 56.02611, 55.99594, 55.96551, 
    55.93482, 55.90387, 55.87266, 55.8412, 55.80947, 55.7775, 55.74526, 
    55.71277, 55.68003, 55.64703, 55.61378, 55.58028, 55.54652, 55.51252, 
    55.47827, 55.44377, 55.40902, 55.37402, 55.33878, 55.30329, 55.26756, 
    55.23158, 55.19535, 55.15889, 55.12218, 55.08524, 55.04805, 55.01062, 
    54.97296, 54.93505, 54.89692, 54.85854, 54.81993, 54.78108, 54.742, 
    54.70269, 54.66314, 54.62336, 54.58335, 54.54312, 54.50265, 54.46196, 
    54.42103, 54.37988, 54.33851, 54.29691, 54.25508, 54.21304, 54.17076, 
    54.12827, 54.08556, 54.04263, 53.99947, 53.9561, 53.91251, 53.86871, 
    53.82469, 53.78045, 53.736, 53.69134, 53.64646, 53.60137, 53.55607, 
    53.51056, 53.46484,
  48.50729, 48.56915, 48.63088, 48.69246, 48.7539, 48.8152, 48.87636, 
    48.93738, 48.99825, 49.05898, 49.11957, 49.18001, 49.2403, 49.30045, 
    49.36045, 49.4203, 49.48, 49.53956, 49.59896, 49.65821, 49.71732, 
    49.77626, 49.83506, 49.8937, 49.95219, 50.01052, 50.0687, 50.12672, 
    50.18458, 50.24229, 50.29983, 50.35722, 50.41444, 50.47151, 50.52841, 
    50.58515, 50.64173, 50.69814, 50.75439, 50.81048, 50.86639, 50.92215, 
    50.97773, 51.03314, 51.08839, 51.14346, 51.19837, 51.2531, 51.30766, 
    51.36205, 51.41626, 51.4703, 51.52417, 51.57786, 51.63137, 51.6847, 
    51.73786, 51.79083, 51.84363, 51.89624, 51.94868, 52.00093, 52.053, 
    52.10488, 52.15658, 52.2081, 52.25943, 52.31057, 52.36152, 52.41228, 
    52.46286, 52.51324, 52.56343, 52.61344, 52.66325, 52.71286, 52.76228, 
    52.81151, 52.86054, 52.90937, 52.95801, 53.00644, 53.05468, 53.10272, 
    53.15056, 53.19819, 53.24562, 53.29286, 53.33988, 53.3867, 53.43332, 
    53.47973, 53.52593, 53.57192, 53.61771, 53.66328, 53.70864, 53.7538, 
    53.79874, 53.84346, 53.88798, 53.93228, 53.97636, 54.02023, 54.06388, 
    54.10731, 54.15052, 54.19352, 54.23629, 54.27884, 54.32117, 54.36327, 
    54.40516, 54.44682, 54.48825, 54.52945, 54.57043, 54.61118, 54.65171, 
    54.692, 54.73206, 54.7719, 54.8115, 54.85086, 54.89, 54.9289, 54.96756, 
    55.00599, 55.04418, 55.08213, 55.11985, 55.15733, 55.19456, 55.23156, 
    55.26831, 55.30483, 55.3411, 55.37712, 55.4129, 55.44844, 55.48373, 
    55.51877, 55.55356, 55.58811, 55.62241, 55.65645, 55.69025, 55.72379, 
    55.75708, 55.79012, 55.82291, 55.85543, 55.88771, 55.91973, 55.95149, 
    55.98299, 56.01424, 56.04522, 56.07595, 56.10641, 56.13662, 56.16656, 
    56.19624, 56.22565, 56.25481, 56.2837, 56.31232, 56.34067, 56.36876, 
    56.39658, 56.42413, 56.45142, 56.47843, 56.50517, 56.53164, 56.55785, 
    56.58377, 56.60943, 56.63481, 56.65992, 56.68475, 56.70931, 56.73359, 
    56.7576, 56.78132, 56.80477, 56.82794, 56.85083, 56.87344, 56.89577, 
    56.91782, 56.93959, 56.96108, 56.98228, 57.0032, 57.02384, 57.04419, 
    57.06426, 57.08404, 57.10353, 57.12275, 57.14167, 57.16031, 57.17865, 
    57.19671, 57.21448, 57.23196, 57.24915, 57.26605, 57.28266, 57.29898, 
    57.315, 57.33074, 57.34618, 57.36133, 57.37618, 57.39074, 57.40501, 
    57.41898, 57.43266, 57.44604, 57.45913, 57.47192, 57.48441, 57.4966, 
    57.50851, 57.52011, 57.53141, 57.54242, 57.55312, 57.56353, 57.57364, 
    57.58345, 57.59296, 57.60217, 57.61108, 57.61969, 57.62799, 57.63601, 
    57.64371, 57.65112, 57.65822, 57.66502, 57.67152, 57.67772, 57.68361, 
    57.68921, 57.6945, 57.69948, 57.70417, 57.70855, 57.71263, 57.7164, 
    57.71987, 57.72304, 57.7259, 57.72846, 57.73072, 57.73267, 57.73432, 
    57.73566, 57.7367, 57.73744, 57.73787, 57.738, 57.73782, 57.73734, 
    57.73656, 57.73547, 57.73408, 57.73238, 57.73038, 57.72808, 57.72547, 
    57.72256, 57.71934, 57.71582, 57.712, 57.70787, 57.70345, 57.69872, 
    57.69368, 57.68834, 57.6827, 57.67676, 57.67051, 57.66396, 57.65712, 
    57.64996, 57.64251, 57.63476, 57.6267, 57.61835, 57.60969, 57.60073, 
    57.59147, 57.58192, 57.57206, 57.5619, 57.55145, 57.5407, 57.52964, 
    57.51829, 57.50664, 57.4947, 57.48245, 57.46991, 57.45708, 57.44394, 
    57.43052, 57.41679, 57.40277, 57.38846, 57.37385, 57.35895, 57.34376, 
    57.32827, 57.31249, 57.29642, 57.28005, 57.2634, 57.24645, 57.22921, 
    57.21169, 57.19387, 57.17577, 57.15738, 57.13869, 57.11972, 57.10047, 
    57.08093, 57.0611, 57.04099, 57.02059, 56.99991, 56.97895, 56.9577, 
    56.93616, 56.91435, 56.89226, 56.86988, 56.84723, 56.82429, 56.80108, 
    56.77758, 56.75381, 56.72977, 56.70544, 56.68084, 56.65596, 56.63081, 
    56.60539, 56.57969, 56.55372, 56.52747, 56.50096, 56.47417, 56.44712, 
    56.41979, 56.3922, 56.36433, 56.3362, 56.3078, 56.27914, 56.25021, 
    56.22102, 56.19156, 56.16184, 56.13186, 56.10161, 56.07111, 56.04034, 
    56.00931, 55.97802, 55.94648, 55.91468, 55.88262, 55.8503, 55.81774, 
    55.78491, 55.75183, 55.7185, 55.68492, 55.65108, 55.617, 55.58266, 
    55.54808, 55.51324, 55.47816, 55.44283, 55.40726, 55.37144, 55.33538, 
    55.29907, 55.26252, 55.22573, 55.18869, 55.15142, 55.1139, 55.07615, 
    55.03815, 54.99993, 54.96146, 54.92276, 54.88382, 54.84465, 54.80525, 
    54.76561, 54.72574, 54.68564, 54.64531, 54.60475, 54.56396, 54.52295, 
    54.48171, 54.44024, 54.39854, 54.35663, 54.31449, 54.27212, 54.22953, 
    54.18673, 54.1437, 54.10045, 54.05699, 54.0133, 53.9694, 53.92529, 
    53.88095, 53.83641, 53.79165, 53.74667, 53.70148, 53.65609, 53.61048, 
    53.56466,
  48.59784, 48.6598, 48.72162, 48.7833, 48.84484, 48.90624, 48.96749, 
    49.02861, 49.08958, 49.15041, 49.21109, 49.27163, 49.33202, 49.39227, 
    49.45236, 49.51231, 49.57211, 49.63177, 49.69127, 49.75062, 49.80982, 
    49.86887, 49.92776, 49.9865, 50.04509, 50.10352, 50.1618, 50.21991, 
    50.27788, 50.33568, 50.39333, 50.45081, 50.50814, 50.5653, 50.62231, 
    50.67915, 50.73582, 50.79234, 50.84869, 50.90487, 50.96089, 51.01674, 
    51.07242, 51.12794, 51.18328, 51.23846, 51.29346, 51.3483, 51.40296, 
    51.45745, 51.51176, 51.5659, 51.61987, 51.67366, 51.72727, 51.7807, 
    51.83396, 51.88704, 51.93993, 51.99265, 52.04518, 52.09753, 52.1497, 
    52.20169, 52.25349, 52.3051, 52.35653, 52.40777, 52.45883, 52.50969, 
    52.56036, 52.61085, 52.66114, 52.71125, 52.76115, 52.81087, 52.86039, 
    52.90971, 52.95884, 53.00778, 53.05651, 53.10505, 53.15339, 53.20152, 
    53.24946, 53.2972, 53.34473, 53.39206, 53.43918, 53.4861, 53.53281, 
    53.57932, 53.62562, 53.67171, 53.71759, 53.76326, 53.80872, 53.85397, 
    53.89901, 53.94384, 53.98845, 54.03284, 54.07702, 54.12098, 54.16473, 
    54.20826, 54.25156, 54.29465, 54.33752, 54.38017, 54.42259, 54.46479, 
    54.50677, 54.54852, 54.59004, 54.63134, 54.67242, 54.71326, 54.75388, 
    54.79426, 54.83442, 54.87434, 54.91403, 54.95349, 54.99271, 55.0317, 
    55.07046, 55.10898, 55.14726, 55.1853, 55.22311, 55.26067, 55.298, 
    55.33508, 55.37192, 55.40852, 55.44488, 55.48099, 55.51686, 55.55247, 
    55.58785, 55.62298, 55.65786, 55.69249, 55.72686, 55.76099, 55.79487, 
    55.8285, 55.86187, 55.89499, 55.92786, 55.96046, 55.99282, 56.02492, 
    56.05676, 56.08834, 56.11966, 56.15073, 56.18153, 56.21207, 56.24235, 
    56.27237, 56.30212, 56.33161, 56.36084, 56.3898, 56.4185, 56.44692, 
    56.47508, 56.50298, 56.5306, 56.55795, 56.58503, 56.61185, 56.63839, 
    56.66466, 56.69065, 56.71637, 56.74182, 56.76699, 56.79189, 56.81651, 
    56.84086, 56.86493, 56.88871, 56.91222, 56.93546, 56.95841, 56.98108, 
    57.00347, 57.02558, 57.04741, 57.06895, 57.09021, 57.11118, 57.13188, 
    57.15228, 57.17241, 57.19224, 57.21179, 57.23105, 57.25002, 57.26871, 
    57.28711, 57.30521, 57.32303, 57.34056, 57.3578, 57.37474, 57.3914, 
    57.40776, 57.42383, 57.43961, 57.45509, 57.47028, 57.48518, 57.49978, 
    57.51408, 57.5281, 57.54181, 57.55523, 57.56835, 57.58117, 57.5937, 
    57.60593, 57.61786, 57.6295, 57.64083, 57.65187, 57.66261, 57.67304, 
    57.68318, 57.69302, 57.70255, 57.71179, 57.72072, 57.72935, 57.73769, 
    57.74572, 57.75344, 57.76087, 57.76799, 57.77481, 57.78133, 57.78755, 
    57.79346, 57.79907, 57.80437, 57.80938, 57.81407, 57.81847, 57.82256, 
    57.82634, 57.82982, 57.833, 57.83587, 57.83844, 57.8407, 57.84266, 
    57.84431, 57.84566, 57.8467, 57.84744, 57.84787, 57.848, 57.84782, 
    57.84734, 57.84655, 57.84546, 57.84407, 57.84237, 57.84036, 57.83805, 
    57.83543, 57.83252, 57.82929, 57.82576, 57.82193, 57.81779, 57.81335, 
    57.80861, 57.80355, 57.7982, 57.79255, 57.78659, 57.78032, 57.77376, 
    57.76689, 57.75972, 57.75224, 57.74447, 57.73639, 57.72801, 57.71933, 
    57.71035, 57.70107, 57.69148, 57.68159, 57.67141, 57.66093, 57.65014, 
    57.63906, 57.62768, 57.616, 57.60402, 57.59174, 57.57917, 57.56629, 
    57.55312, 57.53966, 57.5259, 57.51184, 57.49749, 57.48284, 57.4679, 
    57.45266, 57.43713, 57.42131, 57.40519, 57.38878, 57.37208, 57.35509, 
    57.33781, 57.32023, 57.30237, 57.28421, 57.26577, 57.24704, 57.22802, 
    57.20872, 57.18912, 57.16924, 57.14907, 57.12862, 57.10789, 57.08686, 
    57.06556, 57.04397, 57.0221, 56.99995, 56.97751, 56.9548, 56.9318, 
    56.90852, 56.88497, 56.86114, 56.83702, 56.81264, 56.78797, 56.76303, 
    56.73782, 56.71232, 56.68656, 56.66052, 56.63421, 56.60762, 56.58077, 
    56.55364, 56.52625, 56.49858, 56.47065, 56.44244, 56.41397, 56.38523, 
    56.35624, 56.32697, 56.29743, 56.26764, 56.23758, 56.20726, 56.17667, 
    56.14583, 56.11472, 56.08336, 56.05174, 56.01986, 55.98772, 55.95532, 
    55.92267, 55.88977, 55.85661, 55.8232, 55.78953, 55.75561, 55.72144, 
    55.68702, 55.65236, 55.61744, 55.58227, 55.54686, 55.5112, 55.47529, 
    55.43914, 55.40275, 55.36611, 55.32923, 55.29211, 55.25475, 55.21714, 
    55.1793, 55.14122, 55.1029, 55.06434, 55.02555, 54.98653, 54.94726, 
    54.90777, 54.86804, 54.82808, 54.78789, 54.74747, 54.70681, 54.66594, 
    54.62482, 54.58349, 54.54193, 54.50014, 54.45813, 54.41589, 54.37344, 
    54.33075, 54.28785, 54.24473, 54.20139, 54.15782, 54.11404, 54.07005, 
    54.02583, 53.9814, 53.93676, 53.8919, 53.84683, 53.80155, 53.75605, 
    53.71035, 53.66443,
  48.68832, 48.75037, 48.81229, 48.87407, 48.9357, 48.9972, 49.05855, 
    49.11977, 49.18083, 49.24176, 49.30254, 49.36317, 49.42366, 49.484, 
    49.5442, 49.60425, 49.66415, 49.7239, 49.7835, 49.84295, 49.90225, 
    49.9614, 50.02039, 50.07923, 50.13792, 50.19645, 50.25482, 50.31304, 
    50.3711, 50.429, 50.48675, 50.54434, 50.60176, 50.65903, 50.71613, 
    50.77307, 50.82985, 50.88646, 50.94291, 50.9992, 51.05532, 51.11127, 
    51.16705, 51.22267, 51.27811, 51.33339, 51.3885, 51.44343, 51.49819, 
    51.55278, 51.6072, 51.66144, 51.7155, 51.76939, 51.8231, 51.87664, 51.93, 
    51.98318, 52.03617, 52.08899, 52.14162, 52.19408, 52.24635, 52.29843, 
    52.35033, 52.40205, 52.45358, 52.50492, 52.55607, 52.60704, 52.65781, 
    52.7084, 52.75879, 52.80899, 52.859, 52.90882, 52.95844, 53.00787, 
    53.05709, 53.10613, 53.15496, 53.2036, 53.25203, 53.30027, 53.34831, 
    53.39614, 53.44377, 53.4912, 53.53842, 53.58544, 53.63226, 53.67886, 
    53.72526, 53.77145, 53.81742, 53.8632, 53.90876, 53.9541, 53.99924, 
    54.04416, 54.08886, 54.13336, 54.17763, 54.22169, 54.26553, 54.30916, 
    54.35256, 54.39574, 54.43871, 54.48145, 54.52397, 54.56626, 54.60833, 
    54.65018, 54.6918, 54.73319, 54.77436, 54.8153, 54.856, 54.89648, 
    54.93673, 54.97675, 55.01653, 55.05608, 55.09539, 55.13447, 55.17332, 
    55.21193, 55.2503, 55.28843, 55.32632, 55.36398, 55.40139, 55.43856, 
    55.47549, 55.51218, 55.54862, 55.58482, 55.62077, 55.65648, 55.69194, 
    55.72715, 55.76212, 55.79683, 55.83129, 55.86551, 55.89947, 55.93317, 
    55.96663, 55.99983, 56.03278, 56.06547, 56.0979, 56.13008, 56.162, 
    56.19366, 56.22506, 56.2562, 56.28708, 56.3177, 56.34806, 56.37815, 
    56.40798, 56.43755, 56.46685, 56.49588, 56.52465, 56.55315, 56.58138, 
    56.60935, 56.63704, 56.66447, 56.69162, 56.7185, 56.74511, 56.77145, 
    56.79751, 56.8233, 56.84882, 56.87405, 56.89902, 56.9237, 56.94811, 
    56.97224, 56.99609, 57.01967, 57.04296, 57.06597, 57.0887, 57.11115, 
    57.13332, 57.1552, 57.17681, 57.19812, 57.21916, 57.2399, 57.26036, 
    57.28054, 57.30043, 57.32003, 57.33934, 57.35837, 57.37711, 57.39555, 
    57.41371, 57.43158, 57.44915, 57.46644, 57.48343, 57.50013, 57.51654, 
    57.53265, 57.54847, 57.564, 57.57923, 57.59417, 57.60881, 57.62315, 
    57.6372, 57.65096, 57.66441, 57.67757, 57.69043, 57.70299, 57.71526, 
    57.72722, 57.73888, 57.75025, 57.76132, 57.77208, 57.78255, 57.79272, 
    57.80258, 57.81215, 57.8214, 57.83036, 57.83902, 57.84738, 57.85543, 
    57.86318, 57.87063, 57.87777, 57.88461, 57.89115, 57.89738, 57.90331, 
    57.90893, 57.91425, 57.91927, 57.92398, 57.92838, 57.93248, 57.93628, 
    57.93977, 57.94296, 57.94584, 57.94841, 57.95068, 57.95264, 57.9543, 
    57.95565, 57.9567, 57.95744, 57.95787, 57.958, 57.95782, 57.95734, 
    57.95655, 57.95546, 57.95406, 57.95235, 57.95034, 57.94802, 57.9454, 
    57.94247, 57.93924, 57.9357, 57.93185, 57.9277, 57.92325, 57.91849, 
    57.91343, 57.90806, 57.90239, 57.89641, 57.89013, 57.88355, 57.87666, 
    57.86947, 57.86197, 57.85418, 57.84608, 57.83767, 57.82897, 57.81996, 
    57.81065, 57.80104, 57.79113, 57.78091, 57.7704, 57.75959, 57.74847, 
    57.73706, 57.72535, 57.71333, 57.70102, 57.68841, 57.67551, 57.6623, 
    57.6488, 57.635, 57.6209, 57.60651, 57.59182, 57.57684, 57.56156, 
    57.54599, 57.53012, 57.51396, 57.49751, 57.48076, 57.46372, 57.44639, 
    57.42877, 57.41086, 57.39265, 57.37416, 57.35538, 57.33631, 57.31695, 
    57.2973, 57.27737, 57.25715, 57.23664, 57.21585, 57.19477, 57.17341, 
    57.15176, 57.12983, 57.10762, 57.08513, 57.06235, 57.0393, 57.01596, 
    56.99234, 56.96844, 56.94427, 56.91982, 56.89509, 56.87008, 56.8448, 
    56.81924, 56.79341, 56.7673, 56.74092, 56.71427, 56.68734, 56.66014, 
    56.63268, 56.60494, 56.57693, 56.54866, 56.52012, 56.49131, 56.46223, 
    56.43289, 56.40328, 56.37341, 56.34327, 56.31288, 56.28222, 56.25129, 
    56.22011, 56.18867, 56.15697, 56.12501, 56.09279, 56.06031, 56.02758, 
    55.99459, 55.96135, 55.92786, 55.89411, 55.86011, 55.82586, 55.79136, 
    55.7566, 55.7216, 55.68635, 55.65085, 55.6151, 55.57911, 55.54287, 
    55.50639, 55.46967, 55.4327, 55.39549, 55.35804, 55.32035, 55.28241, 
    55.24424, 55.20584, 55.16719, 55.12831, 55.08919, 55.04984, 55.01025, 
    54.97043, 54.93038, 54.89009, 54.84958, 54.80883, 54.76786, 54.72666, 
    54.68523, 54.64357, 54.60169, 54.55959, 54.51726, 54.4747, 54.43193, 
    54.38893, 54.34571, 54.30227, 54.25861, 54.21474, 54.17064, 54.12634, 
    54.08181, 54.03707, 53.99211, 53.94695, 53.90156, 53.85597, 53.81017, 
    53.76415,
  48.77872, 48.84087, 48.90288, 48.96476, 49.02649, 49.08808, 49.14953, 
    49.21084, 49.27201, 49.33303, 49.39391, 49.45464, 49.51523, 49.57567, 
    49.63597, 49.69611, 49.75611, 49.81596, 49.87566, 49.93521, 49.99461, 
    50.05385, 50.11295, 50.17188, 50.23067, 50.2893, 50.34777, 50.40609, 
    50.46426, 50.52226, 50.5801, 50.63779, 50.69532, 50.75268, 50.80988, 
    50.86693, 50.92381, 50.98052, 51.03707, 51.09346, 51.14967, 51.20573, 
    51.26161, 51.31733, 51.37288, 51.42825, 51.48346, 51.53849, 51.59336, 
    51.64805, 51.70256, 51.7569, 51.81107, 51.86506, 51.91888, 51.97252, 
    52.02597, 52.07925, 52.13235, 52.18527, 52.238, 52.29056, 52.34293, 
    52.39511, 52.44712, 52.49893, 52.55056, 52.60201, 52.65326, 52.70433, 
    52.7552, 52.80589, 52.85638, 52.90668, 52.95679, 53.00671, 53.05643, 
    53.10596, 53.15529, 53.20442, 53.25336, 53.30209, 53.35063, 53.39896, 
    53.4471, 53.49503, 53.54276, 53.59029, 53.63762, 53.68473, 53.73164, 
    53.77835, 53.82484, 53.87113, 53.91721, 53.96308, 54.00874, 54.05418, 
    54.09941, 54.14443, 54.18924, 54.23383, 54.2782, 54.32235, 54.36629, 
    54.41001, 54.45351, 54.49679, 54.53985, 54.58269, 54.6253, 54.66769, 
    54.70985, 54.7518, 54.79351, 54.835, 54.87626, 54.91729, 54.95809, 
    54.99866, 55.039, 55.07911, 55.11898, 55.15863, 55.19803, 55.23721, 
    55.27614, 55.31484, 55.3533, 55.39152, 55.42951, 55.46725, 55.50475, 
    55.54201, 55.57903, 55.61581, 55.65234, 55.68862, 55.72466, 55.76045, 
    55.796, 55.8313, 55.86634, 55.90114, 55.93569, 55.96999, 56.00403, 
    56.03782, 56.07136, 56.10464, 56.13767, 56.17044, 56.20296, 56.23521, 
    56.26722, 56.29895, 56.33044, 56.36166, 56.39261, 56.42331, 56.45374, 
    56.48391, 56.51382, 56.54346, 56.57283, 56.60194, 56.63079, 56.65936, 
    56.68766, 56.7157, 56.74347, 56.77096, 56.79818, 56.82514, 56.85181, 
    56.87822, 56.90435, 56.93021, 56.95579, 56.98109, 57.00613, 57.03088, 
    57.05535, 57.07954, 57.10346, 57.12709, 57.15045, 57.17352, 57.19632, 
    57.21882, 57.24105, 57.26299, 57.28465, 57.30603, 57.32712, 57.34792, 
    57.36844, 57.38867, 57.40861, 57.42826, 57.44763, 57.46671, 57.48549, 
    57.50399, 57.5222, 57.54011, 57.55774, 57.57507, 57.59211, 57.60885, 
    57.62531, 57.64146, 57.65733, 57.6729, 57.68817, 57.70315, 57.71783, 
    57.73222, 57.7463, 57.76009, 57.77359, 57.78678, 57.79968, 57.81227, 
    57.82457, 57.83657, 57.84827, 57.85967, 57.87077, 57.88156, 57.89206, 
    57.90225, 57.91214, 57.92173, 57.93102, 57.94001, 57.94869, 57.95707, 
    57.96514, 57.97291, 57.98038, 57.98755, 57.9944, 58.00096, 58.00721, 
    58.01315, 58.01879, 58.02413, 58.02916, 58.03388, 58.0383, 58.04241, 
    58.04622, 58.04972, 58.05291, 58.0558, 58.05838, 58.06066, 58.06263, 
    58.06429, 58.06564, 58.06669, 58.06743, 58.06787, 58.068, 58.06782, 
    58.06734, 58.06655, 58.06545, 58.06404, 58.06233, 58.06032, 58.05799, 
    58.05536, 58.05243, 58.04918, 58.04564, 58.04178, 58.03762, 58.03315, 
    58.02838, 58.0233, 58.01792, 58.01223, 58.00624, 57.99994, 57.99334, 
    57.98643, 57.97922, 57.9717, 57.96388, 57.95576, 57.94733, 57.9386, 
    57.92957, 57.92023, 57.9106, 57.90066, 57.89042, 57.87988, 57.86903, 
    57.85788, 57.84644, 57.83469, 57.82265, 57.8103, 57.79766, 57.78471, 
    57.77147, 57.75793, 57.74409, 57.72996, 57.71553, 57.7008, 57.68577, 
    57.67045, 57.65484, 57.63893, 57.62272, 57.60622, 57.58943, 57.57235, 
    57.55497, 57.5373, 57.51934, 57.50108, 57.48254, 57.46371, 57.44458, 
    57.42517, 57.40548, 57.38549, 57.36521, 57.34465, 57.3238, 57.30267, 
    57.28125, 57.25954, 57.23755, 57.21528, 57.19273, 57.16989, 57.14677, 
    57.12337, 57.09969, 57.07573, 57.05149, 57.02698, 57.00219, 56.97711, 
    56.95176, 56.92614, 56.90024, 56.87406, 56.84761, 56.82089, 56.7939, 
    56.76663, 56.73909, 56.71128, 56.6832, 56.65486, 56.62624, 56.59736, 
    56.56821, 56.53879, 56.50911, 56.47916, 56.44895, 56.41847, 56.38773, 
    56.35674, 56.32547, 56.29395, 56.26217, 56.23013, 56.19783, 56.16528, 
    56.13247, 56.0994, 56.06607, 56.03249, 55.99866, 55.96458, 55.93024, 
    55.89565, 55.86082, 55.82573, 55.79039, 55.75481, 55.71898, 55.6829, 
    55.64657, 55.61, 55.57319, 55.53614, 55.49884, 55.4613, 55.42352, 
    55.38549, 55.34723, 55.30873, 55.27, 55.23102, 55.19181, 55.15237, 
    55.11269, 55.07278, 55.03263, 54.99226, 54.95165, 54.91081, 54.86975, 
    54.82845, 54.78693, 54.74518, 54.7032, 54.661, 54.61857, 54.57592, 
    54.53305, 54.48996, 54.44664, 54.40311, 54.35936, 54.31538, 54.27119, 
    54.22678, 54.18216, 54.13733, 54.09227, 54.047, 54.00153, 53.95584, 
    53.90993, 53.86382,
  48.86904, 48.93129, 48.9934, 49.05537, 49.1172, 49.17889, 49.24044, 
    49.30184, 49.36311, 49.42423, 49.4852, 49.54604, 49.60672, 49.66726, 
    49.72765, 49.7879, 49.848, 49.90794, 49.96774, 50.02739, 50.08689, 
    50.14623, 50.20543, 50.26447, 50.32335, 50.38208, 50.44065, 50.49907, 
    50.55733, 50.61544, 50.67339, 50.73117, 50.7888, 50.84626, 50.90357, 
    50.96071, 51.01769, 51.0745, 51.13116, 51.18764, 51.24396, 51.30011, 
    51.3561, 51.41192, 51.46757, 51.52304, 51.57835, 51.63349, 51.68845, 
    51.74325, 51.79786, 51.85231, 51.90658, 51.96067, 52.01458, 52.06832, 
    52.12188, 52.17526, 52.22846, 52.28148, 52.33432, 52.38697, 52.43945, 
    52.49173, 52.54384, 52.59576, 52.64749, 52.69903, 52.75039, 52.80156, 
    52.85253, 52.90332, 52.95391, 53.00432, 53.05453, 53.10455, 53.15437, 
    53.20399, 53.25343, 53.30266, 53.35169, 53.40053, 53.44917, 53.4976, 
    53.54584, 53.59387, 53.6417, 53.68933, 53.73675, 53.78397, 53.83098, 
    53.87778, 53.92438, 53.97076, 54.01694, 54.06291, 54.10867, 54.15421, 
    54.19954, 54.24466, 54.28955, 54.33424, 54.37871, 54.42297, 54.467, 
    54.51082, 54.55441, 54.59779, 54.64095, 54.68388, 54.72659, 54.76907, 
    54.81133, 54.85337, 54.89518, 54.93676, 54.97812, 55.01924, 55.06013, 
    55.1008, 55.14123, 55.18143, 55.2214, 55.26114, 55.30063, 55.3399, 
    55.37892, 55.41771, 55.45626, 55.49458, 55.53265, 55.57048, 55.60807, 
    55.64542, 55.68253, 55.71939, 55.75601, 55.79239, 55.82851, 55.86439, 
    55.90002, 55.93541, 55.97054, 56.00542, 56.04005, 56.07444, 56.10857, 
    56.14244, 56.17606, 56.20943, 56.24253, 56.27539, 56.30799, 56.34032, 
    56.3724, 56.40422, 56.43578, 56.46708, 56.49812, 56.52889, 56.5594, 
    56.58965, 56.61963, 56.64935, 56.6788, 56.70798, 56.7369, 56.76554, 
    56.79392, 56.82203, 56.84987, 56.87744, 56.90473, 56.93175, 56.9585, 
    56.98498, 57.01118, 57.0371, 57.06275, 57.08812, 57.11322, 57.13803, 
    57.16257, 57.18683, 57.21081, 57.2345, 57.25792, 57.28106, 57.30391, 
    57.32648, 57.34877, 57.37077, 57.39249, 57.41392, 57.43507, 57.45592, 
    57.4765, 57.49678, 57.51678, 57.53648, 57.5559, 57.57503, 57.59387, 
    57.61242, 57.63068, 57.64864, 57.66631, 57.68369, 57.70078, 57.71757, 
    57.73407, 57.75027, 57.76617, 57.78179, 57.7971, 57.81212, 57.82685, 
    57.84127, 57.8554, 57.86923, 57.88276, 57.89599, 57.90892, 57.92155, 
    57.93389, 57.94592, 57.95765, 57.96908, 57.98021, 57.99104, 58.00156, 
    58.01178, 58.0217, 58.03132, 58.04063, 58.04964, 58.05835, 58.06675, 
    58.07485, 58.08264, 58.09013, 58.09732, 58.10419, 58.11077, 58.11703, 
    58.123, 58.12865, 58.134, 58.13905, 58.14378, 58.14821, 58.15234, 
    58.15615, 58.15966, 58.16287, 58.16576, 58.16835, 58.17064, 58.17261, 
    58.17428, 58.17564, 58.17669, 58.17743, 58.17787, 58.178, 58.17782, 
    58.17733, 58.17654, 58.17544, 58.17403, 58.17232, 58.1703, 58.16796, 
    58.16533, 58.16238, 58.15913, 58.15557, 58.15171, 58.14753, 58.14305, 
    58.13827, 58.13317, 58.12778, 58.12207, 58.11606, 58.10975, 58.10313, 
    58.0962, 58.08897, 58.08143, 58.07359, 58.06544, 58.05699, 58.04824, 
    58.03918, 58.02982, 58.02015, 58.01019, 57.99992, 57.98934, 57.97847, 
    57.96729, 57.95581, 57.94403, 57.93196, 57.91957, 57.90689, 57.89392, 
    57.88064, 57.86706, 57.85318, 57.83901, 57.82454, 57.80977, 57.7947, 
    57.77934, 57.76368, 57.74773, 57.73148, 57.71493, 57.69809, 57.68096, 
    57.66354, 57.64582, 57.62781, 57.6095, 57.59091, 57.57203, 57.55285, 
    57.53339, 57.51363, 57.49359, 57.47326, 57.45264, 57.43174, 57.41055, 
    57.38907, 57.36731, 57.34526, 57.32293, 57.30032, 57.27742, 57.25424, 
    57.23077, 57.20703, 57.18301, 57.15871, 57.13412, 57.10926, 57.08413, 
    57.05871, 57.03302, 57.00705, 56.98081, 56.95429, 56.9275, 56.90043, 
    56.87309, 56.84549, 56.8176, 56.78945, 56.76103, 56.73234, 56.70338, 
    56.67416, 56.64466, 56.61491, 56.58488, 56.5546, 56.52404, 56.49323, 
    56.46215, 56.43081, 56.39921, 56.36735, 56.33523, 56.30285, 56.27021, 
    56.23732, 56.20417, 56.17076, 56.1371, 56.10318, 56.06902, 56.0346, 
    55.99992, 55.965, 55.92982, 55.89441, 55.85873, 55.82281, 55.78665, 
    55.75024, 55.71358, 55.67668, 55.63953, 55.60215, 55.56451, 55.52665, 
    55.48853, 55.45018, 55.41159, 55.37276, 55.3337, 55.2944, 55.25486, 
    55.21509, 55.17509, 55.13485, 55.09438, 55.05368, 55.01275, 54.97159, 
    54.9302, 54.88858, 54.84673, 54.80466, 54.76237, 54.71984, 54.6771, 
    54.63413, 54.59094, 54.54753, 54.5039, 54.46005, 54.41598, 54.37169, 
    54.32719, 54.28247, 54.23753, 54.19238, 54.14702, 54.10144, 54.05565, 
    54.00965, 53.96344,
  48.95928, 49.02163, 49.08383, 49.1459, 49.20783, 49.26962, 49.33126, 
    49.39277, 49.45413, 49.51535, 49.57642, 49.63735, 49.69814, 49.75877, 
    49.81927, 49.87961, 49.93981, 49.99986, 50.05975, 50.1195, 50.1791, 
    50.23854, 50.29783, 50.35697, 50.41596, 50.47479, 50.53346, 50.59198, 
    50.65034, 50.70855, 50.76659, 50.82448, 50.88221, 50.93977, 50.99718, 
    51.05442, 51.1115, 51.16842, 51.22517, 51.28176, 51.33818, 51.39444, 
    51.45052, 51.50644, 51.56219, 51.61777, 51.67318, 51.72842, 51.78349, 
    51.83838, 51.8931, 51.94764, 52.00201, 52.05621, 52.11023, 52.16406, 
    52.21772, 52.27121, 52.32451, 52.37763, 52.43057, 52.48333, 52.5359, 
    52.58829, 52.6405, 52.69252, 52.74435, 52.79599, 52.84745, 52.89872, 
    52.9498, 53.00069, 53.05138, 53.10189, 53.1522, 53.20232, 53.25224, 
    53.30197, 53.3515, 53.40084, 53.44997, 53.49891, 53.54765, 53.59618, 
    53.64452, 53.69265, 53.74059, 53.78831, 53.83583, 53.88315, 53.93026, 
    53.97717, 54.02386, 54.07035, 54.11662, 54.16269, 54.20854, 54.25418, 
    54.29961, 54.34483, 54.38983, 54.43461, 54.47918, 54.52353, 54.56767, 
    54.61158, 54.65527, 54.69874, 54.74199, 54.78502, 54.82783, 54.87041, 
    54.91277, 54.9549, 54.9968, 55.03848, 55.07993, 55.12115, 55.16214, 
    55.20289, 55.24342, 55.28371, 55.32378, 55.3636, 55.40319, 55.44255, 
    55.48167, 55.52055, 55.55919, 55.5976, 55.63576, 55.67368, 55.71136, 
    55.7488, 55.786, 55.82295, 55.85966, 55.89611, 55.93233, 55.9683, 
    56.00402, 56.03949, 56.0747, 56.10967, 56.14439, 56.17886, 56.21307, 
    56.24703, 56.28073, 56.31418, 56.34737, 56.38031, 56.41299, 56.4454, 
    56.47757, 56.50946, 56.5411, 56.57248, 56.6036, 56.63445, 56.66504, 
    56.69536, 56.72542, 56.75521, 56.78474, 56.814, 56.84299, 56.87171, 
    56.90016, 56.92834, 56.95625, 56.98389, 57.01126, 57.03835, 57.06517, 
    57.09171, 57.11798, 57.14397, 57.16969, 57.19513, 57.22029, 57.24517, 
    57.26978, 57.2941, 57.31814, 57.3419, 57.36538, 57.38858, 57.41149, 
    57.43412, 57.45647, 57.47853, 57.50031, 57.5218, 57.543, 57.56392, 
    57.58455, 57.60489, 57.62494, 57.6447, 57.66417, 57.68335, 57.70224, 
    57.72084, 57.73914, 57.75716, 57.77488, 57.7923, 57.80944, 57.82627, 
    57.84282, 57.85907, 57.87502, 57.89067, 57.90603, 57.92109, 57.93586, 
    57.95032, 57.96449, 57.97836, 57.99192, 58.00519, 58.01816, 58.03083, 
    58.0432, 58.05526, 58.06702, 58.07849, 58.08965, 58.10051, 58.11106, 
    58.12131, 58.13126, 58.1409, 58.15024, 58.15928, 58.16801, 58.17643, 
    58.18456, 58.19237, 58.19988, 58.20708, 58.21399, 58.22058, 58.22686, 
    58.23284, 58.23851, 58.24388, 58.24894, 58.25368, 58.25813, 58.26226, 
    58.26609, 58.26961, 58.27282, 58.27573, 58.27832, 58.28061, 58.28259, 
    58.28427, 58.28563, 58.28669, 58.28743, 58.28787, 58.288, 58.28782, 
    58.28733, 58.28654, 58.28543, 58.28402, 58.2823, 58.28027, 58.27794, 
    58.27529, 58.27234, 58.26908, 58.26551, 58.26163, 58.25745, 58.25295, 
    58.24815, 58.24305, 58.23764, 58.23191, 58.22589, 58.21955, 58.21291, 
    58.20597, 58.19872, 58.19115, 58.18329, 58.17512, 58.16665, 58.15787, 
    58.14878, 58.1394, 58.12971, 58.11971, 58.10941, 58.09881, 58.0879, 
    58.07669, 58.06519, 58.05337, 58.04126, 58.02885, 58.01613, 58.00311, 
    57.9898, 57.97618, 57.96227, 57.94805, 57.93354, 57.91873, 57.90362, 
    57.88822, 57.87251, 57.85652, 57.84022, 57.82363, 57.80675, 57.78957, 
    57.77209, 57.75433, 57.73627, 57.71791, 57.69927, 57.68034, 57.66111, 
    57.64159, 57.62178, 57.60168, 57.5813, 57.56063, 57.53967, 57.51842, 
    57.49688, 57.47506, 57.45295, 57.43056, 57.40789, 57.38493, 57.36169, 
    57.33816, 57.31436, 57.29027, 57.2659, 57.24125, 57.21633, 57.19112, 
    57.16564, 57.13988, 57.11384, 57.08753, 57.06094, 57.03408, 57.00695, 
    56.97954, 56.95185, 56.9239, 56.89568, 56.86718, 56.83842, 56.80939, 
    56.78009, 56.75052, 56.72068, 56.69058, 56.66022, 56.62959, 56.59869, 
    56.56754, 56.53612, 56.50444, 56.4725, 56.4403, 56.40783, 56.37511, 
    56.34214, 56.30891, 56.27542, 56.24167, 56.20767, 56.17342, 56.13892, 
    56.10416, 56.06915, 56.03389, 55.99838, 55.96262, 55.92662, 55.89037, 
    55.85387, 55.81712, 55.78013, 55.7429, 55.70542, 55.6677, 55.62974, 
    55.59154, 55.5531, 55.51442, 55.47549, 55.43634, 55.39695, 55.35732, 
    55.31746, 55.27736, 55.23703, 55.19646, 55.15567, 55.11464, 55.07339, 
    55.0319, 54.99019, 54.94825, 54.90608, 54.86369, 54.82107, 54.77823, 
    54.73517, 54.69188, 54.64837, 54.60464, 54.5607, 54.51653, 54.47215, 
    54.42754, 54.38272, 54.33769, 54.29244, 54.24698, 54.2013, 54.15541, 
    54.10931, 54.06301,
  49.04944, 49.11188, 49.17419, 49.23635, 49.29838, 49.36026, 49.42201, 
    49.48361, 49.54507, 49.60639, 49.66756, 49.72859, 49.78947, 49.85021, 
    49.9108, 49.97124, 50.03154, 50.09169, 50.15168, 50.21153, 50.27123, 
    50.33077, 50.39016, 50.4494, 50.50849, 50.56742, 50.62619, 50.68481, 
    50.74328, 50.80158, 50.85973, 50.91772, 50.97554, 51.03321, 51.09072, 
    51.14806, 51.20525, 51.26226, 51.31911, 51.3758, 51.43233, 51.48869, 
    51.54487, 51.60089, 51.65675, 51.71243, 51.76794, 51.82328, 51.87845, 
    51.93344, 51.98826, 52.04291, 52.09739, 52.15168, 52.2058, 52.25974, 
    52.3135, 52.36709, 52.42049, 52.47372, 52.52676, 52.57962, 52.63229, 
    52.68478, 52.73709, 52.78921, 52.84115, 52.89289, 52.94445, 52.99583, 
    53.047, 53.098, 53.1488, 53.1994, 53.24982, 53.30003, 53.35006, 53.39989, 
    53.44952, 53.49896, 53.54819, 53.59723, 53.64607, 53.69471, 53.74314, 
    53.79138, 53.83941, 53.88724, 53.93486, 53.98228, 54.02949, 54.07649, 
    54.12329, 54.16987, 54.21625, 54.26241, 54.30837, 54.35411, 54.39964, 
    54.44495, 54.49005, 54.53493, 54.5796, 54.62405, 54.66828, 54.71229, 
    54.75608, 54.79965, 54.843, 54.88612, 54.92902, 54.9717, 55.01416, 
    55.05638, 55.09838, 55.14015, 55.1817, 55.22301, 55.2641, 55.30495, 
    55.34557, 55.38596, 55.42611, 55.46603, 55.50571, 55.54516, 55.58437, 
    55.62334, 55.66208, 55.70058, 55.73883, 55.77684, 55.81461, 55.85214, 
    55.88943, 55.92647, 55.96326, 55.99981, 56.03611, 56.07217, 56.10798, 
    56.14353, 56.17884, 56.21389, 56.2487, 56.28325, 56.31754, 56.35159, 
    56.38537, 56.4189, 56.45218, 56.4852, 56.51796, 56.55046, 56.5827, 
    56.61468, 56.6464, 56.67786, 56.70905, 56.73998, 56.77065, 56.80105, 
    56.83119, 56.86106, 56.89066, 56.91999, 56.94906, 56.97785, 57.00638, 
    57.03463, 57.06261, 57.09032, 57.11776, 57.14492, 57.17181, 57.19843, 
    57.22477, 57.25083, 57.27661, 57.30212, 57.32735, 57.35229, 57.37696, 
    57.40135, 57.42546, 57.44928, 57.47282, 57.49609, 57.51906, 57.54175, 
    57.56416, 57.58628, 57.60811, 57.62966, 57.65092, 57.67189, 57.69258, 
    57.71297, 57.73308, 57.7529, 57.77242, 57.79166, 57.8106, 57.82925, 
    57.8476, 57.86567, 57.88343, 57.90091, 57.91809, 57.93497, 57.95156, 
    57.96786, 57.98385, 57.99955, 58.01495, 58.03006, 58.04486, 58.05937, 
    58.07357, 58.08748, 58.10109, 58.11439, 58.1274, 58.1401, 58.1525, 
    58.1646, 58.1764, 58.18789, 58.19909, 58.20997, 58.22056, 58.23084, 
    58.24081, 58.25048, 58.25985, 58.26891, 58.27767, 58.28612, 58.29426, 
    58.3021, 58.30963, 58.31686, 58.32377, 58.33038, 58.33669, 58.34268, 
    58.34837, 58.35375, 58.35882, 58.36359, 58.36804, 58.37219, 58.37603, 
    58.37956, 58.38278, 58.38569, 58.3883, 58.39059, 58.39258, 58.39426, 
    58.39562, 58.39668, 58.39743, 58.39787, 58.398, 58.39782, 58.39733, 
    58.39653, 58.39543, 58.39401, 58.39228, 58.39025, 58.38791, 58.38525, 
    58.38229, 58.37902, 58.37544, 58.37156, 58.36736, 58.36285, 58.35804, 
    58.35292, 58.34749, 58.34175, 58.33571, 58.32936, 58.3227, 58.31573, 
    58.30846, 58.30088, 58.29299, 58.2848, 58.2763, 58.2675, 58.25839, 
    58.24897, 58.23925, 58.22923, 58.2189, 58.20827, 58.19733, 58.1861, 
    58.17455, 58.16271, 58.15056, 58.13811, 58.12536, 58.11231, 58.09895, 
    58.0853, 58.07135, 58.05709, 58.04254, 58.02769, 58.01254, 57.99709, 
    57.98134, 57.9653, 57.94896, 57.93232, 57.91539, 57.89817, 57.88065, 
    57.86283, 57.84472, 57.82632, 57.80762, 57.78863, 57.76935, 57.74978, 
    57.72992, 57.70977, 57.68933, 57.6686, 57.64758, 57.62627, 57.60468, 
    57.5828, 57.56063, 57.53818, 57.51545, 57.49242, 57.46912, 57.44553, 
    57.42166, 57.39751, 57.37308, 57.34837, 57.32337, 57.2981, 57.27255, 
    57.24672, 57.22062, 57.19424, 57.16758, 57.14065, 57.11344, 57.08596, 
    57.0582, 57.03018, 57.00188, 56.97332, 56.94448, 56.91537, 56.88599, 
    56.85635, 56.82644, 56.79626, 56.76582, 56.73511, 56.70414, 56.6729, 
    56.6414, 56.60964, 56.57762, 56.54533, 56.51279, 56.47999, 56.44693, 
    56.41362, 56.38004, 56.34622, 56.31213, 56.2778, 56.24321, 56.20836, 
    56.17327, 56.13792, 56.10233, 56.06648, 56.03039, 55.99405, 55.95746, 
    55.92062, 55.88354, 55.84622, 55.80865, 55.77085, 55.7328, 55.6945, 
    55.65597, 55.6172, 55.57819, 55.53894, 55.49945, 55.45973, 55.41977, 
    55.37958, 55.33916, 55.2985, 55.25761, 55.21649, 55.17514, 55.13356, 
    55.09175, 55.04972, 55.00745, 54.96497, 54.92225, 54.87932, 54.83615, 
    54.79277, 54.74917, 54.70534, 54.6613, 54.61703, 54.57255, 54.52785, 
    54.48293, 54.4378, 54.39245, 54.34689, 54.30111, 54.25513, 54.20893, 
    54.16252,
  49.13952, 49.20206, 49.26446, 49.32673, 49.38885, 49.45083, 49.51268, 
    49.57438, 49.63593, 49.69735, 49.75862, 49.81975, 49.88073, 49.94157, 
    50.00226, 50.0628, 50.1232, 50.18344, 50.24354, 50.30349, 50.36329, 
    50.42293, 50.48242, 50.54176, 50.60094, 50.65998, 50.71885, 50.77757, 
    50.83614, 50.89454, 50.95279, 51.01088, 51.06881, 51.12658, 51.18419, 
    51.24163, 51.29892, 51.35603, 51.41299, 51.46978, 51.52641, 51.58286, 
    51.63915, 51.69527, 51.75123, 51.80701, 51.86263, 51.91807, 51.97334, 
    52.02844, 52.08336, 52.13811, 52.19268, 52.24709, 52.30131, 52.35535, 
    52.40922, 52.4629, 52.51641, 52.56974, 52.62288, 52.67584, 52.72862, 
    52.78121, 52.83362, 52.88585, 52.93789, 52.98973, 53.0414, 53.09287, 
    53.14415, 53.19524, 53.24614, 53.29685, 53.34737, 53.39769, 53.44782, 
    53.49775, 53.54748, 53.59702, 53.64636, 53.6955, 53.74444, 53.79318, 
    53.84172, 53.89005, 53.93818, 53.98611, 54.03384, 54.08135, 54.12866, 
    54.17577, 54.22266, 54.26935, 54.31582, 54.36209, 54.40814, 54.45398, 
    54.49961, 54.54502, 54.59022, 54.6352, 54.67997, 54.72451, 54.76884, 
    54.81295, 54.85684, 54.90051, 54.94395, 54.98717, 55.03017, 55.07295, 
    55.1155, 55.15782, 55.19992, 55.24178, 55.28342, 55.32483, 55.36601, 
    55.40696, 55.44767, 55.48816, 55.5284, 55.56842, 55.60819, 55.64774, 
    55.68704, 55.7261, 55.76493, 55.80352, 55.84186, 55.87997, 55.91783, 
    55.95545, 55.99282, 56.02995, 56.06684, 56.10347, 56.13986, 56.17601, 
    56.2119, 56.24754, 56.28294, 56.31808, 56.35297, 56.3876, 56.42198, 
    56.45611, 56.48998, 56.5236, 56.55696, 56.59006, 56.6229, 56.65548, 
    56.68781, 56.71987, 56.75167, 56.78321, 56.81448, 56.84549, 56.87624, 
    56.90672, 56.93693, 56.96687, 56.99655, 57.02596, 57.0551, 57.08397, 
    57.11257, 57.1409, 57.16896, 57.19674, 57.22425, 57.25148, 57.27844, 
    57.30513, 57.33153, 57.35766, 57.38351, 57.40909, 57.43438, 57.4594, 
    57.48413, 57.50859, 57.53276, 57.55665, 57.58025, 57.60358, 57.62661, 
    57.64936, 57.67183, 57.69402, 57.71591, 57.73751, 57.75883, 57.77987, 
    57.80061, 57.82106, 57.84122, 57.86108, 57.88066, 57.89995, 57.91895, 
    57.93764, 57.95605, 57.97417, 57.99199, 58.00951, 58.02674, 58.04367, 
    58.0603, 58.07664, 58.09268, 58.10843, 58.12387, 58.13902, 58.15386, 
    58.16841, 58.18265, 58.1966, 58.21024, 58.22359, 58.23663, 58.24937, 
    58.2618, 58.27394, 58.28577, 58.29729, 58.30852, 58.31944, 58.33005, 
    58.34036, 58.35036, 58.36006, 58.36946, 58.37854, 58.38732, 58.3958, 
    58.40396, 58.41182, 58.41938, 58.42662, 58.43356, 58.44019, 58.44651, 
    58.45252, 58.45823, 58.46362, 58.46871, 58.47349, 58.47796, 58.48212, 
    58.48597, 58.48951, 58.49274, 58.49566, 58.49827, 58.50057, 58.50256, 
    58.50425, 58.50562, 58.50668, 58.50743, 58.50787, 58.508, 58.50782, 
    58.50733, 58.50653, 58.50542, 58.504, 58.50227, 58.50023, 58.49788, 
    58.49522, 58.49225, 58.48897, 58.48538, 58.48148, 58.47727, 58.47275, 
    58.46793, 58.46279, 58.45735, 58.45159, 58.44553, 58.43916, 58.43248, 
    58.4255, 58.4182, 58.4106, 58.40269, 58.39448, 58.38596, 58.37712, 
    58.36799, 58.35855, 58.3488, 58.33875, 58.32839, 58.31773, 58.30676, 
    58.29549, 58.28392, 58.27204, 58.25986, 58.24737, 58.23458, 58.22149, 
    58.2081, 58.19441, 58.18042, 58.16613, 58.15153, 58.13664, 58.12144, 
    58.10595, 58.09016, 58.07408, 58.05769, 58.04101, 58.02403, 58.00676, 
    57.98919, 57.97132, 57.95316, 57.93471, 57.91596, 57.89692, 57.87759, 
    57.85796, 57.83805, 57.81784, 57.79734, 57.77656, 57.75548, 57.73412, 
    57.71246, 57.69053, 57.6683, 57.64579, 57.62299, 57.59991, 57.57654, 
    57.55289, 57.52895, 57.50474, 57.48024, 57.45546, 57.4304, 57.40506, 
    57.37944, 57.35355, 57.32737, 57.30092, 57.2742, 57.24719, 57.21991, 
    57.19236, 57.16454, 57.13644, 57.10807, 57.07942, 57.05051, 57.02133, 
    56.99187, 56.96215, 56.93217, 56.90191, 56.87139, 56.8406, 56.80955, 
    56.77823, 56.74665, 56.71481, 56.68271, 56.65035, 56.61772, 56.58484, 
    56.5517, 56.5183, 56.48464, 56.45073, 56.41656, 56.38214, 56.34746, 
    56.31253, 56.27735, 56.24192, 56.20624, 56.1703, 56.13412, 56.09769, 
    56.06102, 56.02409, 55.98693, 55.94951, 55.91185, 55.87395, 55.83581, 
    55.79743, 55.7588, 55.71994, 55.68084, 55.64149, 55.60192, 55.5621, 
    55.52205, 55.48177, 55.44125, 55.4005, 55.35951, 55.3183, 55.27685, 
    55.23518, 55.19327, 55.15114, 55.10878, 55.0662, 55.02339, 54.98035, 
    54.9371, 54.89362, 54.84991, 54.80599, 54.76184, 54.71748, 54.6729, 
    54.6281, 54.58308, 54.53785, 54.4924, 54.44675, 54.40087, 54.35479, 
    54.30849, 54.26198,
  49.22952, 49.29216, 49.35466, 49.41702, 49.47924, 49.54132, 49.60326, 
    49.66506, 49.72672, 49.78823, 49.84961, 49.91083, 49.97191, 50.03285, 
    50.09364, 50.15428, 50.21478, 50.27512, 50.33532, 50.39537, 50.45526, 
    50.51501, 50.5746, 50.63404, 50.69333, 50.75246, 50.81144, 50.87026, 
    50.92892, 50.98743, 51.04578, 51.10397, 51.162, 51.21987, 51.27758, 
    51.33513, 51.39251, 51.44973, 51.50679, 51.56368, 51.62041, 51.67697, 
    51.73336, 51.78959, 51.84564, 51.90153, 51.95724, 52.01279, 52.06816, 
    52.12336, 52.17839, 52.23324, 52.28792, 52.34242, 52.39675, 52.45089, 
    52.50486, 52.55865, 52.61226, 52.66569, 52.71894, 52.772, 52.82488, 
    52.87758, 52.93009, 52.98242, 53.03456, 53.08651, 53.13828, 53.18985, 
    53.24123, 53.29243, 53.34343, 53.39425, 53.44486, 53.49529, 53.54551, 
    53.59555, 53.64539, 53.69502, 53.74446, 53.7937, 53.84275, 53.89159, 
    53.94023, 53.98867, 54.0369, 54.08493, 54.13275, 54.18037, 54.22778, 
    54.27499, 54.32198, 54.36877, 54.41534, 54.46171, 54.50786, 54.5538, 
    54.59953, 54.64504, 54.69034, 54.73542, 54.78028, 54.82493, 54.86936, 
    54.91357, 54.95755, 55.00132, 55.04486, 55.08818, 55.13128, 55.17415, 
    55.2168, 55.25922, 55.30141, 55.34337, 55.38511, 55.42661, 55.46788, 
    55.50893, 55.54974, 55.59031, 55.63065, 55.67076, 55.71063, 55.75027, 
    55.78966, 55.82882, 55.86774, 55.90642, 55.94485, 55.98305, 56.021, 
    56.05871, 56.09618, 56.1334, 56.17037, 56.2071, 56.24358, 56.27981, 
    56.31579, 56.35152, 56.387, 56.42223, 56.4572, 56.49193, 56.52639, 
    56.56061, 56.59456, 56.62826, 56.66171, 56.69489, 56.72781, 56.76048, 
    56.79288, 56.82503, 56.85691, 56.88853, 56.91988, 56.95097, 56.98179, 
    57.01235, 57.04264, 57.07267, 57.10242, 57.13191, 57.16113, 57.19007, 
    57.21874, 57.24715, 57.27527, 57.30313, 57.33071, 57.35802, 57.38505, 
    57.4118, 57.43828, 57.46448, 57.4904, 57.51604, 57.5414, 57.56649, 
    57.59129, 57.61581, 57.64005, 57.664, 57.68767, 57.71105, 57.73415, 
    57.75697, 57.7795, 57.80173, 57.82369, 57.84536, 57.86673, 57.88782, 
    57.90862, 57.92912, 57.94934, 57.96926, 57.9889, 58.00824, 58.02728, 
    58.04604, 58.0645, 58.08266, 58.10052, 58.1181, 58.13537, 58.15235, 
    58.16903, 58.18542, 58.2015, 58.21729, 58.23278, 58.24796, 58.26285, 
    58.27744, 58.29173, 58.30571, 58.31939, 58.33278, 58.34585, 58.35863, 
    58.3711, 58.38327, 58.39513, 58.40669, 58.41795, 58.4289, 58.43954, 
    58.44988, 58.45991, 58.46964, 58.47906, 58.48817, 58.49698, 58.50547, 
    58.51366, 58.52155, 58.52912, 58.53639, 58.54335, 58.55, 58.55634, 
    58.56236, 58.56808, 58.5735, 58.5786, 58.58339, 58.58787, 58.59204, 
    58.5959, 58.59945, 58.6027, 58.60563, 58.60824, 58.61055, 58.61255, 
    58.61423, 58.61561, 58.61667, 58.61743, 58.61787, 58.618, 58.61782, 
    58.61733, 58.61652, 58.61541, 58.61399, 58.61225, 58.61021, 58.60785, 
    58.60518, 58.6022, 58.59891, 58.59531, 58.5914, 58.58718, 58.58265, 
    58.57781, 58.57266, 58.5672, 58.56143, 58.55535, 58.54896, 58.54227, 
    58.53526, 58.52795, 58.52032, 58.51239, 58.50415, 58.49561, 58.48675, 
    58.47759, 58.46812, 58.45835, 58.44827, 58.43788, 58.42719, 58.41619, 
    58.40488, 58.39328, 58.38136, 58.36915, 58.35663, 58.3438, 58.33068, 
    58.31725, 58.30352, 58.28949, 58.27515, 58.26052, 58.24558, 58.23035, 
    58.21481, 58.19898, 58.18285, 58.16641, 58.14968, 58.13266, 58.11534, 
    58.09772, 58.0798, 58.06159, 58.04309, 58.02429, 58.0052, 57.98581, 
    57.96613, 57.94616, 57.9259, 57.90535, 57.8845, 57.86337, 57.84195, 
    57.82024, 57.79824, 57.77595, 57.75338, 57.73052, 57.70737, 57.68394, 
    57.66023, 57.63623, 57.61195, 57.58738, 57.56254, 57.53741, 57.512, 
    57.48632, 57.46035, 57.43411, 57.40759, 57.38079, 57.35372, 57.32637, 
    57.29874, 57.27084, 57.24267, 57.21423, 57.18551, 57.15652, 57.12726, 
    57.09773, 57.06794, 57.03787, 57.00753, 56.97694, 56.94607, 56.91494, 
    56.88354, 56.85188, 56.81996, 56.78778, 56.75533, 56.72263, 56.68966, 
    56.65643, 56.62295, 56.58921, 56.55521, 56.52096, 56.48645, 56.45169, 
    56.41667, 56.3814, 56.34589, 56.31012, 56.27409, 56.23782, 56.20131, 
    56.16454, 56.12753, 56.09027, 56.05276, 56.01502, 55.97702, 55.93879, 
    55.90031, 55.8616, 55.82264, 55.78345, 55.74401, 55.70434, 55.66443, 
    55.62429, 55.58391, 55.5433, 55.50245, 55.46137, 55.42006, 55.37852, 
    55.33675, 55.29475, 55.25252, 55.21006, 55.16739, 55.12448, 55.08134, 
    55.03799, 54.99441, 54.95061, 54.90659, 54.86235, 54.81788, 54.7732, 
    54.72831, 54.68319, 54.63786, 54.59231, 54.54655, 54.50058, 54.45439, 
    54.40799, 54.36138,
  49.31944, 49.38218, 49.44477, 49.50723, 49.56955, 49.63173, 49.69377, 
    49.75567, 49.81742, 49.87904, 49.94051, 50.00183, 50.06301, 50.12405, 
    50.18494, 50.24568, 50.30628, 50.36672, 50.42702, 50.48717, 50.54716, 
    50.60701, 50.66671, 50.72625, 50.78563, 50.84486, 50.90394, 50.96287, 
    51.02163, 51.08024, 51.13869, 51.19698, 51.25512, 51.31309, 51.3709, 
    51.42855, 51.48603, 51.54336, 51.60052, 51.65751, 51.71434, 51.771, 
    51.8275, 51.88383, 51.93999, 51.99598, 52.0518, 52.10744, 52.16292, 
    52.21822, 52.27335, 52.32831, 52.38309, 52.43769, 52.49212, 52.54637, 
    52.60044, 52.65433, 52.70805, 52.76158, 52.81493, 52.86809, 52.92108, 
    52.97388, 53.02649, 53.07892, 53.13116, 53.18322, 53.23509, 53.28677, 
    53.33826, 53.38955, 53.44066, 53.49157, 53.54229, 53.59282, 53.64315, 
    53.69329, 53.74323, 53.79297, 53.84251, 53.89185, 53.941, 53.98994, 
    54.03868, 54.08722, 54.13556, 54.18369, 54.23161, 54.27934, 54.32685, 
    54.37415, 54.42125, 54.46814, 54.51481, 54.56128, 54.60753, 54.65357, 
    54.6994, 54.74501, 54.79041, 54.83559, 54.88055, 54.9253, 54.96983, 
    55.01413, 55.05822, 55.10208, 55.14572, 55.18914, 55.23233, 55.2753, 
    55.31805, 55.36056, 55.40285, 55.44491, 55.48674, 55.52834, 55.56971, 
    55.61085, 55.65176, 55.69243, 55.73286, 55.77306, 55.81303, 55.85276, 
    55.89225, 55.9315, 55.97051, 56.00928, 56.04781, 56.0861, 56.12414, 
    56.16194, 56.1995, 56.23681, 56.27387, 56.31069, 56.34726, 56.38358, 
    56.41965, 56.45547, 56.49103, 56.52635, 56.56141, 56.59622, 56.63077, 
    56.66507, 56.69911, 56.7329, 56.76642, 56.79969, 56.8327, 56.86545, 
    56.89793, 56.93016, 56.96212, 56.99382, 57.02525, 57.05642, 57.08733, 
    57.11797, 57.14833, 57.17844, 57.20827, 57.23783, 57.26712, 57.29614, 
    57.32489, 57.35337, 57.38157, 57.4095, 57.43716, 57.46453, 57.49163, 
    57.51846, 57.54501, 57.57128, 57.59727, 57.62298, 57.64841, 57.67356, 
    57.69843, 57.72301, 57.74731, 57.77133, 57.79506, 57.81851, 57.84167, 
    57.86455, 57.88714, 57.90944, 57.93146, 57.95318, 57.97462, 57.99576, 
    58.01662, 58.03718, 58.05745, 58.07743, 58.09712, 58.11651, 58.13561, 
    58.15442, 58.17292, 58.19114, 58.20906, 58.22668, 58.244, 58.26103, 
    58.27776, 58.29419, 58.31031, 58.32615, 58.34168, 58.35691, 58.37184, 
    58.38647, 58.40079, 58.41482, 58.42854, 58.44196, 58.45507, 58.46788, 
    58.48039, 58.4926, 58.50449, 58.51609, 58.52737, 58.53835, 58.54903, 
    58.55939, 58.56946, 58.57921, 58.58866, 58.5978, 58.60663, 58.61515, 
    58.62336, 58.63127, 58.63887, 58.64615, 58.65313, 58.6598, 58.66616, 
    58.6722, 58.67794, 58.68337, 58.68848, 58.69329, 58.69778, 58.70197, 
    58.70584, 58.7094, 58.71265, 58.71559, 58.71822, 58.72053, 58.72253, 
    58.72422, 58.7256, 58.72667, 58.72742, 58.72787, 58.728, 58.72782, 
    58.72733, 58.72652, 58.7254, 58.72398, 58.72224, 58.72018, 58.71782, 
    58.71515, 58.71216, 58.70886, 58.70525, 58.70132, 58.69709, 58.69255, 
    58.68769, 58.68253, 58.67706, 58.67127, 58.66517, 58.65876, 58.65205, 
    58.64502, 58.63768, 58.63004, 58.62209, 58.61382, 58.60525, 58.59637, 
    58.58718, 58.57769, 58.56789, 58.55778, 58.54736, 58.53664, 58.52561, 
    58.51427, 58.50263, 58.49068, 58.47844, 58.46588, 58.45302, 58.43985, 
    58.42639, 58.41262, 58.39855, 58.38417, 58.3695, 58.35452, 58.33924, 
    58.32366, 58.30779, 58.29161, 58.27513, 58.25835, 58.24128, 58.22391, 
    58.20624, 58.18828, 58.17002, 58.15146, 58.13261, 58.11346, 58.09402, 
    58.07429, 58.05426, 58.03395, 58.01334, 57.99244, 57.97124, 57.94976, 
    57.92799, 57.90593, 57.88359, 57.86095, 57.83803, 57.81482, 57.79133, 
    57.76755, 57.74349, 57.71914, 57.69451, 57.6696, 57.64441, 57.61893, 
    57.59318, 57.56714, 57.54083, 57.51424, 57.48737, 57.46022, 57.4328, 
    57.4051, 57.37713, 57.34888, 57.32036, 57.29157, 57.2625, 57.23317, 
    57.20357, 57.17369, 57.14355, 57.11314, 57.08245, 57.05151, 57.0203, 
    56.98882, 56.95708, 56.92508, 56.89281, 56.86029, 56.8275, 56.79445, 
    56.76114, 56.72757, 56.69374, 56.65966, 56.62532, 56.59073, 56.55588, 
    56.52078, 56.48542, 56.44982, 56.41396, 56.37785, 56.34149, 56.30488, 
    56.26803, 56.23092, 56.19357, 56.15598, 56.11814, 56.08006, 56.04173, 
    56.00317, 55.96436, 55.9253, 55.88602, 55.84649, 55.80672, 55.76672, 
    55.72648, 55.68601, 55.6453, 55.60436, 55.56318, 55.52178, 55.48014, 
    55.43827, 55.39618, 55.35385, 55.3113, 55.26852, 55.22552, 55.18229, 
    55.13883, 55.09516, 55.05126, 55.00714, 54.9628, 54.91824, 54.87346, 
    54.82846, 54.78324, 54.73781, 54.69217, 54.64631, 54.60023, 54.55394, 
    54.50744, 54.46074,
  49.40928, 49.47211, 49.53481, 49.59737, 49.65978, 49.72206, 49.7842, 
    49.8462, 49.90805, 49.96976, 50.03133, 50.09276, 50.15404, 50.21518, 
    50.27616, 50.33701, 50.3977, 50.45825, 50.51865, 50.57889, 50.63899, 
    50.69894, 50.75873, 50.81837, 50.87786, 50.93719, 50.99638, 51.0554, 
    51.11427, 51.17298, 51.23153, 51.28992, 51.34816, 51.40623, 51.46415, 
    51.5219, 51.57949, 51.63691, 51.69418, 51.75127, 51.8082, 51.86497, 
    51.92157, 51.978, 52.03426, 52.09035, 52.14627, 52.20202, 52.2576, 
    52.31301, 52.36824, 52.4233, 52.47818, 52.53289, 52.58742, 52.64177, 
    52.69595, 52.74995, 52.80376, 52.8574, 52.91085, 52.96412, 53.01721, 
    53.07011, 53.12283, 53.17536, 53.22771, 53.27987, 53.33184, 53.38362, 
    53.43521, 53.48661, 53.53782, 53.58884, 53.63966, 53.69029, 53.74073, 
    53.79097, 53.84101, 53.89085, 53.9405, 53.98994, 54.03919, 54.08824, 
    54.13708, 54.18572, 54.23416, 54.28239, 54.33042, 54.37824, 54.42586, 
    54.47326, 54.52046, 54.56745, 54.61423, 54.66079, 54.70715, 54.75329, 
    54.79922, 54.84493, 54.89043, 54.93571, 54.98077, 55.02562, 55.07024, 
    55.11465, 55.15883, 55.20279, 55.24653, 55.29005, 55.33334, 55.37641, 
    55.41925, 55.46186, 55.50425, 55.54641, 55.58834, 55.63003, 55.6715, 
    55.71273, 55.75373, 55.7945, 55.83503, 55.87533, 55.91539, 55.95521, 
    55.99479, 56.03414, 56.07324, 56.11211, 56.15073, 56.18911, 56.22724, 
    56.26514, 56.30278, 56.34018, 56.37734, 56.41424, 56.4509, 56.48731, 
    56.52347, 56.55938, 56.59503, 56.63044, 56.66558, 56.70048, 56.73512, 
    56.7695, 56.80363, 56.8375, 56.87111, 56.90446, 56.93756, 56.97039, 
    57.00296, 57.03526, 57.06731, 57.09909, 57.1306, 57.16185, 57.19283, 
    57.22355, 57.254, 57.28418, 57.31409, 57.34373, 57.3731, 57.40219, 
    57.43102, 57.45957, 57.48785, 57.51585, 57.54358, 57.57103, 57.5982, 
    57.6251, 57.65172, 57.67806, 57.70412, 57.7299, 57.75539, 57.78061, 
    57.80555, 57.8302, 57.85456, 57.87865, 57.90245, 57.92596, 57.94918, 
    57.97212, 57.99477, 58.01714, 58.03921, 58.06099, 58.08249, 58.10369, 
    58.1246, 58.14523, 58.16555, 58.18559, 58.20533, 58.22477, 58.24393, 
    58.26278, 58.28135, 58.29961, 58.31758, 58.33525, 58.35262, 58.36969, 
    58.38647, 58.40295, 58.41912, 58.435, 58.45057, 58.46585, 58.48082, 
    58.49549, 58.50985, 58.52392, 58.53768, 58.55114, 58.56429, 58.57714, 
    58.58968, 58.60192, 58.61385, 58.62548, 58.6368, 58.64781, 58.65851, 
    58.66891, 58.679, 58.68878, 58.69826, 58.70742, 58.71628, 58.72483, 
    58.73306, 58.74099, 58.74861, 58.75592, 58.76291, 58.7696, 58.77598, 
    58.78204, 58.7878, 58.79324, 58.79837, 58.80319, 58.8077, 58.81189, 
    58.81578, 58.81935, 58.82261, 58.82555, 58.82819, 58.83051, 58.83252, 
    58.83421, 58.83559, 58.83667, 58.83742, 58.83787, 58.838, 58.83782, 
    58.83732, 58.83652, 58.8354, 58.83397, 58.83222, 58.83016, 58.82779, 
    58.82511, 58.82211, 58.8188, 58.81518, 58.81125, 58.807, 58.80245, 
    58.79758, 58.7924, 58.78691, 58.78111, 58.77499, 58.76856, 58.76183, 
    58.75478, 58.74743, 58.73976, 58.73178, 58.7235, 58.7149, 58.70599, 
    58.69678, 58.68726, 58.67743, 58.66729, 58.65684, 58.64608, 58.63503, 
    58.62366, 58.61198, 58.6, 58.58772, 58.57513, 58.56223, 58.54903, 
    58.53552, 58.52171, 58.5076, 58.49319, 58.47847, 58.46345, 58.44813, 
    58.43251, 58.41658, 58.40036, 58.38383, 58.36702, 58.34989, 58.33247, 
    58.31475, 58.29674, 58.27843, 58.25982, 58.24092, 58.22172, 58.20222, 
    58.18244, 58.16236, 58.14198, 58.12132, 58.10036, 58.07911, 58.05757, 
    58.03574, 58.01362, 57.99121, 57.96851, 57.94553, 57.92226, 57.8987, 
    57.87486, 57.85073, 57.82632, 57.80162, 57.77664, 57.75138, 57.72584, 
    57.70002, 57.67391, 57.64753, 57.62086, 57.59392, 57.5667, 57.53921, 
    57.51144, 57.48339, 57.45507, 57.42648, 57.39761, 57.36847, 57.33906, 
    57.30938, 57.27942, 57.2492, 57.21871, 57.18795, 57.15693, 57.12563, 
    57.09408, 57.06226, 57.03017, 56.99782, 56.96521, 56.93234, 56.8992, 
    56.86581, 56.83216, 56.79825, 56.76408, 56.72966, 56.69498, 56.66004, 
    56.62485, 56.58941, 56.55371, 56.51777, 56.48157, 56.44512, 56.40842, 
    56.37148, 56.33428, 56.29684, 56.25916, 56.22123, 56.18305, 56.14463, 
    56.10597, 56.06707, 56.02793, 55.98855, 55.94893, 55.90907, 55.86897, 
    55.82864, 55.78807, 55.74726, 55.70623, 55.66496, 55.62345, 55.58172, 
    55.53975, 55.49756, 55.45514, 55.41249, 55.36961, 55.32651, 55.28318, 
    55.23963, 55.19585, 55.15186, 55.10764, 55.0632, 55.01854, 54.97366, 
    54.92856, 54.88324, 54.83772, 54.79197, 54.74601, 54.69983, 54.65344, 
    54.60684, 54.56003,
  49.49903, 49.56197, 49.62476, 49.68742, 49.74993, 49.81231, 49.87455, 
    49.93664, 49.9986, 50.06041, 50.12208, 50.1836, 50.24498, 50.30622, 
    50.36731, 50.42825, 50.48904, 50.54969, 50.61019, 50.67054, 50.73074, 
    50.79078, 50.85068, 50.91042, 50.97001, 51.02945, 51.08873, 51.14785, 
    51.20683, 51.26564, 51.32429, 51.38279, 51.44112, 51.4993, 51.55732, 
    51.61517, 51.67286, 51.73039, 51.78776, 51.84496, 51.90199, 51.95886, 
    52.01556, 52.07209, 52.12846, 52.18465, 52.24068, 52.29654, 52.35221, 
    52.40773, 52.46306, 52.51822, 52.57321, 52.62802, 52.68266, 52.73711, 
    52.79139, 52.84549, 52.89941, 52.95315, 53.00671, 53.06008, 53.11327, 
    53.16628, 53.2191, 53.27174, 53.32419, 53.37645, 53.42852, 53.48041, 
    53.5321, 53.58361, 53.63492, 53.68604, 53.73697, 53.7877, 53.83824, 
    53.88858, 53.93873, 53.98867, 54.03843, 54.08797, 54.13733, 54.18647, 
    54.23542, 54.28416, 54.3327, 54.38104, 54.42917, 54.47709, 54.52481, 
    54.57232, 54.61962, 54.66671, 54.71358, 54.76025, 54.80671, 54.85295, 
    54.89898, 54.94479, 54.99039, 55.03577, 55.08094, 55.12588, 55.1706, 
    55.21511, 55.2594, 55.30346, 55.3473, 55.39091, 55.4343, 55.47747, 
    55.52041, 55.56312, 55.6056, 55.64786, 55.68988, 55.73168, 55.77324, 
    55.81457, 55.85566, 55.89653, 55.93715, 55.97755, 56.0177, 56.05762, 
    56.09729, 56.13673, 56.17593, 56.21489, 56.2536, 56.29208, 56.33031, 
    56.36829, 56.40603, 56.44352, 56.48077, 56.51776, 56.55451, 56.59101, 
    56.62725, 56.66325, 56.699, 56.73449, 56.76973, 56.80471, 56.83943, 
    56.87391, 56.90812, 56.94207, 56.97577, 57.0092, 57.04238, 57.07529, 
    57.10795, 57.14034, 57.17247, 57.20433, 57.23592, 57.26725, 57.29832, 
    57.32911, 57.35964, 57.3899, 57.41988, 57.4496, 57.47905, 57.50822, 
    57.53712, 57.56575, 57.5941, 57.62218, 57.64998, 57.6775, 57.70475, 
    57.73172, 57.75841, 57.78482, 57.81095, 57.8368, 57.86236, 57.88765, 
    57.91265, 57.93737, 57.9618, 57.98595, 58.00981, 58.03339, 58.05668, 
    58.07968, 58.10239, 58.12482, 58.14695, 58.16879, 58.19035, 58.21161, 
    58.23258, 58.25326, 58.27364, 58.29373, 58.31353, 58.33303, 58.35223, 
    58.37114, 58.38976, 58.40807, 58.42609, 58.44381, 58.46123, 58.47836, 
    58.49518, 58.5117, 58.52792, 58.54384, 58.55946, 58.57478, 58.58979, 
    58.6045, 58.61891, 58.63301, 58.64682, 58.66031, 58.6735, 58.68639, 
    58.69896, 58.71124, 58.7232, 58.73486, 58.74621, 58.75726, 58.76799, 
    58.77842, 58.78854, 58.79835, 58.80785, 58.81704, 58.82592, 58.8345, 
    58.84276, 58.85071, 58.85835, 58.86568, 58.8727, 58.8794, 58.8858, 
    58.89188, 58.89765, 58.90311, 58.90825, 58.91309, 58.91761, 58.92182, 
    58.92571, 58.92929, 58.93256, 58.93552, 58.93816, 58.94049, 58.9425, 
    58.9442, 58.94559, 58.94666, 58.94742, 58.94787, 58.948, 58.94782, 
    58.94732, 58.94651, 58.94539, 58.94395, 58.9422, 58.94014, 58.93776, 
    58.93507, 58.93206, 58.92875, 58.92511, 58.92117, 58.91691, 58.91234, 
    58.90746, 58.90227, 58.89676, 58.89094, 58.88481, 58.87836, 58.8716, 
    58.86454, 58.85716, 58.84947, 58.84147, 58.83316, 58.82454, 58.81561, 
    58.80637, 58.79682, 58.78696, 58.77679, 58.76632, 58.75553, 58.74444, 
    58.73304, 58.72133, 58.70932, 58.69699, 58.68437, 58.67143, 58.6582, 
    58.64465, 58.6308, 58.61665, 58.6022, 58.58744, 58.57237, 58.55701, 
    58.54134, 58.52538, 58.50911, 58.49253, 58.47567, 58.4585, 58.44103, 
    58.42326, 58.4052, 58.38683, 58.36817, 58.34922, 58.32996, 58.31042, 
    58.29057, 58.27044, 58.25001, 58.22928, 58.20827, 58.18696, 58.16536, 
    58.14347, 58.12129, 58.09882, 58.07606, 58.05301, 58.02968, 58.00606, 
    57.98215, 57.95795, 57.93348, 57.90871, 57.88367, 57.85834, 57.83273, 
    57.80683, 57.78066, 57.7542, 57.72747, 57.70046, 57.67317, 57.6456, 
    57.61776, 57.58963, 57.56124, 57.53257, 57.50362, 57.47441, 57.44492, 
    57.41516, 57.38513, 57.35483, 57.32426, 57.29342, 57.26231, 57.23094, 
    57.1993, 57.1674, 57.13523, 57.1028, 57.07011, 57.03715, 57.00393, 
    56.97046, 56.93672, 56.90272, 56.86847, 56.83396, 56.79919, 56.76417, 
    56.72889, 56.69336, 56.65757, 56.62154, 56.58525, 56.54871, 56.51192, 
    56.47489, 56.43761, 56.40007, 56.3623, 56.32428, 56.28601, 56.2475, 
    56.20874, 56.16975, 56.13051, 56.09103, 56.05132, 56.01136, 55.97117, 
    55.93074, 55.89008, 55.84918, 55.80805, 55.76668, 55.72508, 55.68325, 
    55.64119, 55.5989, 55.55638, 55.51363, 55.47065, 55.42746, 55.38403, 
    55.34038, 55.2965, 55.25241, 55.20809, 55.16355, 55.11879, 55.07381, 
    55.02861, 54.98319, 54.93756, 54.89172, 54.84565, 54.79938, 54.75289, 
    54.70618, 54.65927,
  49.58871, 49.65174, 49.71463, 49.77738, 49.84, 49.90247, 49.96481, 50.027, 
    50.08906, 50.15097, 50.21274, 50.27436, 50.33584, 50.39718, 50.45837, 
    50.51941, 50.58031, 50.64106, 50.70166, 50.7621, 50.8224, 50.88255, 
    50.94255, 51.0024, 51.06208, 51.12162, 51.18101, 51.24023, 51.2993, 
    51.35822, 51.41698, 51.47557, 51.53402, 51.59229, 51.65041, 51.70837, 
    51.76616, 51.8238, 51.88126, 51.93857, 51.9957, 52.05268, 52.10948, 
    52.16612, 52.22259, 52.27888, 52.33501, 52.39097, 52.44676, 52.50237, 
    52.55781, 52.61308, 52.66817, 52.72308, 52.77782, 52.83238, 52.88676, 
    52.94097, 52.99499, 53.04884, 53.1025, 53.15598, 53.20927, 53.26238, 
    53.31531, 53.36805, 53.4206, 53.47297, 53.52515, 53.57714, 53.62894, 
    53.68055, 53.73196, 53.78318, 53.83422, 53.88505, 53.93569, 53.98614, 
    54.03639, 54.08644, 54.13629, 54.18594, 54.2354, 54.28465, 54.3337, 
    54.38255, 54.43119, 54.47963, 54.52786, 54.57589, 54.6237, 54.67131, 
    54.71872, 54.76591, 54.81289, 54.85966, 54.90622, 54.95256, 54.99869, 
    55.04461, 55.09031, 55.13578, 55.18105, 55.22609, 55.27092, 55.31553, 
    55.35991, 55.40407, 55.44801, 55.49173, 55.53521, 55.57848, 55.62152, 
    55.66433, 55.70691, 55.74926, 55.79138, 55.83327, 55.87494, 55.91636, 
    55.95755, 55.99851, 56.03923, 56.07972, 56.11997, 56.15998, 56.19976, 
    56.23929, 56.27858, 56.31763, 56.35644, 56.39501, 56.43333, 56.47141, 
    56.50924, 56.54682, 56.58416, 56.62124, 56.65808, 56.69467, 56.73101, 
    56.76709, 56.80293, 56.8385, 56.87383, 56.9089, 56.94371, 56.97827, 
    57.01257, 57.04661, 57.08039, 57.11392, 57.14718, 57.18018, 57.21291, 
    57.24538, 57.2776, 57.30954, 57.34122, 57.37263, 57.40377, 57.43465, 
    57.46525, 57.49559, 57.52566, 57.55545, 57.58498, 57.61422, 57.6432, 
    57.67191, 57.70033, 57.72848, 57.75636, 57.78395, 57.81128, 57.83831, 
    57.86508, 57.89156, 57.91776, 57.94368, 57.96931, 57.99467, 58.01973, 
    58.04452, 58.06902, 58.09324, 58.11716, 58.1408, 58.16415, 58.18722, 
    58.21, 58.23248, 58.25468, 58.27658, 58.29819, 58.31952, 58.34054, 
    58.36128, 58.38172, 58.40186, 58.42171, 58.44127, 58.46053, 58.47949, 
    58.49816, 58.51653, 58.5346, 58.55236, 58.56984, 58.58701, 58.60387, 
    58.62045, 58.63671, 58.65268, 58.66834, 58.6837, 58.69876, 58.71351, 
    58.72796, 58.7421, 58.75594, 58.76948, 58.78271, 58.79563, 58.80824, 
    58.82055, 58.83255, 58.84424, 58.85563, 58.8667, 58.87747, 58.88793, 
    58.89808, 58.90792, 58.91745, 58.92666, 58.93557, 58.94417, 58.95245, 
    58.96043, 58.96809, 58.97544, 58.98248, 58.9892, 58.99562, 59.00172, 
    59.0075, 59.01298, 59.01814, 59.02299, 59.02752, 59.03174, 59.03564, 
    59.03924, 59.04251, 59.04548, 59.04813, 59.05046, 59.05248, 59.05419, 
    59.05558, 59.05666, 59.05742, 59.05787, 59.058, 59.05782, 59.05732, 
    59.05651, 59.05538, 59.05394, 59.05219, 59.05011, 59.04773, 59.04503, 
    59.04202, 59.03869, 59.03505, 59.03109, 59.02682, 59.02224, 59.01734, 
    59.01213, 59.00661, 59.00077, 58.99462, 58.98816, 58.98138, 58.9743, 
    58.9669, 58.95919, 58.95116, 58.94283, 58.93418, 58.92522, 58.91596, 
    58.90638, 58.89649, 58.8863, 58.87579, 58.86497, 58.85385, 58.84241, 
    58.83067, 58.81862, 58.80627, 58.7936, 58.78063, 58.76736, 58.75378, 
    58.73989, 58.7257, 58.7112, 58.6964, 58.68129, 58.66588, 58.65017, 
    58.63416, 58.61784, 58.60123, 58.58431, 58.56709, 58.54957, 58.53176, 
    58.51364, 58.49522, 58.47651, 58.4575, 58.4382, 58.41859, 58.3987, 
    58.37851, 58.35802, 58.33723, 58.31616, 58.2948, 58.27314, 58.25119, 
    58.22894, 58.20641, 58.18359, 58.16048, 58.13708, 58.1134, 58.08942, 
    58.06516, 58.04062, 58.01579, 57.99067, 57.96527, 57.93959, 57.91363, 
    57.88739, 57.86086, 57.83406, 57.80697, 57.77961, 57.75197, 57.72405, 
    57.69585, 57.66738, 57.63864, 57.60962, 57.58032, 57.55076, 57.52092, 
    57.49081, 57.46043, 57.42978, 57.39886, 57.36768, 57.33622, 57.3045, 
    57.27252, 57.24026, 57.20775, 57.17497, 57.14193, 57.10863, 57.07507, 
    57.04124, 57.00716, 56.97282, 56.93822, 56.90337, 56.86826, 56.83289, 
    56.79728, 56.7614, 56.72528, 56.6889, 56.65227, 56.61539, 56.57827, 
    56.54089, 56.50327, 56.4654, 56.42728, 56.38892, 56.35032, 56.31147, 
    56.27238, 56.23305, 56.19348, 56.15367, 56.11362, 56.07333, 56.03281, 
    55.99205, 55.95105, 55.90982, 55.86836, 55.82666, 55.78474, 55.74258, 
    55.70019, 55.65757, 55.61472, 55.57165, 55.52835, 55.48483, 55.44107, 
    55.3971, 55.35291, 55.30848, 55.26384, 55.21898, 55.1739, 55.1286, 
    55.08309, 55.03736, 54.99141, 54.94524, 54.89887, 54.85228, 54.80547, 
    54.75846,
  49.6783, 49.74142, 49.80442, 49.86727, 49.92998, 49.99256, 50.05499, 
    50.11729, 50.17944, 50.24145, 50.30332, 50.36504, 50.42662, 50.48806, 
    50.54935, 50.6105, 50.67149, 50.73234, 50.79304, 50.85359, 50.91399, 
    50.97424, 51.03434, 51.09429, 51.15408, 51.21372, 51.2732, 51.33253, 
    51.39171, 51.45073, 51.50959, 51.56829, 51.62683, 51.68521, 51.74343, 
    51.80149, 51.85939, 51.91713, 51.9747, 52.0321, 52.08934, 52.14642, 
    52.20333, 52.26007, 52.31664, 52.37304, 52.42928, 52.48534, 52.54123, 
    52.59695, 52.65249, 52.70786, 52.76305, 52.81807, 52.87292, 52.92758, 
    52.98207, 53.03638, 53.0905, 53.14445, 53.19822, 53.2518, 53.3052, 
    53.35841, 53.41145, 53.46429, 53.51695, 53.56942, 53.6217, 53.6738, 
    53.7257, 53.77741, 53.82893, 53.88026, 53.9314, 53.98234, 54.03308, 
    54.08363, 54.13398, 54.18414, 54.2341, 54.28385, 54.33341, 54.38276, 
    54.43192, 54.48087, 54.52961, 54.57816, 54.62649, 54.67462, 54.72254, 
    54.77026, 54.81776, 54.86506, 54.91214, 54.95901, 55.00567, 55.05212, 
    55.09835, 55.14436, 55.19016, 55.23575, 55.28111, 55.32626, 55.37119, 
    55.41589, 55.46037, 55.50463, 55.54868, 55.59249, 55.63608, 55.67944, 
    55.72258, 55.76549, 55.80817, 55.85062, 55.89284, 55.93483, 55.97659, 
    56.01811, 56.0594, 56.10045, 56.14127, 56.18185, 56.2222, 56.26231, 
    56.30218, 56.3418, 56.38119, 56.42034, 56.45924, 56.4979, 56.53631, 
    56.57448, 56.6124, 56.65008, 56.68751, 56.72469, 56.76162, 56.79829, 
    56.83472, 56.8709, 56.90682, 56.94249, 56.97791, 57.01306, 57.04796, 
    57.08261, 57.11699, 57.15112, 57.18499, 57.2186, 57.25194, 57.28503, 
    57.31785, 57.3504, 57.38269, 57.41472, 57.44648, 57.47797, 57.5092, 
    57.54015, 57.57084, 57.60126, 57.6314, 57.66128, 57.69088, 57.72021, 
    57.74926, 57.77804, 57.80654, 57.83477, 57.86272, 57.89039, 57.91778, 
    57.94489, 57.97173, 57.99828, 58.02455, 58.05054, 58.07624, 58.10167, 
    58.1268, 58.15165, 58.17622, 58.2005, 58.22449, 58.2482, 58.27162, 
    58.29475, 58.31758, 58.34013, 58.36239, 58.38435, 58.40602, 58.42741, 
    58.44849, 58.46928, 58.48978, 58.50999, 58.52989, 58.5495, 58.56882, 
    58.58783, 58.60655, 58.62497, 58.64309, 58.66091, 58.67843, 58.69565, 
    58.71257, 58.72918, 58.74549, 58.76151, 58.77721, 58.79262, 58.80772, 
    58.82251, 58.83701, 58.85119, 58.86507, 58.87864, 58.89191, 58.90487, 
    58.91752, 58.92986, 58.94189, 58.95362, 58.96504, 58.97615, 58.98695, 
    58.99743, 59.00761, 59.01748, 59.02703, 59.03628, 59.04521, 59.05383, 
    59.06215, 59.07014, 59.07782, 59.0852, 59.09225, 59.099, 59.10543, 
    59.11155, 59.11736, 59.12284, 59.12802, 59.13288, 59.13743, 59.14166, 
    59.14558, 59.14918, 59.15247, 59.15544, 59.1581, 59.16044, 59.16247, 
    59.16418, 59.16557, 59.16665, 59.16742, 59.16787, 59.168, 59.16782, 
    59.16732, 59.1665, 59.16537, 59.16393, 59.16217, 59.16009, 59.1577, 
    59.15499, 59.15197, 59.14863, 59.14498, 59.14101, 59.13673, 59.13213, 
    59.12722, 59.122, 59.11646, 59.1106, 59.10443, 59.09795, 59.09116, 
    59.08405, 59.07663, 59.0689, 59.06085, 59.05249, 59.04382, 59.03484, 
    59.02554, 59.01594, 59.00602, 58.9958, 58.98526, 58.97441, 58.96325, 
    58.95179, 58.94001, 58.92793, 58.91553, 58.90284, 58.88983, 58.87651, 
    58.86289, 58.84896, 58.83473, 58.82019, 58.80535, 58.7902, 58.77475, 
    58.759, 58.74294, 58.72657, 58.70991, 58.69294, 58.67568, 58.65811, 
    58.64024, 58.62207, 58.60361, 58.58484, 58.56578, 58.54642, 58.52676, 
    58.50681, 58.48656, 58.46601, 58.44518, 58.42405, 58.40262, 58.3809, 
    58.35889, 58.33659, 58.31399, 58.29111, 58.26793, 58.24447, 58.22072, 
    58.19668, 58.17236, 58.14774, 58.12284, 58.09766, 58.0722, 58.04644, 
    58.02041, 57.9941, 57.9675, 57.94062, 57.91346, 57.88603, 57.85831, 
    57.83032, 57.80205, 57.7735, 57.74468, 57.71558, 57.68621, 57.65657, 
    57.62665, 57.59647, 57.56601, 57.53527, 57.50428, 57.47301, 57.44147, 
    57.40967, 57.37761, 57.34527, 57.31267, 57.27981, 57.24669, 57.2133, 
    57.17965, 57.14574, 57.11157, 57.07714, 57.04246, 57.00752, 56.97232, 
    56.93687, 56.90116, 56.86519, 56.82898, 56.79251, 56.75579, 56.71882, 
    56.6816, 56.64414, 56.60642, 56.56846, 56.53025, 56.4918, 56.4531, 
    56.41416, 56.37498, 56.33555, 56.29589, 56.25598, 56.21584, 56.17545, 
    56.13483, 56.09398, 56.05288, 56.01155, 55.96999, 55.9282, 55.88617, 
    55.84392, 55.80143, 55.75871, 55.71577, 55.6726, 55.6292, 55.58557, 
    55.54172, 55.49765, 55.45335, 55.40883, 55.36409, 55.31913, 55.27395, 
    55.22855, 55.18293, 55.1371, 55.09105, 55.04478, 54.9983, 54.95161, 
    54.90471, 54.85759,
  49.7678, 49.83103, 49.89412, 49.95707, 50.01988, 50.08256, 50.14509, 
    50.20749, 50.26974, 50.33185, 50.39382, 50.45564, 50.51733, 50.57886, 
    50.64025, 50.7015, 50.7626, 50.82354, 50.88435, 50.945, 51.0055, 
    51.06585, 51.12605, 51.1861, 51.246, 51.30574, 51.36533, 51.42476, 
    51.48404, 51.54316, 51.60212, 51.66092, 51.71957, 51.77805, 51.83638, 
    51.89454, 51.95254, 52.01038, 52.06805, 52.12556, 52.18291, 52.24009, 
    52.2971, 52.35394, 52.41062, 52.46713, 52.52346, 52.57963, 52.63562, 
    52.69145, 52.7471, 52.80257, 52.85787, 52.91299, 52.96794, 53.02271, 
    53.0773, 53.13171, 53.18595, 53.24, 53.29387, 53.34756, 53.40106, 
    53.45438, 53.50752, 53.56047, 53.61323, 53.66581, 53.71819, 53.77039, 
    53.8224, 53.87422, 53.92584, 53.97728, 54.02851, 54.07956, 54.13041, 
    54.18106, 54.23152, 54.28178, 54.33184, 54.3817, 54.43136, 54.48082, 
    54.53008, 54.57913, 54.62798, 54.67662, 54.72506, 54.7733, 54.82132, 
    54.86914, 54.91675, 54.96415, 55.01133, 55.05831, 55.10507, 55.15162, 
    55.19795, 55.24407, 55.28997, 55.33566, 55.38112, 55.42637, 55.47139, 
    55.5162, 55.56079, 55.60515, 55.64929, 55.6932, 55.73689, 55.78035, 
    55.82359, 55.8666, 55.90938, 55.95193, 55.99425, 56.03633, 56.07819, 
    56.11981, 56.1612, 56.20235, 56.24327, 56.28395, 56.32439, 56.36459, 
    56.40455, 56.44428, 56.48376, 56.523, 56.562, 56.60075, 56.63926, 
    56.67752, 56.71553, 56.7533, 56.79082, 56.82809, 56.86512, 56.90189, 
    56.9384, 56.97467, 57.01068, 57.04644, 57.08194, 57.11719, 57.15218, 
    57.18691, 57.22139, 57.2556, 57.28955, 57.32325, 57.35668, 57.38985, 
    57.42275, 57.45539, 57.48777, 57.51987, 57.55172, 57.58329, 57.6146, 
    57.64564, 57.6764, 57.7069, 57.73713, 57.76708, 57.79676, 57.82616, 
    57.85529, 57.88415, 57.91273, 57.94103, 57.96905, 57.9968, 58.02426, 
    58.05145, 58.07835, 58.10498, 58.13132, 58.15738, 58.18316, 58.20864, 
    58.23385, 58.25877, 58.28341, 58.30775, 58.33181, 58.35558, 58.37906, 
    58.40226, 58.42516, 58.44777, 58.47009, 58.49211, 58.51385, 58.53529, 
    58.55643, 58.57728, 58.59784, 58.6181, 58.63806, 58.65772, 58.67709, 
    58.69616, 58.71493, 58.7334, 58.75158, 58.76944, 58.78701, 58.80428, 
    58.82125, 58.83791, 58.85427, 58.87033, 58.88608, 58.90153, 58.91667, 
    58.93151, 58.94604, 58.96027, 58.97419, 58.9878, 59.0011, 59.0141, 
    59.02679, 59.03917, 59.05124, 59.063, 59.07445, 59.08559, 59.09642, 
    59.10693, 59.11714, 59.12704, 59.13662, 59.14589, 59.15485, 59.1635, 
    59.17183, 59.17986, 59.18756, 59.19495, 59.20203, 59.2088, 59.21525, 
    59.22139, 59.22721, 59.23271, 59.2379, 59.24278, 59.24734, 59.25159, 
    59.25552, 59.25913, 59.26242, 59.2654, 59.26807, 59.27042, 59.27245, 
    59.27417, 59.27557, 59.27665, 59.27742, 59.27787, 59.278, 59.27782, 
    59.27732, 59.2765, 59.27537, 59.27392, 59.27215, 59.27007, 59.26767, 
    59.26495, 59.26192, 59.25858, 59.25491, 59.25093, 59.24664, 59.24203, 
    59.2371, 59.23186, 59.22631, 59.22044, 59.21425, 59.20775, 59.20094, 
    59.19381, 59.18636, 59.17861, 59.17054, 59.16215, 59.15346, 59.14445, 
    59.13513, 59.12549, 59.11555, 59.10529, 59.09472, 59.08384, 59.07265, 
    59.06116, 59.04935, 59.03723, 59.0248, 59.01206, 58.99902, 58.98566, 
    58.972, 58.95804, 58.94376, 58.92918, 58.9143, 58.89911, 58.88361, 
    58.86781, 58.8517, 58.8353, 58.81858, 58.80157, 58.78426, 58.76664, 
    58.74872, 58.7305, 58.71198, 58.69316, 58.67405, 58.65463, 58.63492, 
    58.61491, 58.5946, 58.574, 58.5531, 58.53191, 58.51043, 58.48865, 
    58.46658, 58.44421, 58.42155, 58.39861, 58.37537, 58.35184, 58.32803, 
    58.30392, 58.27953, 58.25485, 58.22989, 58.20463, 58.1791, 58.15328, 
    58.12717, 58.10078, 58.07412, 58.04717, 58.01994, 57.99243, 57.96464, 
    57.93657, 57.90822, 57.8796, 57.8507, 57.82153, 57.79208, 57.76236, 
    57.73236, 57.7021, 57.67155, 57.64074, 57.60966, 57.57832, 57.5467, 
    57.51482, 57.48266, 57.45024, 57.41756, 57.38462, 57.35141, 57.31794, 
    57.2842, 57.25021, 57.21595, 57.18143, 57.14666, 57.11163, 57.07634, 
    57.0408, 57.005, 56.96895, 56.93264, 56.89608, 56.85928, 56.82222, 
    56.7849, 56.74734, 56.70954, 56.67148, 56.63318, 56.59464, 56.55584, 
    56.51681, 56.47753, 56.43801, 56.39825, 56.35825, 56.318, 56.27753, 
    56.23681, 56.19585, 56.15467, 56.11324, 56.07158, 56.02969, 55.98757, 
    55.94521, 55.90263, 55.85981, 55.81676, 55.77349, 55.73, 55.68627, 
    55.64232, 55.59815, 55.55375, 55.50913, 55.46429, 55.41922, 55.37394, 
    55.32844, 55.28272, 55.23679, 55.19064, 55.14427, 55.09769, 55.05089, 
    55.00388, 54.95666,
  49.85722, 49.92055, 49.98374, 50.04679, 50.1097, 50.17247, 50.23511, 
    50.2976, 50.35995, 50.42216, 50.48423, 50.54616, 50.60794, 50.66958, 
    50.73107, 50.79242, 50.85361, 50.91467, 50.97557, 51.03632, 51.09693, 
    51.15738, 51.21769, 51.27784, 51.33783, 51.39768, 51.45737, 51.5169, 
    51.57628, 51.63551, 51.69457, 51.75348, 51.81223, 51.87082, 51.92924, 
    51.98751, 52.04561, 52.10356, 52.16133, 52.21895, 52.2764, 52.33368, 
    52.3908, 52.44775, 52.50453, 52.56114, 52.61758, 52.67385, 52.72995, 
    52.78588, 52.84163, 52.89721, 52.95261, 53.00784, 53.06289, 53.11777, 
    53.17247, 53.22698, 53.28132, 53.33548, 53.38945, 53.44324, 53.49685, 
    53.55028, 53.60352, 53.65657, 53.70944, 53.76212, 53.81462, 53.86692, 
    53.91903, 53.97095, 54.02269, 54.07422, 54.12557, 54.17672, 54.22767, 
    54.27843, 54.32899, 54.37936, 54.42952, 54.47949, 54.52925, 54.57882, 
    54.62818, 54.67733, 54.72629, 54.77504, 54.82358, 54.87192, 54.92004, 
    54.96796, 55.01568, 55.06318, 55.11047, 55.15754, 55.20441, 55.25106, 
    55.2975, 55.34372, 55.38972, 55.43551, 55.48108, 55.52642, 55.57156, 
    55.61646, 55.66115, 55.70561, 55.74985, 55.79387, 55.83765, 55.88122, 
    55.92455, 55.96766, 56.01054, 56.05319, 56.09561, 56.13779, 56.17974, 
    56.22147, 56.26295, 56.3042, 56.34521, 56.38599, 56.42653, 56.46683, 
    56.50689, 56.54671, 56.58628, 56.62562, 56.66471, 56.70356, 56.74216, 
    56.78052, 56.81863, 56.85649, 56.8941, 56.93147, 56.96858, 57.00544, 
    57.04205, 57.0784, 57.11451, 57.15036, 57.18595, 57.22128, 57.25636, 
    57.29118, 57.32574, 57.36005, 57.39408, 57.42786, 57.46138, 57.49464, 
    57.52763, 57.56035, 57.59281, 57.625, 57.65693, 57.68858, 57.71997, 
    57.75109, 57.78194, 57.81252, 57.84282, 57.87285, 57.90261, 57.93209, 
    57.9613, 57.99023, 58.01889, 58.04726, 58.07536, 58.10318, 58.13073, 
    58.15799, 58.18496, 58.21166, 58.23807, 58.2642, 58.29005, 58.31561, 
    58.34089, 58.36587, 58.39058, 58.41499, 58.43911, 58.46295, 58.4865, 
    58.50975, 58.53271, 58.55539, 58.57777, 58.59986, 58.62165, 58.64315, 
    58.66436, 58.68526, 58.70588, 58.72619, 58.74621, 58.76593, 58.78535, 
    58.80448, 58.8233, 58.84183, 58.86005, 58.87797, 58.89559, 58.91291, 
    58.92992, 58.94663, 58.96304, 58.97914, 58.99494, 59.01043, 59.02562, 
    59.0405, 59.05507, 59.06934, 59.0833, 59.09695, 59.11029, 59.12333, 
    59.13605, 59.14847, 59.16057, 59.17237, 59.18385, 59.19502, 59.20588, 
    59.21643, 59.22667, 59.2366, 59.24621, 59.2555, 59.26449, 59.27316, 
    59.28152, 59.28957, 59.29729, 59.30471, 59.31181, 59.3186, 59.32507, 
    59.33122, 59.33706, 59.34258, 59.34779, 59.35268, 59.35725, 59.36151, 
    59.36545, 59.36907, 59.37238, 59.37537, 59.37804, 59.3804, 59.38243, 
    59.38416, 59.38556, 59.38665, 59.38741, 59.38787, 59.388, 59.38781, 
    59.38731, 59.38649, 59.38536, 59.3839, 59.38213, 59.38005, 59.37764, 
    59.37492, 59.37188, 59.36852, 59.36485, 59.36086, 59.35655, 59.35192, 
    59.34698, 59.34173, 59.33615, 59.33027, 59.32406, 59.31754, 59.31071, 
    59.30356, 59.29609, 59.28831, 59.28022, 59.27181, 59.26309, 59.25406, 
    59.24471, 59.23505, 59.22507, 59.21479, 59.20419, 59.19328, 59.18205, 
    59.17052, 59.15868, 59.14652, 59.13406, 59.12128, 59.1082, 59.09481, 
    59.08111, 59.0671, 59.05279, 59.03817, 59.02324, 59.008, 58.99246, 
    58.97662, 58.96046, 58.94401, 58.92725, 58.91019, 58.89282, 58.87516, 
    58.85719, 58.83892, 58.82035, 58.80148, 58.7823, 58.76283, 58.74306, 
    58.723, 58.70264, 58.68198, 58.66102, 58.63977, 58.61823, 58.59638, 
    58.57425, 58.55182, 58.5291, 58.50609, 58.48279, 58.4592, 58.43531, 
    58.41114, 58.38668, 58.36194, 58.33691, 58.31158, 58.28598, 58.26009, 
    58.23391, 58.20745, 58.18071, 58.15369, 58.12639, 58.0988, 58.07094, 
    58.0428, 58.01437, 57.98568, 57.9567, 57.92745, 57.89792, 57.86812, 
    57.83804, 57.8077, 57.77708, 57.74619, 57.71503, 57.68359, 57.65189, 
    57.61993, 57.58769, 57.55519, 57.52242, 57.48939, 57.4561, 57.42254, 
    57.38872, 57.35464, 57.32029, 57.28569, 57.25083, 57.21571, 57.18033, 
    57.1447, 57.10881, 57.07267, 57.03627, 56.99962, 56.96272, 56.92557, 
    56.88817, 56.85051, 56.81261, 56.77447, 56.73607, 56.69743, 56.65854, 
    56.61942, 56.58004, 56.54042, 56.50057, 56.46047, 56.42013, 56.37956, 
    56.33874, 56.29769, 56.2564, 56.21488, 56.17313, 56.13113, 56.08891, 
    56.04646, 56.00377, 55.96086, 55.91771, 55.87434, 55.83075, 55.78692, 
    55.74287, 55.69859, 55.65409, 55.60938, 55.56443, 55.51927, 55.47388, 
    55.42828, 55.38246, 55.33642, 55.29016, 55.24369, 55.19701, 55.15011, 
    55.103, 55.05568,
  49.94656, 50.00998, 50.07327, 50.13642, 50.19943, 50.26231, 50.32504, 
    50.38763, 50.45009, 50.5124, 50.57457, 50.6366, 50.69848, 50.76022, 
    50.82181, 50.88326, 50.94456, 51.00571, 51.06671, 51.12757, 51.18827, 
    51.24883, 51.30923, 51.36949, 51.42959, 51.48954, 51.54933, 51.60897, 
    51.66845, 51.72778, 51.78695, 51.84595, 51.90481, 51.9635, 52.02203, 
    52.0804, 52.13861, 52.19666, 52.25454, 52.31226, 52.36981, 52.4272, 
    52.48442, 52.54147, 52.59836, 52.65508, 52.71162, 52.768, 52.8242, 
    52.88023, 52.93609, 52.99178, 53.04728, 53.10262, 53.15778, 53.21275, 
    53.26756, 53.32218, 53.37662, 53.43089, 53.48497, 53.53886, 53.59258, 
    53.64611, 53.69946, 53.75262, 53.80559, 53.85838, 53.91097, 53.96338, 
    54.0156, 54.06763, 54.11946, 54.17111, 54.22256, 54.27381, 54.32487, 
    54.37574, 54.4264, 54.47687, 54.52714, 54.57721, 54.62708, 54.67675, 
    54.72622, 54.77548, 54.82454, 54.87339, 54.92204, 54.97048, 55.01871, 
    55.06673, 55.11455, 55.16215, 55.20955, 55.25673, 55.3037, 55.35045, 
    55.39699, 55.44331, 55.48942, 55.53531, 55.58098, 55.62643, 55.67166, 
    55.71667, 55.76146, 55.80602, 55.85036, 55.89448, 55.93837, 55.98203, 
    56.02547, 56.06868, 56.11166, 56.1544, 56.19692, 56.2392, 56.28126, 
    56.32307, 56.36466, 56.40601, 56.44712, 56.48799, 56.52863, 56.56902, 
    56.60918, 56.6491, 56.68877, 56.7282, 56.76739, 56.80633, 56.84502, 
    56.88348, 56.92168, 56.95963, 56.99734, 57.03479, 57.072, 57.10896, 
    57.14566, 57.1821, 57.2183, 57.25423, 57.28992, 57.32534, 57.36051, 
    57.39542, 57.43007, 57.46446, 57.49858, 57.53245, 57.56606, 57.5994, 
    57.63247, 57.66528, 57.69782, 57.7301, 57.76211, 57.79385, 57.82532, 
    57.85652, 57.88745, 57.91811, 57.94849, 57.9786, 58.00844, 58.038, 
    58.06729, 58.09629, 58.12503, 58.15348, 58.18166, 58.20955, 58.23717, 
    58.2645, 58.29155, 58.31832, 58.3448, 58.37101, 58.39692, 58.42255, 
    58.4479, 58.47295, 58.49772, 58.52221, 58.5464, 58.5703, 58.59391, 
    58.61723, 58.64026, 58.66299, 58.68544, 58.70759, 58.72944, 58.751, 
    58.77227, 58.79324, 58.81391, 58.83428, 58.85435, 58.87413, 58.89361, 
    58.91279, 58.93166, 58.95024, 58.96851, 58.98649, 59.00416, 59.02152, 
    59.03859, 59.05535, 59.0718, 59.08795, 59.10379, 59.11933, 59.13456, 
    59.14948, 59.1641, 59.17841, 59.19241, 59.2061, 59.21948, 59.23255, 
    59.24531, 59.25776, 59.2699, 59.28173, 59.29325, 59.30445, 59.31535, 
    59.32593, 59.33619, 59.34615, 59.35579, 59.36512, 59.37413, 59.38282, 
    59.39121, 59.39928, 59.40703, 59.41446, 59.42159, 59.42839, 59.43488, 
    59.44105, 59.44691, 59.45245, 59.45767, 59.46257, 59.46716, 59.47143, 
    59.47538, 59.47902, 59.48233, 59.48533, 59.48801, 59.49038, 59.49242, 
    59.49414, 59.49555, 59.49664, 59.49741, 59.49786, 59.498, 59.49781, 
    59.49731, 59.49649, 59.49535, 59.49389, 59.49212, 59.49002, 59.48761, 
    59.48488, 59.48183, 59.47846, 59.47478, 59.47078, 59.46645, 59.46182, 
    59.45686, 59.45159, 59.446, 59.44009, 59.43387, 59.42733, 59.42048, 
    59.41331, 59.40582, 59.39802, 59.3899, 59.38147, 59.37272, 59.36366, 
    59.35429, 59.34459, 59.33459, 59.32428, 59.31364, 59.3027, 59.29145, 
    59.27988, 59.26801, 59.25581, 59.24331, 59.2305, 59.21738, 59.20395, 
    59.19021, 59.17617, 59.16181, 59.14714, 59.13217, 59.11689, 59.10131, 
    59.08541, 59.06922, 59.05272, 59.03591, 59.0188, 59.00138, 58.98367, 
    58.96564, 58.94732, 58.9287, 58.90977, 58.89055, 58.87103, 58.8512, 
    58.83108, 58.81066, 58.78994, 58.76892, 58.74761, 58.72601, 58.70411, 
    58.68191, 58.65942, 58.63664, 58.61356, 58.59019, 58.56654, 58.54259, 
    58.51835, 58.49382, 58.46901, 58.44391, 58.41852, 58.39284, 58.36688, 
    58.34063, 58.3141, 58.28729, 58.26019, 58.23281, 58.20516, 58.17722, 
    58.149, 58.1205, 58.09172, 58.06267, 58.03334, 58.00374, 57.97386, 
    57.9437, 57.91327, 57.88258, 57.8516, 57.82036, 57.78885, 57.75706, 
    57.72501, 57.69269, 57.66011, 57.62725, 57.59414, 57.56076, 57.52711, 
    57.49321, 57.45903, 57.4246, 57.38991, 57.35497, 57.31976, 57.28429, 
    57.24857, 57.21259, 57.17635, 57.13987, 57.10313, 57.06613, 57.02889, 
    56.99139, 56.95365, 56.91565, 56.87741, 56.83892, 56.80019, 56.7612, 
    56.72198, 56.68251, 56.6428, 56.60284, 56.56265, 56.52222, 56.48154, 
    56.44063, 56.39948, 56.3581, 56.31647, 56.27462, 56.23253, 56.19021, 
    56.14766, 56.10487, 56.06186, 56.01861, 55.97514, 55.93144, 55.88752, 
    55.84336, 55.79899, 55.75439, 55.70956, 55.66452, 55.61926, 55.57377, 
    55.52806, 55.48214, 55.436, 55.38964, 55.34307, 55.29628, 55.24928, 
    55.20206, 55.15464,
  50.03581, 50.09933, 50.16272, 50.22597, 50.28908, 50.35205, 50.41489, 
    50.47758, 50.54013, 50.60255, 50.66482, 50.72694, 50.78893, 50.85077, 
    50.91246, 50.97401, 51.03541, 51.09667, 51.15778, 51.21873, 51.27954, 
    51.3402, 51.40071, 51.46106, 51.52127, 51.58131, 51.64121, 51.70095, 
    51.76054, 51.81997, 51.87924, 51.93835, 51.99731, 52.05611, 52.11474, 
    52.17322, 52.23153, 52.28968, 52.34767, 52.40549, 52.46315, 52.52064, 
    52.57796, 52.63512, 52.69212, 52.74894, 52.80559, 52.86207, 52.91838, 
    52.97451, 53.03048, 53.08627, 53.14188, 53.19732, 53.25258, 53.30767, 
    53.36258, 53.4173, 53.47186, 53.52622, 53.58041, 53.63441, 53.68823, 
    53.74187, 53.79532, 53.84859, 53.90167, 53.95456, 54.00726, 54.05978, 
    54.1121, 54.16423, 54.21618, 54.26793, 54.31948, 54.37084, 54.422, 
    54.47298, 54.52375, 54.57432, 54.6247, 54.67487, 54.72485, 54.77462, 
    54.82419, 54.87356, 54.92272, 54.97168, 55.02043, 55.06898, 55.11731, 
    55.16544, 55.21336, 55.26107, 55.30857, 55.35585, 55.40292, 55.44978, 
    55.49643, 55.54285, 55.58906, 55.63505, 55.68083, 55.72638, 55.77171, 
    55.81683, 55.86171, 55.90638, 55.95082, 55.99504, 56.03903, 56.0828, 
    56.12634, 56.16964, 56.21272, 56.25557, 56.29819, 56.34057, 56.38272, 
    56.42464, 56.46632, 56.50777, 56.54898, 56.58995, 56.63068, 56.67118, 
    56.71143, 56.75144, 56.79121, 56.83074, 56.87002, 56.90906, 56.94785, 
    56.98639, 57.02469, 57.06274, 57.10054, 57.13809, 57.17538, 57.21243, 
    57.24923, 57.28576, 57.32205, 57.35808, 57.39385, 57.42937, 57.46462, 
    57.49962, 57.53436, 57.56884, 57.60305, 57.637, 57.6707, 57.70412, 
    57.73728, 57.77018, 57.80281, 57.83517, 57.86726, 57.89908, 57.93064, 
    57.96192, 57.99293, 58.02367, 58.05413, 58.08432, 58.11424, 58.14388, 
    58.17325, 58.20234, 58.23114, 58.25967, 58.28793, 58.3159, 58.34359, 
    58.37099, 58.39812, 58.42496, 58.45152, 58.47779, 58.50378, 58.52948, 
    58.55489, 58.58002, 58.60485, 58.62941, 58.65366, 58.67763, 58.70131, 
    58.7247, 58.74779, 58.77059, 58.79309, 58.8153, 58.83722, 58.85884, 
    58.88017, 58.90119, 58.92192, 58.94235, 58.96249, 58.98232, 59.00185, 
    59.02108, 59.04002, 59.05864, 59.07697, 59.09499, 59.11272, 59.13013, 
    59.14724, 59.16405, 59.18055, 59.19675, 59.21264, 59.22822, 59.2435, 
    59.25846, 59.27312, 59.28747, 59.30151, 59.31524, 59.32866, 59.34177, 
    59.35457, 59.36705, 59.37923, 59.39109, 59.40265, 59.41388, 59.42481, 
    59.43542, 59.44572, 59.4557, 59.46537, 59.47472, 59.48376, 59.49249, 
    59.50089, 59.50898, 59.51676, 59.52422, 59.53136, 59.53819, 59.54469, 
    59.55088, 59.55676, 59.56231, 59.56755, 59.57247, 59.57707, 59.58135, 
    59.58532, 59.58896, 59.59229, 59.59529, 59.59798, 59.60035, 59.6024, 
    59.60413, 59.60555, 59.60664, 59.60741, 59.60786, 59.608, 59.60781, 
    59.60731, 59.60649, 59.60534, 59.60388, 59.6021, 59.6, 59.59758, 
    59.59484, 59.59178, 59.58841, 59.58471, 59.58069, 59.57636, 59.57171, 
    59.56674, 59.56145, 59.55585, 59.54992, 59.54368, 59.53712, 59.53025, 
    59.52306, 59.51555, 59.50772, 59.49958, 59.49112, 59.48235, 59.47326, 
    59.46386, 59.45414, 59.44411, 59.43376, 59.4231, 59.41212, 59.40084, 
    59.38924, 59.37733, 59.3651, 59.35257, 59.33972, 59.32656, 59.31309, 
    59.29931, 59.28522, 59.27082, 59.25611, 59.2411, 59.22578, 59.21014, 
    59.19421, 59.17796, 59.16141, 59.14456, 59.1274, 59.10993, 59.09216, 
    59.07409, 59.05572, 59.03704, 59.01806, 58.99878, 58.9792, 58.95932, 
    58.93914, 58.91866, 58.89789, 58.87681, 58.85544, 58.83377, 58.81181, 
    58.78955, 58.767, 58.74416, 58.72102, 58.69758, 58.67386, 58.64985, 
    58.62554, 58.60094, 58.57606, 58.55089, 58.52543, 58.49968, 58.47365, 
    58.44733, 58.42073, 58.39384, 58.36668, 58.33922, 58.31149, 58.28347, 
    58.25518, 58.2266, 58.19775, 58.16862, 58.13921, 58.10953, 58.07957, 
    58.04933, 58.01883, 57.98804, 57.95699, 57.92566, 57.89407, 57.8622, 
    57.83007, 57.79766, 57.76499, 57.73206, 57.69885, 57.66539, 57.63165, 
    57.59766, 57.5634, 57.52888, 57.4941, 57.45906, 57.42376, 57.38821, 
    57.35239, 57.31633, 57.28, 57.24342, 57.20659, 57.1695, 57.13216, 
    57.09458, 57.05674, 57.01865, 56.98031, 56.94173, 56.9029, 56.86382, 
    56.8245, 56.78493, 56.74513, 56.70508, 56.66479, 56.62426, 56.58348, 
    56.54247, 56.50123, 56.45974, 56.41803, 56.37607, 56.33388, 56.29146, 
    56.24881, 56.20592, 56.16281, 56.11946, 56.07589, 56.03209, 55.98806, 
    55.94381, 55.89933, 55.85463, 55.8097, 55.76456, 55.71919, 55.6736, 
    55.62779, 55.58176, 55.53552, 55.48906, 55.44238, 55.39549, 55.34839, 
    55.30107, 55.25354,
  50.12497, 50.18859, 50.25208, 50.31543, 50.37864, 50.44172, 50.50465, 
    50.56744, 50.6301, 50.69261, 50.75498, 50.81721, 50.8793, 50.94124, 
    51.00303, 51.06468, 51.12619, 51.18754, 51.24875, 51.30981, 51.37072, 
    51.43148, 51.4921, 51.55256, 51.61286, 51.67301, 51.73301, 51.79286, 
    51.85255, 51.91208, 51.97145, 52.03067, 52.08973, 52.14863, 52.20737, 
    52.26595, 52.32437, 52.38263, 52.44072, 52.49865, 52.55641, 52.61401, 
    52.67144, 52.7287, 52.78579, 52.84272, 52.89948, 52.95606, 53.01248, 
    53.06872, 53.12479, 53.18069, 53.2364, 53.29195, 53.34732, 53.40251, 
    53.45752, 53.51236, 53.56701, 53.62149, 53.67578, 53.72989, 53.78382, 
    53.83756, 53.89112, 53.94449, 53.99768, 54.05067, 54.10349, 54.15611, 
    54.20853, 54.26077, 54.31282, 54.36468, 54.41634, 54.4678, 54.51908, 
    54.57015, 54.62103, 54.67171, 54.72219, 54.77247, 54.82255, 54.87243, 
    54.9221, 54.97158, 55.02085, 55.06991, 55.11877, 55.16742, 55.21586, 
    55.26409, 55.31212, 55.35993, 55.40753, 55.45492, 55.5021, 55.54906, 
    55.5958, 55.64233, 55.68865, 55.73474, 55.78062, 55.82627, 55.87171, 
    55.91693, 55.96192, 56.00669, 56.05123, 56.09555, 56.13964, 56.18351, 
    56.22715, 56.27056, 56.31374, 56.35669, 56.3994, 56.44189, 56.48414, 
    56.52615, 56.56794, 56.60948, 56.65079, 56.69186, 56.73269, 56.77328, 
    56.81363, 56.85374, 56.89361, 56.93323, 56.97261, 57.01174, 57.05063, 
    57.08927, 57.12766, 57.16581, 57.2037, 57.24134, 57.27873, 57.31587, 
    57.35276, 57.38939, 57.42577, 57.46189, 57.49775, 57.53336, 57.5687, 
    57.60379, 57.63862, 57.67318, 57.70749, 57.74153, 57.77531, 57.80882, 
    57.84206, 57.87505, 57.90776, 57.9402, 57.97238, 58.00429, 58.03593, 
    58.06729, 58.09838, 58.1292, 58.15975, 58.19003, 58.22002, 58.24974, 
    58.27918, 58.30835, 58.33723, 58.36584, 58.39417, 58.42222, 58.44998, 
    58.47746, 58.50466, 58.53158, 58.55821, 58.58455, 58.61061, 58.63638, 
    58.66187, 58.68707, 58.71197, 58.73659, 58.76091, 58.78495, 58.80869, 
    58.83214, 58.8553, 58.87817, 58.90073, 58.92301, 58.94498, 58.96667, 
    58.98805, 59.00914, 59.02993, 59.05042, 59.07061, 59.0905, 59.11008, 
    59.12937, 59.14835, 59.16704, 59.18542, 59.20349, 59.22126, 59.23873, 
    59.25589, 59.27275, 59.2893, 59.30554, 59.32148, 59.3371, 59.35242, 
    59.36743, 59.38213, 59.39652, 59.4106, 59.42437, 59.43784, 59.45098, 
    59.46382, 59.47634, 59.48855, 59.50045, 59.51204, 59.52331, 59.53426, 
    59.54491, 59.55524, 59.56525, 59.57494, 59.58433, 59.59339, 59.60214, 
    59.61057, 59.61869, 59.62649, 59.63397, 59.64113, 59.64798, 59.6545, 
    59.66071, 59.6666, 59.67217, 59.67743, 59.68236, 59.68697, 59.69127, 
    59.69525, 59.6989, 59.70224, 59.70525, 59.70795, 59.71033, 59.71239, 
    59.71412, 59.71554, 59.71663, 59.71741, 59.71786, 59.718, 59.71782, 
    59.71731, 59.71648, 59.71534, 59.71387, 59.71208, 59.70997, 59.70755, 
    59.7048, 59.70173, 59.69835, 59.69464, 59.69061, 59.68627, 59.6816, 
    59.67662, 59.67131, 59.66569, 59.65975, 59.65349, 59.64692, 59.64002, 
    59.6328, 59.62527, 59.61742, 59.60926, 59.60078, 59.59198, 59.58286, 
    59.57343, 59.56369, 59.55362, 59.54324, 59.53255, 59.52155, 59.51022, 
    59.49859, 59.48664, 59.47438, 59.46181, 59.44893, 59.43573, 59.42222, 
    59.4084, 59.39427, 59.37983, 59.36508, 59.35002, 59.33465, 59.31897, 
    59.30299, 59.2867, 59.2701, 59.2532, 59.23599, 59.21847, 59.20065, 
    59.18253, 59.1641, 59.14537, 59.12634, 59.10701, 59.08737, 59.06743, 
    59.0472, 59.02666, 59.00582, 58.98469, 58.96326, 58.94153, 58.91951, 
    58.89718, 58.87457, 58.85166, 58.82845, 58.80495, 58.78117, 58.75708, 
    58.73271, 58.70805, 58.6831, 58.65786, 58.63233, 58.60651, 58.58041, 
    58.55402, 58.52734, 58.50038, 58.47314, 58.44561, 58.4178, 58.38971, 
    58.36134, 58.33268, 58.30375, 58.27454, 58.24506, 58.21529, 58.18525, 
    58.15494, 58.12435, 58.09349, 58.06235, 58.03094, 57.99926, 57.96731, 
    57.93509, 57.9026, 57.86985, 57.83682, 57.80354, 57.76998, 57.73616, 
    57.70208, 57.66773, 57.63313, 57.59826, 57.56313, 57.52774, 57.49209, 
    57.45619, 57.42003, 57.38361, 57.34694, 57.31001, 57.27283, 57.2354, 
    57.19772, 57.15979, 57.1216, 57.08318, 57.04449, 57.00557, 56.9664, 
    56.92698, 56.88732, 56.84741, 56.80727, 56.76688, 56.72625, 56.68538, 
    56.64427, 56.60292, 56.56134, 56.51952, 56.47747, 56.43518, 56.39266, 
    56.34991, 56.30692, 56.26371, 56.22026, 56.17659, 56.13269, 56.08855, 
    56.0442, 55.99962, 55.95482, 55.90979, 55.86454, 55.81907, 55.77338, 
    55.72747, 55.68134, 55.63499, 55.58842, 55.54165, 55.49465, 55.44744, 
    55.40002, 55.35238,
  50.21405, 50.27777, 50.34136, 50.40481, 50.46812, 50.53129, 50.59433, 
    50.65722, 50.71998, 50.78259, 50.84506, 50.90739, 50.96958, 51.03162, 
    51.09352, 51.15527, 51.21688, 51.27834, 51.33965, 51.40081, 51.46182, 
    51.52269, 51.5834, 51.64396, 51.70437, 51.76463, 51.82473, 51.88468, 
    51.94447, 52.00411, 52.06359, 52.12291, 52.18208, 52.24108, 52.29993, 
    52.35861, 52.41713, 52.47549, 52.53369, 52.59172, 52.64959, 52.70729, 
    52.76483, 52.8222, 52.8794, 52.93643, 52.99329, 53.04998, 53.10651, 
    53.16285, 53.21903, 53.27503, 53.33086, 53.38651, 53.44198, 53.49728, 
    53.5524, 53.60734, 53.6621, 53.71668, 53.77108, 53.8253, 53.87933, 
    53.93318, 53.98684, 54.04033, 54.09362, 54.14672, 54.19963, 54.25237, 
    54.3049, 54.35725, 54.4094, 54.46136, 54.51313, 54.5647, 54.61608, 
    54.66726, 54.71825, 54.76903, 54.81962, 54.87, 54.92019, 54.97018, 
    55.01996, 55.06953, 55.11891, 55.16808, 55.21704, 55.2658, 55.31435, 
    55.36268, 55.41081, 55.45873, 55.50644, 55.55393, 55.60121, 55.64828, 
    55.69513, 55.74176, 55.78818, 55.83438, 55.88036, 55.92612, 55.97166, 
    56.01698, 56.06207, 56.10694, 56.15159, 56.19601, 56.2402, 56.28417, 
    56.32791, 56.37142, 56.4147, 56.45775, 56.50057, 56.54316, 56.58551, 
    56.62762, 56.66951, 56.71115, 56.75256, 56.79372, 56.83466, 56.87534, 
    56.91579, 56.956, 56.99596, 57.03568, 57.07516, 57.11439, 57.15337, 
    57.19211, 57.23059, 57.26883, 57.30682, 57.34456, 57.38204, 57.41927, 
    57.45625, 57.49298, 57.52945, 57.56566, 57.60161, 57.63731, 57.67274, 
    57.70792, 57.74284, 57.7775, 57.81189, 57.84602, 57.87988, 57.91348, 
    57.94682, 57.97989, 58.01268, 58.04522, 58.07748, 58.10947, 58.14119, 
    58.17264, 58.20381, 58.23471, 58.26534, 58.2957, 58.32577, 58.35557, 
    58.38509, 58.41434, 58.4433, 58.47199, 58.50039, 58.52851, 58.55635, 
    58.58391, 58.61119, 58.63818, 58.66488, 58.6913, 58.71743, 58.74327, 
    58.76883, 58.79409, 58.81907, 58.84375, 58.86814, 58.89225, 58.91606, 
    58.93958, 58.9628, 58.98573, 59.00836, 59.0307, 59.05273, 59.07448, 
    59.09592, 59.11707, 59.13792, 59.15847, 59.17871, 59.19866, 59.2183, 
    59.23764, 59.25668, 59.27542, 59.29385, 59.31198, 59.3298, 59.34732, 
    59.36453, 59.38144, 59.39803, 59.41432, 59.43031, 59.44598, 59.46134, 
    59.47639, 59.49114, 59.50557, 59.5197, 59.5335, 59.547, 59.56019, 
    59.57306, 59.58562, 59.59787, 59.60981, 59.62143, 59.63273, 59.64372, 
    59.65439, 59.66475, 59.67479, 59.68452, 59.69393, 59.70302, 59.7118, 
    59.72025, 59.72839, 59.73621, 59.74372, 59.7509, 59.75777, 59.76431, 
    59.77054, 59.77645, 59.78204, 59.7873, 59.79226, 59.79688, 59.80119, 
    59.80518, 59.80885, 59.81219, 59.81522, 59.81792, 59.8203, 59.82237, 
    59.82411, 59.82553, 59.82663, 59.82741, 59.82787, 59.828, 59.82781, 
    59.8273, 59.82648, 59.82533, 59.82386, 59.82206, 59.81995, 59.81752, 
    59.81476, 59.81168, 59.80828, 59.80457, 59.80053, 59.79617, 59.79149, 
    59.7865, 59.78117, 59.77554, 59.76958, 59.7633, 59.7567, 59.74979, 
    59.74255, 59.735, 59.72713, 59.71894, 59.71043, 59.7016, 59.69246, 
    59.683, 59.67323, 59.66313, 59.65273, 59.642, 59.63096, 59.61961, 
    59.60794, 59.59595, 59.58366, 59.57105, 59.55812, 59.54489, 59.53134, 
    59.51748, 59.50331, 59.48883, 59.47403, 59.45893, 59.44352, 59.4278, 
    59.41177, 59.39543, 59.37878, 59.36183, 59.34457, 59.327, 59.30914, 
    59.29096, 59.27248, 59.25369, 59.2346, 59.21521, 59.19552, 59.17553, 
    59.15524, 59.13464, 59.11375, 59.09255, 59.07106, 59.04927, 59.02718, 
    59.0048, 58.98212, 58.95914, 58.93587, 58.91231, 58.88845, 58.86431, 
    58.83987, 58.81514, 58.79012, 58.7648, 58.7392, 58.71331, 58.68714, 
    58.66068, 58.63393, 58.60689, 58.57957, 58.55197, 58.52409, 58.49592, 
    58.46747, 58.43874, 58.40973, 58.38044, 58.35088, 58.32103, 58.29091, 
    58.26052, 58.22984, 58.1989, 58.16768, 58.13619, 58.10442, 58.07239, 
    58.04008, 58.00751, 57.97467, 57.94156, 57.90818, 57.87454, 57.84064, 
    57.80647, 57.77203, 57.73734, 57.70238, 57.66716, 57.63168, 57.59594, 
    57.55995, 57.52369, 57.48719, 57.45042, 57.4134, 57.37613, 57.3386, 
    57.30083, 57.2628, 57.22452, 57.186, 57.14722, 57.1082, 57.06893, 
    57.02942, 56.98966, 56.94966, 56.90941, 56.86892, 56.8282, 56.78723, 
    56.74602, 56.70458, 56.6629, 56.62098, 56.57882, 56.53643, 56.49381, 
    56.45096, 56.40787, 56.36456, 56.32101, 56.27723, 56.23323, 56.189, 
    56.14454, 56.09986, 56.05495, 56.00982, 55.96447, 55.9189, 55.8731, 
    55.82708, 55.78085, 55.7344, 55.68773, 55.64085, 55.59375, 55.54643, 
    55.49891, 55.45116,
  50.30304, 50.36686, 50.43055, 50.49409, 50.55751, 50.62078, 50.68392, 
    50.74691, 50.80977, 50.87249, 50.93506, 50.99749, 51.05978, 51.12192, 
    51.18392, 51.24577, 51.30748, 51.36905, 51.43046, 51.49172, 51.55284, 
    51.61381, 51.67463, 51.73529, 51.7958, 51.85616, 51.91637, 51.97642, 
    52.03632, 52.09606, 52.15564, 52.21507, 52.27434, 52.33345, 52.3924, 
    52.45119, 52.50982, 52.56828, 52.62658, 52.68472, 52.74269, 52.8005, 
    52.85814, 52.91562, 52.97292, 53.03006, 53.08703, 53.14383, 53.20045, 
    53.25691, 53.31319, 53.3693, 53.42523, 53.48099, 53.53657, 53.59198, 
    53.6472, 53.70225, 53.75712, 53.8118, 53.86631, 53.92063, 53.97477, 
    54.02873, 54.0825, 54.13609, 54.18948, 54.24269, 54.29572, 54.34855, 
    54.4012, 54.45365, 54.50591, 54.55798, 54.60985, 54.66153, 54.71302, 
    54.76431, 54.8154, 54.86629, 54.91698, 54.96748, 55.01777, 55.06786, 
    55.11774, 55.16743, 55.21691, 55.26619, 55.31525, 55.36412, 55.41277, 
    55.46121, 55.50945, 55.55747, 55.60528, 55.65288, 55.70027, 55.74744, 
    55.79439, 55.84113, 55.88765, 55.93396, 55.98004, 56.02591, 56.07155, 
    56.11697, 56.16217, 56.20714, 56.25189, 56.29642, 56.34071, 56.38478, 
    56.42863, 56.47224, 56.51562, 56.55877, 56.60169, 56.64437, 56.68683, 
    56.72905, 56.77103, 56.81277, 56.85428, 56.89555, 56.93657, 56.97736, 
    57.01791, 57.05821, 57.09827, 57.13809, 57.17767, 57.21699, 57.25607, 
    57.2949, 57.33348, 57.37182, 57.4099, 57.44773, 57.48531, 57.52264, 
    57.55971, 57.59653, 57.63309, 57.66939, 57.70544, 57.74123, 57.77676, 
    57.81202, 57.84703, 57.88177, 57.91626, 57.95047, 57.98443, 58.01812, 
    58.05154, 58.08469, 58.11758, 58.15019, 58.18254, 58.21461, 58.24642, 
    58.27795, 58.30921, 58.3402, 58.37091, 58.40134, 58.4315, 58.46138, 
    58.49098, 58.52031, 58.54935, 58.57811, 58.60659, 58.63479, 58.66271, 
    58.69034, 58.71769, 58.74475, 58.77153, 58.79802, 58.82422, 58.85014, 
    58.87576, 58.9011, 58.92614, 58.9509, 58.97536, 58.99953, 59.02341, 
    59.04699, 59.07028, 59.09327, 59.11597, 59.13837, 59.16047, 59.18228, 
    59.20378, 59.22499, 59.2459, 59.2665, 59.28681, 59.30681, 59.32651, 
    59.34591, 59.365, 59.38379, 59.40228, 59.42046, 59.43834, 59.4559, 
    59.47316, 59.49012, 59.50676, 59.5231, 59.53913, 59.55484, 59.57026, 
    59.58535, 59.60014, 59.61461, 59.62878, 59.64263, 59.65617, 59.6694, 
    59.6823, 59.6949, 59.70719, 59.71915, 59.73081, 59.74215, 59.75317, 
    59.76387, 59.77426, 59.78434, 59.79409, 59.80353, 59.81264, 59.82145, 
    59.82993, 59.83809, 59.84594, 59.85346, 59.86067, 59.86756, 59.87412, 
    59.88037, 59.8863, 59.8919, 59.89718, 59.90215, 59.90679, 59.91111, 
    59.91511, 59.91879, 59.92215, 59.92518, 59.92789, 59.93028, 59.93235, 
    59.9341, 59.93552, 59.93663, 59.9374, 59.93786, 59.938, 59.93781, 
    59.9373, 59.93647, 59.93532, 59.93384, 59.93204, 59.92992, 59.92748, 
    59.92472, 59.92163, 59.91823, 59.9145, 59.91045, 59.90607, 59.90138, 
    59.89637, 59.89103, 59.88538, 59.8794, 59.8731, 59.86649, 59.85955, 
    59.85229, 59.84472, 59.83682, 59.82861, 59.82008, 59.81123, 59.80206, 
    59.79257, 59.78276, 59.77264, 59.7622, 59.75145, 59.74038, 59.72898, 
    59.71728, 59.70527, 59.69293, 59.68028, 59.66732, 59.65405, 59.64046, 
    59.62656, 59.61235, 59.59782, 59.58298, 59.56784, 59.55238, 59.53661, 
    59.52053, 59.50415, 59.48745, 59.47045, 59.45314, 59.43553, 59.4176, 
    59.39938, 59.38084, 59.362, 59.34286, 59.32341, 59.30367, 59.28362, 
    59.26326, 59.24261, 59.22165, 59.2004, 59.17885, 59.15699, 59.13485, 
    59.1124, 59.08965, 59.06662, 59.04328, 59.01965, 58.99573, 58.97151, 
    58.947, 58.9222, 58.89711, 58.87173, 58.84606, 58.8201, 58.79385, 
    58.76731, 58.74049, 58.71338, 58.68599, 58.65831, 58.63035, 58.6021, 
    58.57358, 58.54477, 58.51569, 58.48632, 58.45667, 58.42675, 58.39655, 
    58.36607, 58.33531, 58.30429, 58.27298, 58.24141, 58.20956, 58.17744, 
    58.14505, 58.11239, 58.07946, 58.04627, 58.01281, 57.97908, 57.94508, 
    57.91082, 57.8763, 57.84151, 57.80646, 57.77115, 57.73558, 57.69975, 
    57.66367, 57.62732, 57.59072, 57.55386, 57.51675, 57.47939, 57.44176, 
    57.40389, 57.36577, 57.3274, 57.28878, 57.2499, 57.21078, 57.17142, 
    57.13181, 57.09195, 57.05185, 57.01151, 56.97093, 56.9301, 56.88903, 
    56.84773, 56.80618, 56.7644, 56.72238, 56.68013, 56.63764, 56.59492, 
    56.55196, 56.50877, 56.46535, 56.42171, 56.37783, 56.33372, 56.28939, 
    56.24483, 56.20004, 56.15503, 56.1098, 56.06434, 56.01867, 55.97277, 
    55.92665, 55.88031, 55.83375, 55.78698, 55.73999, 55.69278, 55.64537, 
    55.59773, 55.54989,
  50.39194, 50.45586, 50.51965, 50.5833, 50.64681, 50.71019, 50.77342, 
    50.83652, 50.89948, 50.96229, 51.02497, 51.0875, 51.14989, 51.21214, 
    51.27423, 51.33619, 51.398, 51.45967, 51.52118, 51.58255, 51.64377, 
    51.70484, 51.76576, 51.82653, 51.88715, 51.94761, 52.00792, 52.06808, 
    52.12808, 52.18793, 52.24762, 52.30715, 52.36652, 52.42574, 52.48479, 
    52.54368, 52.60242, 52.66099, 52.71939, 52.77764, 52.83572, 52.89363, 
    52.95138, 53.00896, 53.06637, 53.12362, 53.18069, 53.23759, 53.29433, 
    53.35089, 53.40728, 53.46349, 53.51953, 53.5754, 53.63108, 53.6866, 
    53.74193, 53.79708, 53.85206, 53.90685, 53.96146, 54.0159, 54.07014, 
    54.12421, 54.17809, 54.23178, 54.28528, 54.3386, 54.39173, 54.44468, 
    54.49743, 54.54998, 54.60235, 54.65453, 54.70651, 54.7583, 54.80989, 
    54.86128, 54.91248, 54.96348, 55.01428, 55.06488, 55.11528, 55.16548, 
    55.21547, 55.26526, 55.31485, 55.36423, 55.41341, 55.46237, 55.51113, 
    55.55968, 55.60802, 55.65615, 55.70407, 55.75177, 55.79926, 55.84654, 
    55.8936, 55.94044, 55.98707, 56.03348, 56.07967, 56.12564, 56.17138, 
    56.21691, 56.26221, 56.30729, 56.35214, 56.39677, 56.44117, 56.48534, 
    56.52929, 56.573, 56.61649, 56.65974, 56.70276, 56.74555, 56.7881, 
    56.83042, 56.8725, 56.91434, 56.95595, 56.99732, 57.03845, 57.07933, 
    57.11998, 57.16038, 57.20054, 57.24046, 57.28013, 57.31955, 57.35873, 
    57.39766, 57.43633, 57.47476, 57.51294, 57.55087, 57.58854, 57.62596, 
    57.66313, 57.70004, 57.73669, 57.77309, 57.80923, 57.84511, 57.88073, 
    57.91609, 57.95118, 57.98602, 58.02059, 58.0549, 58.08894, 58.12271, 
    58.15622, 58.18946, 58.22244, 58.25514, 58.28757, 58.31974, 58.35162, 
    58.38324, 58.41458, 58.44565, 58.47644, 58.50696, 58.5372, 58.56716, 
    58.59684, 58.62624, 58.65537, 58.68421, 58.71277, 58.74104, 58.76904, 
    58.79675, 58.82417, 58.85131, 58.87816, 58.90472, 58.931, 58.95699, 
    58.98268, 59.00809, 59.0332, 59.05803, 59.08256, 59.1068, 59.13074, 
    59.15439, 59.17775, 59.2008, 59.22356, 59.24603, 59.26819, 59.29006, 
    59.31163, 59.33289, 59.35386, 59.37453, 59.39489, 59.41495, 59.43471, 
    59.45416, 59.47331, 59.49216, 59.5107, 59.52893, 59.54686, 59.56447, 
    59.58178, 59.59879, 59.61548, 59.63187, 59.64794, 59.66371, 59.67916, 
    59.6943, 59.70913, 59.72365, 59.73786, 59.75175, 59.76533, 59.77859, 
    59.79154, 59.80418, 59.8165, 59.8285, 59.84019, 59.85156, 59.86261, 
    59.87335, 59.88377, 59.89388, 59.90366, 59.91312, 59.92227, 59.9311, 
    59.93961, 59.94779, 59.95566, 59.96321, 59.97044, 59.97734, 59.98393, 
    59.9902, 59.99614, 60.00176, 60.00706, 60.01204, 60.01669, 60.02103, 
    60.02504, 60.02873, 60.0321, 60.03514, 60.03786, 60.04026, 60.04234, 
    60.04409, 60.04552, 60.04662, 60.04741, 60.04786, 60.048, 60.04781, 
    60.0473, 60.04647, 60.04531, 60.04383, 60.04203, 60.0399, 60.03745, 
    60.03468, 60.03159, 60.02817, 60.02443, 60.02037, 60.01598, 60.01127, 
    60.00624, 60.00089, 59.99522, 59.98922, 59.98291, 59.97627, 59.96931, 
    59.96204, 59.95444, 59.94652, 59.93828, 59.92972, 59.92085, 59.91165, 
    59.90213, 59.8923, 59.88214, 59.87167, 59.86089, 59.84978, 59.83836, 
    59.82662, 59.81457, 59.8022, 59.78951, 59.77652, 59.7632, 59.74957, 
    59.73563, 59.72137, 59.70681, 59.69193, 59.67673, 59.66123, 59.64542, 
    59.6293, 59.61286, 59.59612, 59.57907, 59.56171, 59.54404, 59.52607, 
    59.50778, 59.4892, 59.4703, 59.4511, 59.4316, 59.4118, 59.39169, 
    59.37128, 59.35056, 59.32955, 59.30824, 59.28662, 59.26471, 59.24249, 
    59.21998, 59.19717, 59.17407, 59.15067, 59.12697, 59.10298, 59.0787, 
    59.05412, 59.02925, 59.00409, 58.97864, 58.95289, 58.92686, 58.90054, 
    58.87393, 58.84703, 58.81985, 58.79238, 58.76463, 58.73659, 58.70827, 
    58.67966, 58.65078, 58.62161, 58.59217, 58.56244, 58.53243, 58.50215, 
    58.47159, 58.44075, 58.40965, 58.37826, 58.3466, 58.31467, 58.28246, 
    58.24998, 58.21724, 58.18423, 58.15094, 58.11739, 58.08357, 58.04949, 
    58.01514, 57.98053, 57.94565, 57.91051, 57.87511, 57.83945, 57.80353, 
    57.76735, 57.73091, 57.69422, 57.65726, 57.62006, 57.5826, 57.54489, 
    57.50692, 57.4687, 57.43023, 57.39151, 57.35255, 57.31333, 57.27387, 
    57.23416, 57.19421, 57.15401, 57.11357, 57.07288, 57.03196, 56.99079, 
    56.94939, 56.90774, 56.86586, 56.82374, 56.78138, 56.73879, 56.69597, 
    56.65291, 56.60962, 56.5661, 56.52235, 56.47837, 56.43416, 56.38972, 
    56.34506, 56.30017, 56.25506, 56.20972, 56.16416, 56.11838, 56.07238, 
    56.02615, 55.97971, 55.93305, 55.88617, 55.83908, 55.79177, 55.74424, 
    55.6965, 55.64855,
  50.48075, 50.54478, 50.60866, 50.67241, 50.73602, 50.7995, 50.86284, 
    50.92604, 50.98909, 51.05201, 51.11479, 51.17742, 51.23991, 51.30226, 
    51.36447, 51.42653, 51.48844, 51.55021, 51.61182, 51.6733, 51.73462, 
    51.7958, 51.85682, 51.91769, 51.97841, 52.03898, 52.0994, 52.15966, 
    52.21976, 52.27971, 52.3395, 52.39914, 52.45862, 52.51794, 52.5771, 
    52.6361, 52.69494, 52.75362, 52.81213, 52.87048, 52.92867, 52.98668, 
    53.04454, 53.10222, 53.15974, 53.21709, 53.27428, 53.33129, 53.38813, 
    53.44479, 53.50129, 53.55761, 53.61376, 53.66973, 53.72552, 53.78114, 
    53.83658, 53.89185, 53.94693, 54.00183, 54.05655, 54.11108, 54.16544, 
    54.21961, 54.2736, 54.3274, 54.38101, 54.43444, 54.48767, 54.54073, 
    54.59358, 54.64625, 54.69873, 54.75101, 54.8031, 54.85499, 54.90669, 
    54.95819, 55.0095, 55.0606, 55.11151, 55.16222, 55.21273, 55.26303, 
    55.31313, 55.36303, 55.41272, 55.46221, 55.51149, 55.56057, 55.60943, 
    55.65809, 55.70654, 55.75477, 55.8028, 55.85061, 55.8982, 55.94558, 
    55.99275, 56.0397, 56.08643, 56.13294, 56.17924, 56.22531, 56.27116, 
    56.31679, 56.3622, 56.40738, 56.45234, 56.49707, 56.54157, 56.58585, 
    56.62989, 56.67371, 56.7173, 56.76065, 56.80378, 56.84667, 56.88932, 
    56.93174, 56.97392, 57.01587, 57.05758, 57.09904, 57.14027, 57.18126, 
    57.222, 57.26251, 57.30276, 57.34278, 57.38255, 57.42207, 57.46134, 
    57.50037, 57.53914, 57.57767, 57.61594, 57.65396, 57.69173, 57.72925, 
    57.76651, 57.80351, 57.84026, 57.87675, 57.91298, 57.94896, 57.98466, 
    58.02011, 58.05531, 58.09023, 58.12489, 58.15929, 58.19342, 58.22728, 
    58.26088, 58.29421, 58.32727, 58.36006, 58.39258, 58.42482, 58.4568, 
    58.4885, 58.51992, 58.55108, 58.58195, 58.61255, 58.64287, 58.67291, 
    58.70268, 58.73216, 58.76136, 58.79028, 58.81892, 58.84727, 58.87534, 
    58.90313, 58.93063, 58.95784, 58.98477, 59.01141, 59.03775, 59.06381, 
    59.08958, 59.11506, 59.14025, 59.16514, 59.18974, 59.21405, 59.23806, 
    59.26177, 59.28519, 59.30832, 59.33114, 59.35367, 59.3759, 59.39783, 
    59.41946, 59.44078, 59.46181, 59.48254, 59.50296, 59.52308, 59.54289, 
    59.5624, 59.58161, 59.60051, 59.6191, 59.63739, 59.65536, 59.67303, 
    59.6904, 59.70745, 59.72419, 59.74063, 59.75675, 59.77256, 59.78806, 
    59.80325, 59.81812, 59.83268, 59.84693, 59.86086, 59.87448, 59.88778, 
    59.90077, 59.91344, 59.9258, 59.93784, 59.94957, 59.96097, 59.97206, 
    59.98283, 59.99328, 60.00341, 60.01322, 60.02272, 60.03189, 60.04074, 
    60.04928, 60.05749, 60.06538, 60.07295, 60.0802, 60.08713, 60.09373, 
    60.10002, 60.10598, 60.11162, 60.11694, 60.12193, 60.1266, 60.13095, 
    60.13497, 60.13867, 60.14205, 60.1451, 60.14783, 60.15023, 60.15232, 
    60.15408, 60.15551, 60.15662, 60.1574, 60.15786, 60.158, 60.15781, 
    60.1573, 60.15646, 60.1553, 60.15382, 60.15201, 60.14988, 60.14742, 
    60.14464, 60.14154, 60.13811, 60.13436, 60.13028, 60.12588, 60.12116, 
    60.11612, 60.11075, 60.10506, 60.09905, 60.09271, 60.08606, 60.07908, 
    60.07178, 60.06416, 60.05621, 60.04795, 60.03936, 60.03046, 60.02124, 
    60.01169, 60.00183, 59.99165, 59.98114, 59.97033, 59.95919, 59.94773, 
    59.93596, 59.92387, 59.91146, 59.89874, 59.8857, 59.87235, 59.85868, 
    59.8447, 59.8304, 59.81579, 59.80087, 59.78563, 59.77008, 59.75422, 
    59.73805, 59.72157, 59.70477, 59.68767, 59.67026, 59.65254, 59.63451, 
    59.61618, 59.59754, 59.57859, 59.55934, 59.53978, 59.51992, 59.49975, 
    59.47928, 59.45851, 59.43743, 59.41606, 59.39438, 59.3724, 59.35013, 
    59.32755, 59.30468, 59.28151, 59.25804, 59.23428, 59.21022, 59.18587, 
    59.16122, 59.13628, 59.11105, 59.08553, 59.05971, 59.0336, 59.00721, 
    58.98053, 58.95356, 58.9263, 58.89875, 58.87092, 58.84281, 58.81441, 
    58.78572, 58.75676, 58.72752, 58.69799, 58.66818, 58.6381, 58.60773, 
    58.57709, 58.54617, 58.51497, 58.4835, 58.45176, 58.41974, 58.38745, 
    58.35489, 58.32206, 58.28896, 58.25558, 58.22195, 58.18804, 58.15387, 
    58.11943, 58.08472, 58.04976, 58.01453, 57.97903, 57.94328, 57.90727, 
    57.87099, 57.83447, 57.79768, 57.76063, 57.72333, 57.68578, 57.64796, 
    57.60991, 57.57159, 57.53302, 57.49421, 57.45515, 57.41583, 57.37627, 
    57.33646, 57.29641, 57.25611, 57.21558, 57.17479, 57.13377, 57.0925, 
    57.05099, 57.00925, 56.96727, 56.92505, 56.88259, 56.8399, 56.79697, 
    56.75381, 56.71042, 56.6668, 56.62294, 56.57886, 56.53455, 56.49001, 
    56.44524, 56.40025, 56.35503, 56.30959, 56.26392, 56.21804, 56.17193, 
    56.1256, 56.07905, 56.03229, 55.9853, 55.9381, 55.89069, 55.84306, 
    55.79521, 55.74715,
  50.56948, 50.6336, 50.69759, 50.76144, 50.82515, 50.88873, 50.95216, 
    51.01546, 51.07862, 51.14164, 51.20452, 51.26726, 51.32985, 51.3923, 
    51.45461, 51.51677, 51.57879, 51.64066, 51.70238, 51.76396, 51.82538, 
    51.88666, 51.94779, 52.00877, 52.06959, 52.13026, 52.19078, 52.25115, 
    52.31136, 52.37141, 52.43131, 52.49105, 52.55064, 52.61006, 52.66933, 
    52.72844, 52.78738, 52.84616, 52.90478, 52.96324, 53.02153, 53.07965, 
    53.13762, 53.19541, 53.25304, 53.31049, 53.36778, 53.4249, 53.48185, 
    53.53862, 53.59522, 53.65165, 53.7079, 53.76398, 53.81989, 53.87561, 
    53.93116, 53.98653, 54.04172, 54.09673, 54.15156, 54.2062, 54.26067, 
    54.31495, 54.36904, 54.42295, 54.47667, 54.5302, 54.58355, 54.6367, 
    54.68967, 54.74245, 54.79503, 54.84742, 54.89962, 54.95162, 55.00343, 
    55.05503, 55.10645, 55.15766, 55.20868, 55.25949, 55.31011, 55.36052, 
    55.41073, 55.46074, 55.51054, 55.56013, 55.60952, 55.6587, 55.70767, 
    55.75644, 55.80499, 55.85333, 55.90146, 55.94938, 55.99708, 56.04457, 
    56.09184, 56.1389, 56.18573, 56.23235, 56.27875, 56.32493, 56.37088, 
    56.41662, 56.46213, 56.50742, 56.55248, 56.59731, 56.64192, 56.6863, 
    56.73045, 56.77437, 56.81806, 56.86152, 56.90475, 56.94774, 56.99049, 
    57.03302, 57.0753, 57.11735, 57.15915, 57.20072, 57.24205, 57.28314, 
    57.32398, 57.36459, 57.40494, 57.44505, 57.48492, 57.52454, 57.56391, 
    57.60303, 57.64191, 57.68053, 57.7189, 57.75702, 57.79488, 57.83249, 
    57.86985, 57.90695, 57.94379, 57.98037, 58.0167, 58.05276, 58.08857, 
    58.12411, 58.15939, 58.1944, 58.22916, 58.26365, 58.29787, 58.33182, 
    58.36551, 58.39892, 58.43207, 58.46495, 58.49755, 58.52988, 58.56194, 
    58.59373, 58.62524, 58.65648, 58.68744, 58.71812, 58.74852, 58.77864, 
    58.80849, 58.83805, 58.86733, 58.89633, 58.92505, 58.95348, 58.98163, 
    59.00949, 59.03706, 59.06435, 59.09135, 59.11806, 59.14449, 59.17062, 
    59.19646, 59.22201, 59.24727, 59.27223, 59.2969, 59.32128, 59.34536, 
    59.36914, 59.39263, 59.41582, 59.43871, 59.4613, 59.48359, 59.50558, 
    59.52728, 59.54866, 59.56975, 59.59054, 59.61102, 59.6312, 59.65107, 
    59.67064, 59.6899, 59.70885, 59.7275, 59.74583, 59.76387, 59.78159, 
    59.799, 59.8161, 59.8329, 59.84938, 59.86555, 59.8814, 59.89695, 
    59.91218, 59.9271, 59.9417, 59.95599, 59.96997, 59.98363, 59.99697, 
    60.01, 60.02271, 60.0351, 60.04718, 60.05894, 60.07037, 60.0815, 60.0923, 
    60.10278, 60.11294, 60.12279, 60.13231, 60.14151, 60.15039, 60.15895, 
    60.16719, 60.1751, 60.1827, 60.18997, 60.19691, 60.20354, 60.20984, 
    60.21582, 60.22148, 60.22681, 60.23182, 60.2365, 60.24086, 60.2449, 
    60.24861, 60.252, 60.25506, 60.2578, 60.26021, 60.2623, 60.26406, 
    60.2655, 60.26661, 60.2674, 60.26786, 60.268, 60.26781, 60.2673, 
    60.26646, 60.26529, 60.26381, 60.26199, 60.25985, 60.25739, 60.2546, 
    60.25148, 60.24805, 60.24429, 60.2402, 60.23579, 60.23105, 60.22599, 
    60.22061, 60.2149, 60.20887, 60.20251, 60.19584, 60.18884, 60.18151, 
    60.17387, 60.1659, 60.15762, 60.14901, 60.14008, 60.13082, 60.12125, 
    60.11136, 60.10114, 60.09061, 60.07976, 60.06859, 60.0571, 60.04529, 
    60.03316, 60.02072, 60.00796, 59.99488, 59.98149, 59.96778, 59.95375, 
    59.93941, 59.92476, 59.90979, 59.89451, 59.87892, 59.86301, 59.84679, 
    59.83026, 59.81342, 59.79627, 59.7788, 59.76104, 59.74295, 59.72457, 
    59.70587, 59.68687, 59.66756, 59.64795, 59.62803, 59.6078, 59.58727, 
    59.56644, 59.5453, 59.52386, 59.50212, 59.48008, 59.45774, 59.4351, 
    59.41217, 59.38893, 59.3654, 59.34157, 59.31744, 59.29302, 59.2683, 
    59.24329, 59.21799, 59.19239, 59.16651, 59.14033, 59.11386, 59.0871, 
    59.06005, 59.03272, 59.0051, 58.9772, 58.949, 58.92052, 58.89176, 
    58.86272, 58.83339, 58.80378, 58.7739, 58.74373, 58.71328, 58.68256, 
    58.65155, 58.62027, 58.58872, 58.55689, 58.52479, 58.49241, 58.45976, 
    58.42684, 58.39365, 58.3602, 58.32647, 58.29247, 58.25821, 58.22368, 
    58.18888, 58.15383, 58.1185, 58.08292, 58.04707, 58.01097, 57.9746, 
    57.93798, 57.9011, 57.86396, 57.82656, 57.78891, 57.75101, 57.71285, 
    57.67444, 57.63578, 57.59686, 57.5577, 57.51829, 57.47863, 57.43872, 
    57.39857, 57.35818, 57.31754, 57.27666, 57.23553, 57.19416, 57.15256, 
    57.11071, 57.06863, 57.02631, 56.98375, 56.94095, 56.89793, 56.85466, 
    56.81117, 56.76744, 56.72348, 56.6793, 56.63488, 56.59024, 56.54536, 
    56.50027, 56.45495, 56.4094, 56.36363, 56.31764, 56.27142, 56.22499, 
    56.17834, 56.13147, 56.08438, 56.03707, 55.98955, 55.94181, 55.89386, 
    55.8457,
  50.65811, 50.72233, 50.78642, 50.85037, 50.91419, 50.97786, 51.0414, 
    51.1048, 51.16806, 51.23119, 51.29417, 51.35701, 51.4197, 51.48226, 
    51.54467, 51.60693, 51.66905, 51.73102, 51.79285, 51.85453, 51.91606, 
    51.97744, 52.03867, 52.09975, 52.16068, 52.22146, 52.28209, 52.34256, 
    52.40287, 52.46303, 52.52304, 52.58288, 52.64257, 52.7021, 52.76147, 
    52.82069, 52.87974, 52.93863, 52.99735, 53.05592, 53.11431, 53.17255, 
    53.23061, 53.28851, 53.34624, 53.40381, 53.4612, 53.51843, 53.57549, 
    53.63237, 53.68908, 53.74561, 53.80198, 53.85816, 53.91417, 53.97001, 
    54.02566, 54.08114, 54.13644, 54.19156, 54.24649, 54.30125, 54.35582, 
    54.4102, 54.46441, 54.51842, 54.57225, 54.62589, 54.67935, 54.73261, 
    54.78569, 54.83857, 54.89126, 54.94376, 54.99607, 55.04818, 55.10009, 
    55.15181, 55.20333, 55.25465, 55.30578, 55.3567, 55.40742, 55.45794, 
    55.50826, 55.55837, 55.60828, 55.65799, 55.70748, 55.75677, 55.80585, 
    55.85472, 55.90338, 55.95183, 56.00006, 56.04809, 56.0959, 56.14349, 
    56.19087, 56.23803, 56.28498, 56.3317, 56.3782, 56.42449, 56.47055, 
    56.51639, 56.56201, 56.6074, 56.65257, 56.69751, 56.74222, 56.7867, 
    56.83096, 56.87498, 56.91877, 56.96233, 57.00566, 57.04876, 57.09162, 
    57.13424, 57.17662, 57.21877, 57.26068, 57.30235, 57.34378, 57.38497, 
    57.42591, 57.46662, 57.50708, 57.54729, 57.58725, 57.62697, 57.66644, 
    57.70566, 57.74463, 57.78335, 57.82182, 57.86003, 57.89799, 57.9357, 
    57.97315, 58.01034, 58.04728, 58.08396, 58.12038, 58.15653, 58.19243, 
    58.22807, 58.26344, 58.29855, 58.33339, 58.36797, 58.40228, 58.43632, 
    58.4701, 58.5036, 58.53683, 58.5698, 58.60249, 58.63491, 58.66706, 
    58.69893, 58.73053, 58.76184, 58.79289, 58.82365, 58.85414, 58.88435, 
    58.91427, 58.94392, 58.97328, 59.00236, 59.03115, 59.05966, 59.08789, 
    59.11583, 59.14348, 59.17085, 59.19792, 59.2247, 59.2512, 59.27741, 
    59.30332, 59.32894, 59.35427, 59.37931, 59.40405, 59.42849, 59.45264, 
    59.47649, 59.50004, 59.5233, 59.54625, 59.56891, 59.59127, 59.61332, 
    59.63508, 59.65653, 59.67768, 59.69852, 59.71906, 59.7393, 59.75923, 
    59.77885, 59.79817, 59.81718, 59.83588, 59.85427, 59.87236, 59.89013, 
    59.9076, 59.92475, 59.94159, 59.95812, 59.97434, 59.99024, 60.00583, 
    60.02111, 60.03607, 60.05072, 60.06505, 60.07907, 60.09277, 60.10615, 
    60.11922, 60.13197, 60.1444, 60.15651, 60.1683, 60.17978, 60.19093, 
    60.20177, 60.21228, 60.22247, 60.23235, 60.2419, 60.25113, 60.26003, 
    60.26862, 60.27688, 60.28482, 60.29244, 60.29973, 60.3067, 60.31335, 
    60.31967, 60.32566, 60.33134, 60.33669, 60.34171, 60.34641, 60.35078, 
    60.35483, 60.35855, 60.36195, 60.36502, 60.36777, 60.37019, 60.37228, 
    60.37405, 60.37549, 60.37661, 60.3774, 60.37786, 60.378, 60.37781, 
    60.3773, 60.37645, 60.37529, 60.37379, 60.37197, 60.36983, 60.36736, 
    60.36456, 60.36143, 60.35799, 60.35421, 60.35011, 60.34569, 60.34094, 
    60.33586, 60.33046, 60.32474, 60.31869, 60.31232, 60.30562, 60.2986, 
    60.29125, 60.28358, 60.2756, 60.26728, 60.25864, 60.24969, 60.24041, 
    60.2308, 60.22088, 60.21064, 60.20007, 60.18919, 60.17798, 60.16646, 
    60.15461, 60.14245, 60.12997, 60.11717, 60.10406, 60.09062, 60.07687, 
    60.06281, 60.04842, 60.03373, 60.01871, 60.00339, 59.98775, 59.97179, 
    59.95553, 59.93895, 59.92206, 59.90485, 59.88734, 59.86952, 59.85138, 
    59.83294, 59.81419, 59.79514, 59.77577, 59.7561, 59.73612, 59.71584, 
    59.69524, 59.67435, 59.65316, 59.63166, 59.60986, 59.58775, 59.56535, 
    59.54264, 59.51964, 59.49634, 59.47274, 59.44884, 59.42464, 59.40015, 
    59.37537, 59.35028, 59.32491, 59.29924, 59.27328, 59.24703, 59.22049, 
    59.19366, 59.16653, 59.13913, 59.11143, 59.08344, 59.05517, 59.02662, 
    58.99778, 58.96865, 58.93924, 58.90955, 58.87959, 58.84933, 58.81881, 
    58.78799, 58.75691, 58.72555, 58.6939, 58.66199, 58.6298, 58.59734, 
    58.56461, 58.5316, 58.49832, 58.46477, 58.43095, 58.39687, 58.36251, 
    58.3279, 58.29301, 58.25786, 58.22245, 58.18677, 58.15083, 58.11463, 
    58.07817, 58.04145, 58.00448, 57.96724, 57.92975, 57.89201, 57.854, 
    57.81575, 57.77724, 57.73848, 57.69947, 57.66021, 57.6207, 57.58095, 
    57.54094, 57.50069, 57.46019, 57.41946, 57.37847, 57.33725, 57.29578, 
    57.25407, 57.21212, 57.16994, 57.12751, 57.08485, 57.04196, 56.99883, 
    56.95546, 56.91186, 56.86803, 56.82397, 56.77968, 56.73516, 56.69041, 
    56.64544, 56.60023, 56.55481, 56.50916, 56.46328, 56.41718, 56.37086, 
    56.32433, 56.27757, 56.23059, 56.18339, 56.13598, 56.08835, 56.04051, 
    55.99245, 55.94418,
  50.74665, 50.81098, 50.87516, 50.93922, 51.00313, 51.06691, 51.13055, 
    51.19405, 51.25742, 51.32064, 51.38372, 51.44667, 51.50946, 51.57212, 
    51.63463, 51.697, 51.75922, 51.8213, 51.88323, 51.94501, 52.00665, 
    52.06813, 52.12947, 52.19066, 52.25169, 52.31257, 52.3733, 52.43388, 
    52.4943, 52.55457, 52.61468, 52.67463, 52.73442, 52.79406, 52.85354, 
    52.91286, 52.97201, 53.03101, 53.08984, 53.14851, 53.20702, 53.26535, 
    53.32353, 53.38154, 53.43938, 53.49705, 53.55455, 53.61189, 53.66905, 
    53.72604, 53.78286, 53.8395, 53.89597, 53.95226, 54.00838, 54.06432, 
    54.12009, 54.17567, 54.23108, 54.2863, 54.34135, 54.39621, 54.45089, 
    54.50539, 54.5597, 54.61382, 54.66776, 54.72151, 54.77508, 54.82845, 
    54.88163, 54.93462, 54.98743, 55.04003, 55.09245, 55.14466, 55.19669, 
    55.24852, 55.30014, 55.35158, 55.40281, 55.45384, 55.50467, 55.5553, 
    55.60572, 55.65594, 55.70596, 55.75577, 55.80538, 55.85477, 55.90396, 
    55.95294, 56.00171, 56.05026, 56.09861, 56.14674, 56.19466, 56.24236, 
    56.28984, 56.33711, 56.38416, 56.43099, 56.4776, 56.52399, 56.57016, 
    56.61611, 56.66183, 56.70732, 56.7526, 56.79764, 56.84246, 56.88705, 
    56.93141, 56.97554, 57.01943, 57.0631, 57.10653, 57.14973, 57.19269, 
    57.23541, 57.2779, 57.32015, 57.36216, 57.40394, 57.44547, 57.48676, 
    57.5278, 57.5686, 57.60916, 57.64947, 57.68954, 57.72935, 57.76892, 
    57.80824, 57.84731, 57.88613, 57.92469, 57.96301, 58.00106, 58.03886, 
    58.07641, 58.1137, 58.15073, 58.1875, 58.22402, 58.26027, 58.29626, 
    58.33199, 58.36745, 58.40265, 58.43758, 58.47225, 58.50666, 58.54079, 
    58.57465, 58.60825, 58.64157, 58.67463, 58.70741, 58.73991, 58.77214, 
    58.8041, 58.83578, 58.86719, 58.89831, 58.92916, 58.95973, 58.99002, 
    59.02003, 59.04975, 59.0792, 59.10836, 59.13723, 59.16582, 59.19412, 
    59.22214, 59.24987, 59.27731, 59.30446, 59.33133, 59.35789, 59.38417, 
    59.41016, 59.43586, 59.46125, 59.48636, 59.51117, 59.53569, 59.5599, 
    59.58382, 59.60744, 59.63076, 59.65379, 59.67651, 59.69893, 59.72105, 
    59.74287, 59.76438, 59.78559, 59.8065, 59.8271, 59.84739, 59.86738, 
    59.88706, 59.90643, 59.9255, 59.94426, 59.9627, 59.98084, 59.99866, 
    60.01618, 60.03339, 60.05028, 60.06686, 60.08312, 60.09907, 60.11471, 
    60.13003, 60.14504, 60.15973, 60.17411, 60.18816, 60.2019, 60.21533, 
    60.22844, 60.24122, 60.25369, 60.26584, 60.27767, 60.28917, 60.30036, 
    60.31123, 60.32178, 60.332, 60.3419, 60.35148, 60.36074, 60.36967, 
    60.37828, 60.38657, 60.39454, 60.40218, 60.40949, 60.41648, 60.42315, 
    60.42949, 60.4355, 60.4412, 60.44656, 60.4516, 60.45631, 60.4607, 
    60.46476, 60.46849, 60.4719, 60.47498, 60.47774, 60.48016, 60.48227, 
    60.48404, 60.48549, 60.4866, 60.4874, 60.48786, 60.488, 60.48781, 
    60.48729, 60.48645, 60.48528, 60.48378, 60.48196, 60.4798, 60.47732, 
    60.47452, 60.47139, 60.46793, 60.46414, 60.46003, 60.45559, 60.45082, 
    60.44573, 60.44032, 60.43457, 60.42851, 60.42212, 60.4154, 60.40836, 
    60.40099, 60.3933, 60.38528, 60.37695, 60.36828, 60.35929, 60.34999, 
    60.34036, 60.3304, 60.32013, 60.30953, 60.29861, 60.28738, 60.27582, 
    60.26394, 60.25174, 60.23922, 60.22638, 60.21323, 60.19975, 60.18596, 
    60.17185, 60.15743, 60.14269, 60.12763, 60.11226, 60.09657, 60.08057, 
    60.06425, 60.04763, 60.03069, 60.01343, 59.99586, 59.97799, 59.9598, 
    59.94131, 59.9225, 59.90339, 59.88396, 59.86423, 59.8442, 59.82386, 
    59.80321, 59.78225, 59.761, 59.73943, 59.71757, 59.6954, 59.67294, 
    59.65017, 59.62709, 59.60373, 59.58006, 59.55609, 59.53183, 59.50727, 
    59.48241, 59.45726, 59.43181, 59.40607, 59.38004, 59.35371, 59.3271, 
    59.30019, 59.27299, 59.2455, 59.21773, 59.18967, 59.16132, 59.13268, 
    59.10376, 59.07456, 59.04507, 59.0153, 58.98525, 58.95491, 58.9243, 
    58.89341, 58.86224, 58.83079, 58.79906, 58.76706, 58.73479, 58.70224, 
    58.66941, 58.63632, 58.60295, 58.56931, 58.53541, 58.50123, 58.46679, 
    58.43208, 58.3971, 58.36186, 58.32635, 58.29058, 58.25455, 58.21826, 
    58.18171, 58.14489, 58.10782, 58.07049, 58.0329, 57.99506, 57.95696, 
    57.91861, 57.88, 57.84115, 57.80204, 57.76268, 57.72307, 57.68322, 
    57.64311, 57.60276, 57.56216, 57.52132, 57.48024, 57.43892, 57.39735, 
    57.35553, 57.31348, 57.2712, 57.22867, 57.18591, 57.14291, 57.09967, 
    57.05621, 57.0125, 56.96857, 56.9244, 56.88001, 56.83538, 56.79053, 
    56.74545, 56.70014, 56.65461, 56.60885, 56.56287, 56.51667, 56.47025, 
    56.4236, 56.37673, 56.32965, 56.28234, 56.23483, 56.18709, 56.13914, 
    56.09098, 56.0426,
  50.83511, 50.89953, 50.96382, 51.02797, 51.09199, 51.15587, 51.21961, 
    51.28322, 51.34668, 51.41001, 51.47319, 51.53624, 51.59914, 51.6619, 
    51.72451, 51.78699, 51.84931, 51.91149, 51.97353, 52.03542, 52.09715, 
    52.15874, 52.22018, 52.28148, 52.34261, 52.4036, 52.46444, 52.52512, 
    52.58564, 52.64602, 52.70623, 52.76629, 52.82619, 52.88593, 52.94552, 
    53.00494, 53.06421, 53.12331, 53.18225, 53.24102, 53.29964, 53.35809, 
    53.41637, 53.47448, 53.53243, 53.59021, 53.64782, 53.70526, 53.76253, 
    53.81963, 53.87655, 53.9333, 53.98988, 54.04629, 54.10252, 54.15857, 
    54.21444, 54.27013, 54.32565, 54.38098, 54.43613, 54.4911, 54.54589, 
    54.6005, 54.65492, 54.70915, 54.7632, 54.81706, 54.87073, 54.92421, 
    54.9775, 55.03061, 55.08352, 55.13623, 55.18876, 55.24109, 55.29322, 
    55.34515, 55.39689, 55.44843, 55.49977, 55.55091, 55.60185, 55.65259, 
    55.70312, 55.75345, 55.80358, 55.8535, 55.90321, 55.95271, 56.00201, 
    56.0511, 56.09997, 56.14864, 56.19709, 56.24533, 56.29335, 56.34116, 
    56.38875, 56.43613, 56.48328, 56.53022, 56.57694, 56.62344, 56.66971, 
    56.71576, 56.76159, 56.80719, 56.85257, 56.89772, 56.94265, 56.98734, 
    57.0318, 57.07603, 57.12004, 57.16381, 57.20734, 57.25064, 57.29371, 
    57.33654, 57.37913, 57.42148, 57.4636, 57.50547, 57.5471, 57.58849, 
    57.62964, 57.67054, 57.7112, 57.75161, 57.79178, 57.8317, 57.87136, 
    57.91078, 57.94995, 57.98886, 58.02753, 58.06593, 58.10409, 58.14199, 
    58.17963, 58.21702, 58.25414, 58.29101, 58.32762, 58.36396, 58.40005, 
    58.43587, 58.47143, 58.50672, 58.54174, 58.57651, 58.611, 58.64522, 
    58.67918, 58.71286, 58.74627, 58.77942, 58.81228, 58.84488, 58.8772, 
    58.90924, 58.94101, 58.9725, 59.00371, 59.03464, 59.0653, 59.09566, 
    59.12576, 59.15556, 59.18509, 59.21433, 59.24329, 59.27195, 59.30033, 
    59.32843, 59.35624, 59.38375, 59.41098, 59.43792, 59.46457, 59.49092, 
    59.51698, 59.54275, 59.56822, 59.5934, 59.61828, 59.64286, 59.66715, 
    59.69114, 59.71482, 59.73821, 59.7613, 59.78409, 59.80658, 59.82876, 
    59.85064, 59.87222, 59.89349, 59.91446, 59.93512, 59.95547, 59.97551, 
    59.99525, 60.01468, 60.03381, 60.05262, 60.07112, 60.08931, 60.10719, 
    60.12476, 60.14201, 60.15895, 60.17558, 60.19189, 60.2079, 60.22358, 
    60.23895, 60.254, 60.26873, 60.28315, 60.29725, 60.31104, 60.3245, 
    60.33765, 60.35047, 60.36298, 60.37516, 60.38702, 60.39857, 60.40979, 
    60.42069, 60.43127, 60.44152, 60.45145, 60.46106, 60.47035, 60.47931, 
    60.48795, 60.49626, 60.50425, 60.51191, 60.51925, 60.52626, 60.53295, 
    60.53931, 60.54535, 60.55105, 60.55643, 60.56149, 60.56622, 60.57061, 
    60.57469, 60.57843, 60.58185, 60.58494, 60.58771, 60.59014, 60.59225, 
    60.59402, 60.59548, 60.5966, 60.59739, 60.59786, 60.598, 60.59781, 
    60.59729, 60.59644, 60.59527, 60.59377, 60.59193, 60.58978, 60.58729, 
    60.58448, 60.58133, 60.57787, 60.57407, 60.56994, 60.56549, 60.56071, 
    60.5556, 60.55017, 60.54441, 60.53833, 60.53191, 60.52518, 60.51811, 
    60.51072, 60.50301, 60.49497, 60.4866, 60.47792, 60.4689, 60.45956, 
    60.44991, 60.43992, 60.42962, 60.41899, 60.40804, 60.39676, 60.38517, 
    60.37325, 60.36102, 60.34846, 60.33559, 60.32239, 60.30888, 60.29504, 
    60.2809, 60.26643, 60.25164, 60.23654, 60.22112, 60.20539, 60.18933, 
    60.17297, 60.1563, 60.13931, 60.122, 60.10438, 60.08645, 60.06821, 
    60.04966, 60.0308, 60.01163, 59.99215, 59.97237, 59.95227, 59.93187, 
    59.91116, 59.89014, 59.86882, 59.8472, 59.82527, 59.80304, 59.78051, 
    59.75767, 59.73454, 59.7111, 59.68736, 59.66333, 59.63899, 59.61436, 
    59.58944, 59.56421, 59.53869, 59.51288, 59.48677, 59.46037, 59.43368, 
    59.4067, 59.37942, 59.35186, 59.32401, 59.29586, 59.26744, 59.23872, 
    59.20972, 59.18044, 59.15087, 59.12102, 59.09088, 59.06047, 59.02977, 
    58.99879, 58.96754, 58.936, 58.90419, 58.8721, 58.83974, 58.8071, 
    58.77419, 58.741, 58.70755, 58.67382, 58.63983, 58.60556, 58.57103, 
    58.53622, 58.50116, 58.46582, 58.43022, 58.39436, 58.35823, 58.32185, 
    58.28519, 58.24829, 58.21112, 58.17369, 58.13601, 58.09807, 58.05988, 
    58.02143, 57.98272, 57.94377, 57.90456, 57.8651, 57.8254, 57.78544, 
    57.74524, 57.70478, 57.66409, 57.62315, 57.58196, 57.54053, 57.49886, 
    57.45695, 57.4148, 57.37241, 57.32978, 57.28691, 57.24381, 57.20047, 
    57.1569, 57.11309, 57.06905, 57.02478, 56.98029, 56.93555, 56.89059, 
    56.84541, 56.8, 56.75436, 56.7085, 56.66241, 56.6161, 56.56956, 56.52281, 
    56.47584, 56.42865, 56.38124, 56.33361, 56.28577, 56.23771, 56.18944, 
    56.14095,
  50.92347, 50.98799, 51.05238, 51.11663, 51.18076, 51.24474, 51.30858, 
    51.37229, 51.43586, 51.49928, 51.56257, 51.62572, 51.68872, 51.75159, 
    51.8143, 51.87688, 51.93931, 52.00159, 52.06373, 52.12572, 52.18757, 
    52.24926, 52.31081, 52.3722, 52.43345, 52.49454, 52.55548, 52.61627, 
    52.6769, 52.73738, 52.7977, 52.85786, 52.91787, 52.97772, 53.03741, 
    53.09695, 53.15631, 53.21552, 53.27457, 53.33345, 53.39217, 53.45073, 
    53.50912, 53.56734, 53.6254, 53.68328, 53.741, 53.79855, 53.85593, 
    53.91314, 53.97017, 54.02703, 54.08372, 54.14023, 54.19657, 54.25273, 
    54.30871, 54.36451, 54.42014, 54.47558, 54.53084, 54.58592, 54.64082, 
    54.69553, 54.75006, 54.80441, 54.85856, 54.91253, 54.96631, 55.01991, 
    55.07331, 55.12652, 55.17954, 55.23236, 55.285, 55.33743, 55.38968, 
    55.44172, 55.49357, 55.54522, 55.59667, 55.64791, 55.69896, 55.74981, 
    55.80045, 55.85089, 55.90113, 55.95116, 56.00098, 56.05059, 56.09999, 
    56.14919, 56.19817, 56.24695, 56.29551, 56.34385, 56.39199, 56.4399, 
    56.4876, 56.53508, 56.58235, 56.62939, 56.67622, 56.72282, 56.76921, 
    56.81536, 56.8613, 56.90701, 56.95249, 56.99775, 57.04277, 57.08757, 
    57.13214, 57.17648, 57.22059, 57.26446, 57.3081, 57.35151, 57.39468, 
    57.43761, 57.4803, 57.52276, 57.56498, 57.60696, 57.64869, 57.69018, 
    57.73143, 57.77243, 57.81319, 57.85371, 57.89397, 57.93399, 57.97375, 
    58.01328, 58.05254, 58.09156, 58.13032, 58.16882, 58.20708, 58.24507, 
    58.28281, 58.32029, 58.35752, 58.39448, 58.43118, 58.46762, 58.5038, 
    58.53971, 58.57537, 58.61075, 58.64587, 58.68072, 58.71531, 58.74962, 
    58.78367, 58.81744, 58.85094, 58.88417, 58.91713, 58.94981, 58.98222, 
    59.01435, 59.0462, 59.07778, 59.10908, 59.14009, 59.17083, 59.20129, 
    59.23146, 59.26135, 59.29095, 59.32028, 59.34931, 59.37806, 59.40652, 
    59.4347, 59.46258, 59.49018, 59.51748, 59.5445, 59.57122, 59.59764, 
    59.62378, 59.64962, 59.67516, 59.70041, 59.72536, 59.75002, 59.77438, 
    59.79843, 59.82219, 59.84565, 59.8688, 59.89165, 59.91421, 59.93645, 
    59.9584, 59.98004, 60.00137, 60.0224, 60.04312, 60.06353, 60.08364, 
    60.10344, 60.12292, 60.1421, 60.16097, 60.17953, 60.19777, 60.21571, 
    60.23332, 60.25063, 60.26762, 60.2843, 60.30066, 60.31671, 60.33244, 
    60.34785, 60.36295, 60.37773, 60.39219, 60.40634, 60.42016, 60.43367, 
    60.44685, 60.45971, 60.47226, 60.48448, 60.49638, 60.50796, 60.51921, 
    60.53015, 60.54076, 60.55104, 60.561, 60.57064, 60.57996, 60.58895, 
    60.59761, 60.60595, 60.61396, 60.62165, 60.62901, 60.63604, 60.64275, 
    60.64913, 60.65518, 60.66091, 60.66631, 60.67138, 60.67612, 60.68053, 
    60.68462, 60.68837, 60.6918, 60.6949, 60.69767, 60.70012, 60.70223, 
    60.70401, 60.70547, 60.7066, 60.70739, 60.70786, 60.708, 60.70781, 
    60.70729, 60.70644, 60.70526, 60.70375, 60.70192, 60.69975, 60.69726, 
    60.69444, 60.69128, 60.6878, 60.68399, 60.67986, 60.67539, 60.67059, 
    60.66547, 60.66002, 60.65425, 60.64814, 60.64171, 60.63495, 60.62786, 
    60.62045, 60.61272, 60.60465, 60.59626, 60.58755, 60.57851, 60.56914, 
    60.55945, 60.54944, 60.5391, 60.52844, 60.51746, 60.50615, 60.49452, 
    60.48257, 60.47029, 60.4577, 60.44479, 60.43155, 60.418, 60.40412, 
    60.38993, 60.37542, 60.36058, 60.34544, 60.32998, 60.31419, 60.2981, 
    60.28168, 60.26495, 60.24791, 60.23056, 60.21289, 60.19491, 60.17661, 
    60.158, 60.13909, 60.11986, 60.10033, 60.08048, 60.06033, 60.03986, 
    60.01909, 59.99802, 59.97663, 59.95495, 59.93296, 59.91066, 59.88806, 
    59.86516, 59.84196, 59.81845, 59.79465, 59.77054, 59.74614, 59.72144, 
    59.69644, 59.67114, 59.64555, 59.61967, 59.59349, 59.56701, 59.54024, 
    59.51318, 59.48583, 59.45819, 59.43026, 59.40204, 59.37354, 59.34474, 
    59.31566, 59.28629, 59.25664, 59.22671, 59.19649, 59.16599, 59.13521, 
    59.10415, 59.0728, 59.04118, 59.00928, 58.97711, 58.94466, 58.91194, 
    58.87894, 58.84566, 58.81212, 58.7783, 58.74421, 58.70985, 58.67523, 
    58.64034, 58.60517, 58.56974, 58.53405, 58.4981, 58.46188, 58.42539, 
    58.38865, 58.35165, 58.31438, 58.27686, 58.23908, 58.20104, 58.16275, 
    58.1242, 58.0854, 58.04634, 58.00704, 57.96748, 57.92768, 57.88762, 
    57.84731, 57.80676, 57.76596, 57.72492, 57.68364, 57.64211, 57.60033, 
    57.55832, 57.51606, 57.47357, 57.43084, 57.38786, 57.34466, 57.30122, 
    57.25754, 57.21363, 57.16948, 57.12511, 57.08051, 57.03567, 56.9906, 
    56.94531, 56.89979, 56.85405, 56.80808, 56.76188, 56.71547, 56.66883, 
    56.62197, 56.57489, 56.52759, 56.48007, 56.43234, 56.38439, 56.33622, 
    56.28784, 56.23925,
  51.01173, 51.07636, 51.14085, 51.20521, 51.26943, 51.33351, 51.39746, 
    51.46127, 51.52494, 51.58847, 51.65186, 51.71511, 51.77822, 51.84118, 
    51.90401, 51.96669, 52.02922, 52.09161, 52.15385, 52.21595, 52.2779, 
    52.33969, 52.40134, 52.46284, 52.5242, 52.5854, 52.64644, 52.70733, 
    52.76807, 52.82866, 52.88908, 52.94936, 53.00947, 53.06943, 53.12922, 
    53.18886, 53.24834, 53.30766, 53.36681, 53.4258, 53.48463, 53.54329, 
    53.60179, 53.66012, 53.71828, 53.77628, 53.83411, 53.89177, 53.94925, 
    54.00657, 54.06371, 54.12068, 54.17747, 54.2341, 54.29054, 54.34681, 
    54.4029, 54.45881, 54.51455, 54.5701, 54.62547, 54.68066, 54.73567, 
    54.79049, 54.84513, 54.89959, 54.95385, 55.00793, 55.06182, 55.11552, 
    55.16904, 55.22235, 55.27549, 55.32842, 55.38116, 55.43371, 55.48606, 
    55.53822, 55.59017, 55.64193, 55.69349, 55.74485, 55.79601, 55.84697, 
    55.89772, 55.94827, 55.99861, 56.04875, 56.09868, 56.1484, 56.19791, 
    56.24722, 56.29631, 56.34519, 56.39386, 56.44232, 56.49056, 56.53858, 
    56.58639, 56.63398, 56.68135, 56.72851, 56.77544, 56.82215, 56.86864, 
    56.91491, 56.96095, 57.00676, 57.05235, 57.09772, 57.14285, 57.18776, 
    57.23243, 57.27687, 57.32109, 57.36507, 57.40881, 57.45232, 57.49559, 
    57.53863, 57.58143, 57.62399, 57.66631, 57.70839, 57.75023, 57.79182, 
    57.83317, 57.87428, 57.91514, 57.95575, 57.99612, 58.03624, 58.07611, 
    58.11572, 58.15509, 58.1942, 58.23306, 58.27167, 58.31002, 58.34811, 
    58.38595, 58.42353, 58.46085, 58.49791, 58.53471, 58.57124, 58.60751, 
    58.64352, 58.67927, 58.71475, 58.74996, 58.7849, 58.81958, 58.85399, 
    58.88812, 58.92199, 58.95558, 58.9889, 59.02195, 59.05472, 59.08721, 
    59.11943, 59.15137, 59.18303, 59.21442, 59.24552, 59.27634, 59.30688, 
    59.33714, 59.36711, 59.3968, 59.4262, 59.45532, 59.48415, 59.51269, 
    59.54094, 59.5689, 59.59658, 59.62396, 59.65105, 59.67785, 59.70435, 
    59.73056, 59.75647, 59.78209, 59.80741, 59.83244, 59.85716, 59.88159, 
    59.90571, 59.92954, 59.95306, 59.97629, 59.99921, 60.02182, 60.04414, 
    60.06614, 60.08784, 60.10924, 60.13033, 60.15112, 60.17159, 60.19175, 
    60.21161, 60.23116, 60.25039, 60.26931, 60.28792, 60.30622, 60.32421, 
    60.34188, 60.35924, 60.37628, 60.39301, 60.40942, 60.42552, 60.4413, 
    60.45676, 60.4719, 60.48672, 60.50123, 60.51542, 60.52928, 60.54282, 
    60.55605, 60.56895, 60.58154, 60.59379, 60.60573, 60.61734, 60.62864, 
    60.6396, 60.65024, 60.66056, 60.67056, 60.68022, 60.68956, 60.69858, 
    60.70727, 60.71563, 60.72367, 60.73138, 60.73877, 60.74582, 60.75255, 
    60.75895, 60.76502, 60.77076, 60.77618, 60.78126, 60.78602, 60.79045, 
    60.79454, 60.79831, 60.80175, 60.80486, 60.80764, 60.81009, 60.81221, 
    60.814, 60.81546, 60.81659, 60.81739, 60.81786, 60.818, 60.81781, 
    60.81729, 60.81643, 60.81525, 60.81374, 60.8119, 60.80973, 60.80722, 
    60.80439, 60.80123, 60.79774, 60.79392, 60.78977, 60.78529, 60.78048, 
    60.77534, 60.76987, 60.76408, 60.75796, 60.75151, 60.74472, 60.73762, 
    60.73018, 60.72242, 60.71433, 60.70592, 60.69717, 60.68811, 60.67871, 
    60.66899, 60.65895, 60.64858, 60.63789, 60.62687, 60.61553, 60.60386, 
    60.59188, 60.57957, 60.56693, 60.55398, 60.5407, 60.52711, 60.51319, 
    60.49895, 60.4844, 60.46952, 60.45433, 60.43882, 60.42299, 60.40685, 
    60.39038, 60.37361, 60.35651, 60.33911, 60.32138, 60.30335, 60.285, 
    60.26634, 60.24737, 60.22808, 60.20849, 60.18858, 60.16837, 60.14785, 
    60.12702, 60.10588, 60.08443, 60.06268, 60.04063, 60.01826, 59.9956, 
    59.97263, 59.94936, 59.92579, 59.90192, 59.87774, 59.85327, 59.8285, 
    59.80342, 59.77806, 59.75239, 59.72643, 59.70018, 59.67363, 59.64679, 
    59.61965, 59.59222, 59.5645, 59.53649, 59.50819, 59.47961, 59.45073, 
    59.42157, 59.39212, 59.36239, 59.33237, 59.30207, 59.27148, 59.24062, 
    59.20947, 59.17804, 59.14634, 59.11435, 59.08209, 59.04955, 59.01674, 
    58.98365, 58.95029, 58.91665, 58.88274, 58.84856, 58.81411, 58.7794, 
    58.74441, 58.70915, 58.67363, 58.63784, 58.6018, 58.56548, 58.5289, 
    58.49206, 58.45496, 58.4176, 58.37998, 58.34211, 58.30397, 58.26558, 
    58.22693, 58.18803, 58.14888, 58.10947, 58.06982, 58.02991, 57.98975, 
    57.94934, 57.90869, 57.86779, 57.82665, 57.78526, 57.74363, 57.70175, 
    57.65963, 57.61728, 57.57468, 57.53184, 57.48877, 57.44545, 57.40191, 
    57.35812, 57.31411, 57.26986, 57.22538, 57.18067, 57.13573, 57.09056, 
    57.04516, 56.99953, 56.95368, 56.9076, 56.8613, 56.81478, 56.76803, 
    56.72106, 56.67387, 56.62647, 56.57884, 56.531, 56.48294, 56.43467, 
    56.38618, 56.33747,
  51.09991, 51.16463, 51.22923, 51.29369, 51.35801, 51.4222, 51.48624, 
    51.55016, 51.61393, 51.67756, 51.74105, 51.80441, 51.86762, 51.93069, 
    51.99361, 52.0564, 52.11904, 52.18153, 52.24388, 52.30608, 52.36813, 
    52.43004, 52.49179, 52.5534, 52.61486, 52.67616, 52.73731, 52.79831, 
    52.85915, 52.91985, 52.98038, 53.04076, 53.10098, 53.16105, 53.22095, 
    53.28069, 53.34028, 53.3997, 53.45897, 53.51807, 53.577, 53.63577, 
    53.69438, 53.75282, 53.81109, 53.86919, 53.92713, 53.9849, 54.04249, 
    54.09991, 54.15717, 54.21425, 54.27115, 54.32788, 54.38444, 54.44081, 
    54.49702, 54.55304, 54.60888, 54.66454, 54.72002, 54.77533, 54.83044, 
    54.88538, 54.94012, 54.99469, 55.04906, 55.10325, 55.15726, 55.21107, 
    55.26469, 55.31812, 55.37136, 55.4244, 55.47726, 55.52991, 55.58237, 
    55.63464, 55.68671, 55.73858, 55.79025, 55.84172, 55.89299, 55.94405, 
    55.99492, 56.04557, 56.09602, 56.14627, 56.19631, 56.24614, 56.29577, 
    56.34518, 56.39438, 56.44337, 56.49215, 56.54072, 56.58907, 56.6372, 
    56.68512, 56.73281, 56.7803, 56.82756, 56.8746, 56.92142, 56.96801, 
    57.01439, 57.06054, 57.10646, 57.15216, 57.19763, 57.24287, 57.28788, 
    57.33266, 57.37721, 57.42153, 57.46561, 57.50946, 57.55308, 57.59646, 
    57.6396, 57.6825, 57.72517, 57.76759, 57.80978, 57.85172, 57.89341, 
    57.93487, 57.97607, 58.01704, 58.05775, 58.09822, 58.13844, 58.17841, 
    58.21813, 58.2576, 58.29681, 58.33577, 58.37447, 58.41292, 58.45111, 
    58.48905, 58.52672, 58.56414, 58.6013, 58.63819, 58.67482, 58.71119, 
    58.7473, 58.78313, 58.81871, 58.85401, 58.88905, 58.92382, 58.95832, 
    58.99255, 59.0265, 59.06018, 59.09359, 59.12673, 59.15959, 59.19217, 
    59.22448, 59.25651, 59.28826, 59.31973, 59.35091, 59.38182, 59.41245, 
    59.44278, 59.47284, 59.50261, 59.5321, 59.56129, 59.59021, 59.61883, 
    59.64716, 59.6752, 59.70295, 59.73042, 59.75758, 59.78445, 59.81103, 
    59.83731, 59.8633, 59.889, 59.91439, 59.93948, 59.96428, 59.98878, 
    60.01297, 60.03687, 60.06046, 60.08375, 60.10674, 60.12942, 60.1518, 
    60.17387, 60.19564, 60.2171, 60.23825, 60.25909, 60.27963, 60.29985, 
    60.31977, 60.33937, 60.35866, 60.37764, 60.39631, 60.41466, 60.4327, 
    60.45043, 60.46784, 60.48493, 60.50171, 60.51817, 60.53432, 60.55014, 
    60.56565, 60.58084, 60.59571, 60.61026, 60.62449, 60.63839, 60.65198, 
    60.66525, 60.67818, 60.69081, 60.7031, 60.71508, 60.72673, 60.73805, 
    60.74905, 60.75972, 60.77007, 60.7801, 60.78979, 60.79917, 60.80821, 
    60.81693, 60.82532, 60.83338, 60.84111, 60.84852, 60.85559, 60.86235, 
    60.86876, 60.87486, 60.88062, 60.88605, 60.89115, 60.89592, 60.90036, 
    60.90447, 60.90825, 60.9117, 60.91482, 60.91761, 60.92007, 60.9222, 
    60.92399, 60.92545, 60.92659, 60.92739, 60.92786, 60.928, 60.92781, 
    60.92728, 60.92643, 60.92524, 60.92373, 60.92188, 60.9197, 60.91719, 
    60.91435, 60.91118, 60.90768, 60.90384, 60.89968, 60.89519, 60.89036, 
    60.88521, 60.87973, 60.87391, 60.86777, 60.8613, 60.8545, 60.84737, 
    60.83991, 60.83213, 60.82401, 60.81557, 60.8068, 60.79771, 60.78828, 
    60.77853, 60.76846, 60.75806, 60.74733, 60.73628, 60.7249, 60.7132, 
    60.70118, 60.68883, 60.67616, 60.66317, 60.64985, 60.63622, 60.62225, 
    60.60798, 60.59338, 60.57846, 60.56322, 60.54766, 60.53178, 60.51559, 
    60.49908, 60.48225, 60.4651, 60.44764, 60.42987, 60.41178, 60.39338, 
    60.37466, 60.35563, 60.33629, 60.31664, 60.29667, 60.2764, 60.25582, 
    60.23492, 60.21373, 60.19222, 60.1704, 60.14828, 60.12585, 60.10312, 
    60.08009, 60.05675, 60.03311, 60.00917, 59.98492, 59.96038, 59.93554, 
    59.91039, 59.88495, 59.85921, 59.83318, 59.80685, 59.78022, 59.7533, 
    59.72609, 59.69859, 59.67079, 59.6427, 59.61432, 59.58565, 59.55669, 
    59.52745, 59.49792, 59.46811, 59.438, 59.40762, 59.37695, 59.346, 
    59.31477, 59.28325, 59.25146, 59.21939, 59.18704, 59.15441, 59.12151, 
    59.08833, 59.05487, 59.02115, 58.98715, 58.95288, 58.91833, 58.88353, 
    58.84845, 58.8131, 58.77748, 58.7416, 58.70546, 58.66904, 58.63237, 
    58.59544, 58.55824, 58.52078, 58.48306, 58.44509, 58.40686, 58.36837, 
    58.32962, 58.29062, 58.25137, 58.21186, 58.1721, 58.1321, 58.09184, 
    58.05133, 58.01057, 57.96957, 57.92833, 57.88683, 57.8451, 57.80312, 
    57.7609, 57.71843, 57.67573, 57.63279, 57.58961, 57.5462, 57.50254, 
    57.45866, 57.41454, 57.37018, 57.32559, 57.28078, 57.23573, 57.19045, 
    57.14494, 57.09921, 57.05325, 57.00707, 56.96066, 56.91403, 56.86717, 
    56.8201, 56.7728, 56.72528, 56.67755, 56.6296, 56.58143, 56.53305, 
    56.48445, 56.43564,
  51.18799, 51.25282, 51.31751, 51.38207, 51.4465, 51.51078, 51.57494, 
    51.63895, 51.70282, 51.76656, 51.83016, 51.89362, 51.95693, 52.0201, 
    52.08313, 52.14602, 52.20877, 52.27136, 52.33382, 52.39612, 52.45828, 
    52.52029, 52.58215, 52.64386, 52.70543, 52.76683, 52.82809, 52.8892, 
    52.95015, 53.01095, 53.07159, 53.13208, 53.19241, 53.25257, 53.31259, 
    53.37244, 53.43213, 53.49166, 53.55104, 53.61024, 53.66929, 53.72817, 
    53.78688, 53.84543, 53.90381, 53.96202, 54.02007, 54.07795, 54.13565, 
    54.19318, 54.25055, 54.30773, 54.36475, 54.42159, 54.47825, 54.53474, 
    54.59105, 54.64718, 54.70314, 54.75891, 54.8145, 54.86991, 54.92514, 
    54.98018, 55.03504, 55.08971, 55.1442, 55.1985, 55.25261, 55.30654, 
    55.36027, 55.41381, 55.46716, 55.52032, 55.57328, 55.62605, 55.67862, 
    55.731, 55.78317, 55.83515, 55.88693, 55.93851, 55.98989, 56.04107, 
    56.09204, 56.14281, 56.19337, 56.24373, 56.29388, 56.34382, 56.39355, 
    56.44308, 56.49239, 56.54149, 56.59038, 56.63905, 56.68751, 56.73576, 
    56.78378, 56.83159, 56.87918, 56.92655, 56.9737, 57.02063, 57.06733, 
    57.11381, 57.16007, 57.2061, 57.2519, 57.29748, 57.34283, 57.38795, 
    57.43283, 57.47749, 57.52192, 57.56611, 57.61007, 57.65379, 57.69727, 
    57.74052, 57.78352, 57.82629, 57.86882, 57.91111, 57.95315, 57.99495, 
    58.03651, 58.07782, 58.11889, 58.15971, 58.20028, 58.2406, 58.28067, 
    58.32048, 58.36005, 58.39936, 58.43843, 58.47723, 58.51578, 58.55407, 
    58.5921, 58.62988, 58.66739, 58.70464, 58.74163, 58.77836, 58.81483, 
    58.85102, 58.88696, 58.92263, 58.95803, 58.99316, 59.02802, 59.06261, 
    59.09693, 59.13098, 59.16475, 59.19825, 59.23148, 59.26443, 59.2971, 
    59.32949, 59.36161, 59.39345, 59.425, 59.45628, 59.48727, 59.51798, 
    59.5484, 59.57854, 59.6084, 59.63797, 59.66725, 59.69624, 59.72494, 
    59.75335, 59.78148, 59.80931, 59.83685, 59.86409, 59.89104, 59.91769, 
    59.94405, 59.97012, 59.99588, 60.02135, 60.04652, 60.07138, 60.09595, 
    60.12022, 60.14418, 60.16785, 60.1912, 60.21426, 60.23701, 60.25945, 
    60.28159, 60.30342, 60.32494, 60.34615, 60.36706, 60.38765, 60.40794, 
    60.42791, 60.44757, 60.46693, 60.48596, 60.50468, 60.52309, 60.54119, 
    60.55896, 60.57643, 60.59357, 60.6104, 60.62691, 60.6431, 60.65898, 
    60.67453, 60.68977, 60.70468, 60.71928, 60.73355, 60.7475, 60.76113, 
    60.77443, 60.78741, 60.80007, 60.81241, 60.82442, 60.8361, 60.84746, 
    60.85849, 60.8692, 60.87959, 60.88964, 60.89937, 60.90877, 60.91784, 
    60.92658, 60.935, 60.94308, 60.95084, 60.95827, 60.96537, 60.97214, 
    60.97858, 60.98469, 60.99047, 60.99591, 61.00103, 61.00582, 61.01027, 
    61.0144, 61.01819, 61.02165, 61.02478, 61.02758, 61.03004, 61.03218, 
    61.03398, 61.03545, 61.03658, 61.03739, 61.03786, 61.038, 61.03781, 
    61.03728, 61.03643, 61.03524, 61.03371, 61.03186, 61.02967, 61.02716, 
    61.02431, 61.02113, 61.01761, 61.01377, 61.00959, 61.00508, 61.00024, 
    60.99508, 60.98957, 60.98375, 60.97758, 60.97109, 60.96427, 60.95712, 
    60.94964, 60.94183, 60.93369, 60.92522, 60.91642, 60.9073, 60.89785, 
    60.88807, 60.87796, 60.86753, 60.85677, 60.84569, 60.83427, 60.82254, 
    60.81048, 60.79809, 60.78538, 60.77235, 60.75899, 60.74532, 60.73131, 
    60.71699, 60.70235, 60.68738, 60.6721, 60.65649, 60.64056, 60.62432, 
    60.60776, 60.59088, 60.57368, 60.55618, 60.53835, 60.5202, 60.50174, 
    60.48297, 60.46389, 60.44448, 60.42477, 60.40475, 60.38442, 60.36377, 
    60.34282, 60.32156, 60.29998, 60.27811, 60.25592, 60.23343, 60.21063, 
    60.18753, 60.16412, 60.14041, 60.1164, 60.09209, 60.06747, 60.04255, 
    60.01734, 59.99183, 59.96601, 59.9399, 59.9135, 59.8868, 59.8598, 
    59.83251, 59.80492, 59.77705, 59.74888, 59.72042, 59.69167, 59.66264, 
    59.63331, 59.60369, 59.5738, 59.54361, 59.51314, 59.48239, 59.45135, 
    59.42003, 59.38843, 59.35655, 59.32439, 59.29195, 59.25924, 59.22624, 
    59.19297, 59.15943, 59.12561, 59.09152, 59.05716, 59.02253, 58.98762, 
    58.95245, 58.917, 58.88129, 58.84532, 58.80907, 58.77257, 58.7358, 
    58.69877, 58.66147, 58.62392, 58.5861, 58.54803, 58.5097, 58.47111, 
    58.43226, 58.39317, 58.35381, 58.31421, 58.27435, 58.23423, 58.19387, 
    58.15327, 58.11241, 58.0713, 58.02995, 57.98836, 57.94652, 57.90443, 
    57.86211, 57.81955, 57.77674, 57.73369, 57.69041, 57.64688, 57.60313, 
    57.55913, 57.5149, 57.47044, 57.42575, 57.38083, 57.33567, 57.29029, 
    57.24467, 57.19883, 57.15277, 57.10648, 57.05996, 57.01322, 56.96626, 
    56.91907, 56.87167, 56.82404, 56.7762, 56.72814, 56.67986, 56.63137, 
    56.58266, 56.53374,
  51.27598, 51.3409, 51.4057, 51.47036, 51.53489, 51.59928, 51.66354, 
    51.72765, 51.79163, 51.85547, 51.91917, 51.98273, 52.04615, 52.10943, 
    52.17256, 52.23555, 52.2984, 52.36111, 52.42366, 52.48607, 52.54834, 
    52.61045, 52.67242, 52.73424, 52.79591, 52.85742, 52.91879, 52.98, 
    53.04106, 53.10196, 53.16271, 53.2233, 53.28374, 53.34402, 53.40414, 
    53.4641, 53.5239, 53.58354, 53.64302, 53.70234, 53.76149, 53.82048, 
    53.8793, 53.93796, 53.99645, 54.05477, 54.11292, 54.17091, 54.22873, 
    54.28637, 54.34384, 54.40114, 54.45826, 54.51521, 54.57199, 54.62859, 
    54.68501, 54.74125, 54.79731, 54.8532, 54.9089, 54.96442, 55.01976, 
    55.07491, 55.12988, 55.18467, 55.23926, 55.29367, 55.3479, 55.40193, 
    55.45577, 55.50943, 55.56289, 55.61615, 55.66923, 55.72211, 55.77479, 
    55.82727, 55.87957, 55.93166, 55.98355, 56.03524, 56.08673, 56.13801, 
    56.1891, 56.23997, 56.29065, 56.34112, 56.39138, 56.44143, 56.49128, 
    56.54091, 56.59033, 56.63954, 56.68854, 56.73732, 56.78589, 56.83424, 
    56.88238, 56.9303, 56.978, 57.02548, 57.07273, 57.11977, 57.16658, 
    57.21318, 57.25954, 57.30568, 57.35159, 57.39728, 57.44273, 57.48796, 
    57.53296, 57.57772, 57.62225, 57.66655, 57.71061, 57.75444, 57.79803, 
    57.84138, 57.88449, 57.92737, 57.97, 58.01239, 58.05454, 58.09645, 
    58.13811, 58.17952, 58.22069, 58.26161, 58.30228, 58.3427, 58.38288, 
    58.4228, 58.46247, 58.50188, 58.54104, 58.57994, 58.61859, 58.65698, 
    58.69511, 58.73299, 58.7706, 58.80795, 58.84504, 58.88186, 58.91842, 
    58.95472, 58.99075, 59.02651, 59.062, 59.09723, 59.13219, 59.16687, 
    59.20128, 59.23542, 59.26929, 59.30288, 59.3362, 59.36924, 59.402, 
    59.43448, 59.46669, 59.49861, 59.53025, 59.56161, 59.59269, 59.62349, 
    59.654, 59.68422, 59.71416, 59.74381, 59.77317, 59.80225, 59.83103, 
    59.85952, 59.88773, 59.91563, 59.94325, 59.97057, 59.9976, 60.02433, 
    60.05077, 60.0769, 60.10275, 60.12828, 60.15353, 60.17847, 60.20311, 
    60.22744, 60.25148, 60.27521, 60.29864, 60.32176, 60.34457, 60.36708, 
    60.38929, 60.41118, 60.43277, 60.45404, 60.47501, 60.49567, 60.51601, 
    60.53605, 60.55577, 60.57518, 60.59427, 60.61305, 60.63151, 60.64966, 
    60.66749, 60.68501, 60.70221, 60.71909, 60.73565, 60.75189, 60.76781, 
    60.78341, 60.79869, 60.81365, 60.82829, 60.84261, 60.8566, 60.87027, 
    60.88361, 60.89664, 60.90934, 60.92171, 60.93375, 60.94547, 60.95687, 
    60.96794, 60.97868, 60.98909, 60.99918, 61.00893, 61.01836, 61.02747, 
    61.03624, 61.04468, 61.05279, 61.06057, 61.06802, 61.07515, 61.08194, 
    61.08839, 61.09452, 61.10032, 61.10579, 61.11092, 61.11572, 61.12019, 
    61.12432, 61.12813, 61.1316, 61.13474, 61.13755, 61.14002, 61.14216, 
    61.14396, 61.14544, 61.14658, 61.14738, 61.14786, 61.148, 61.1478, 
    61.14728, 61.14642, 61.14523, 61.1437, 61.14184, 61.13965, 61.13712, 
    61.13427, 61.13107, 61.12755, 61.12369, 61.1195, 61.11498, 61.11013, 
    61.10494, 61.09943, 61.09357, 61.08739, 61.08088, 61.07404, 61.06687, 
    61.05936, 61.05153, 61.04337, 61.03487, 61.02605, 61.0169, 61.00741, 
    60.9976, 60.98746, 60.977, 60.96621, 60.95509, 60.94364, 60.93187, 
    60.91977, 60.90735, 60.8946, 60.88153, 60.86813, 60.85441, 60.84036, 
    60.826, 60.81131, 60.7963, 60.78096, 60.76531, 60.74934, 60.73305, 
    60.71643, 60.6995, 60.68226, 60.66469, 60.64681, 60.62861, 60.6101, 
    60.59127, 60.57213, 60.55267, 60.5329, 60.51282, 60.49242, 60.47172, 
    60.4507, 60.42937, 60.40774, 60.3858, 60.36354, 60.34098, 60.31812, 
    60.29495, 60.27148, 60.2477, 60.22361, 60.19923, 60.17454, 60.14956, 
    60.12426, 60.09868, 60.07279, 60.0466, 60.02012, 59.99334, 59.96627, 
    59.9389, 59.91124, 59.88329, 59.85504, 59.8265, 59.79767, 59.76855, 
    59.73914, 59.70944, 59.67946, 59.64919, 59.61864, 59.5878, 59.55667, 
    59.52527, 59.49358, 59.46161, 59.42936, 59.39684, 59.36403, 59.33094, 
    59.29758, 59.26395, 59.23004, 59.19586, 59.1614, 59.12667, 59.09168, 
    59.05641, 59.02087, 58.98507, 58.949, 58.91266, 58.87606, 58.83919, 
    58.80206, 58.76467, 58.72701, 58.6891, 58.65093, 58.6125, 58.57381, 
    58.53486, 58.49566, 58.45621, 58.4165, 58.37654, 58.33633, 58.29587, 
    58.25515, 58.2142, 58.17299, 58.13153, 58.08983, 58.04789, 58.0057, 
    57.96327, 57.9206, 57.87769, 57.83454, 57.79115, 57.74752, 57.70366, 
    57.65956, 57.61522, 57.57065, 57.52585, 57.48082, 57.43556, 57.39006, 
    57.34435, 57.2984, 57.25222, 57.20582, 57.15919, 57.11235, 57.06527, 
    57.01798, 56.97047, 56.92273, 56.87478, 56.82661, 56.77822, 56.72962, 
    56.68081, 56.63177,
  51.36387, 51.4289, 51.4938, 51.55856, 51.62319, 51.68768, 51.75204, 
    51.81626, 51.88034, 51.94429, 52.00809, 52.07175, 52.13528, 52.19866, 
    52.2619, 52.32499, 52.38795, 52.45076, 52.51342, 52.57594, 52.63831, 
    52.70053, 52.7626, 52.82452, 52.8863, 52.94792, 53.00939, 53.07071, 
    53.13188, 53.19289, 53.25374, 53.31445, 53.37499, 53.43538, 53.49561, 
    53.55567, 53.61558, 53.67533, 53.73492, 53.79434, 53.8536, 53.9127, 
    53.97163, 54.0304, 54.089, 54.14743, 54.2057, 54.26379, 54.32172, 
    54.37947, 54.43705, 54.49446, 54.55169, 54.60875, 54.66564, 54.72235, 
    54.77888, 54.83523, 54.89141, 54.9474, 55.00322, 55.05885, 55.1143, 
    55.16956, 55.22464, 55.27954, 55.33425, 55.38877, 55.4431, 55.49725, 
    55.5512, 55.60497, 55.65854, 55.71192, 55.7651, 55.81809, 55.87089, 
    55.92348, 55.97588, 56.02809, 56.08009, 56.13189, 56.18349, 56.23489, 
    56.28608, 56.33707, 56.38786, 56.43844, 56.48881, 56.53897, 56.58893, 
    56.63867, 56.68821, 56.73753, 56.78664, 56.83553, 56.88421, 56.93267, 
    56.98092, 57.02895, 57.07676, 57.12434, 57.17171, 57.21886, 57.26578, 
    57.31248, 57.35895, 57.4052, 57.45122, 57.49701, 57.54258, 57.58791, 
    57.63301, 57.67789, 57.72253, 57.76693, 57.8111, 57.85503, 57.89873, 
    57.94219, 57.98541, 58.02839, 58.07113, 58.11362, 58.15588, 58.19789, 
    58.23965, 58.28117, 58.32244, 58.36347, 58.40424, 58.44477, 58.48504, 
    58.52506, 58.56483, 58.60435, 58.64361, 58.68261, 58.72136, 58.75985, 
    58.79808, 58.83606, 58.87377, 58.91122, 58.9484, 58.98532, 59.02198, 
    59.05837, 59.0945, 59.13036, 59.16595, 59.20127, 59.23632, 59.2711, 
    59.3056, 59.33983, 59.37379, 59.40747, 59.44088, 59.47401, 59.50686, 
    59.53944, 59.57173, 59.60374, 59.63547, 59.66692, 59.69809, 59.72897, 
    59.75956, 59.78987, 59.81989, 59.84963, 59.87907, 59.90823, 59.9371, 
    59.96567, 59.99395, 60.02194, 60.04964, 60.07703, 60.10414, 60.13095, 
    60.15746, 60.18367, 60.20959, 60.2352, 60.26052, 60.28553, 60.31024, 
    60.33465, 60.35876, 60.38256, 60.40605, 60.42924, 60.45213, 60.4747, 
    60.49697, 60.51893, 60.54058, 60.56192, 60.58295, 60.60367, 60.62408, 
    60.64417, 60.66395, 60.68341, 60.70256, 60.7214, 60.73992, 60.75813, 
    60.77601, 60.79358, 60.81083, 60.82776, 60.84437, 60.86066, 60.87663, 
    60.89228, 60.90761, 60.92262, 60.9373, 60.95166, 60.96569, 60.9794, 
    60.99279, 61.00586, 61.01859, 61.031, 61.04309, 61.05484, 61.06627, 
    61.07737, 61.08815, 61.09859, 61.10871, 61.1185, 61.12796, 61.13709, 
    61.14589, 61.15435, 61.16249, 61.1703, 61.17777, 61.18492, 61.19173, 
    61.19821, 61.20435, 61.21017, 61.21565, 61.2208, 61.22562, 61.2301, 
    61.23425, 61.23807, 61.24155, 61.2447, 61.24751, 61.24999, 61.25214, 
    61.25395, 61.25543, 61.25657, 61.25738, 61.25786, 61.258, 61.2578, 
    61.25728, 61.25642, 61.25522, 61.25369, 61.25182, 61.24962, 61.24709, 
    61.24422, 61.24102, 61.23748, 61.23362, 61.22941, 61.22488, 61.22001, 
    61.21481, 61.20927, 61.2034, 61.1972, 61.19067, 61.18381, 61.17661, 
    61.16909, 61.16122, 61.15304, 61.14452, 61.13567, 61.12648, 61.11697, 
    61.10713, 61.09697, 61.08647, 61.07564, 61.06449, 61.05301, 61.04119, 
    61.02906, 61.0166, 61.00381, 60.9907, 60.97726, 60.96349, 60.94941, 
    60.935, 60.92026, 60.9052, 60.88983, 60.87413, 60.8581, 60.84176, 
    60.8251, 60.80812, 60.79082, 60.7732, 60.75526, 60.73701, 60.71844, 
    60.69956, 60.68036, 60.66084, 60.64101, 60.62087, 60.60041, 60.57965, 
    60.55857, 60.53718, 60.51548, 60.49347, 60.47115, 60.44853, 60.42559, 
    60.40236, 60.37881, 60.35496, 60.33081, 60.30635, 60.28159, 60.25653, 
    60.23117, 60.20551, 60.17955, 60.15329, 60.12673, 60.09987, 60.07272, 
    60.04527, 60.01753, 59.9895, 59.96117, 59.93255, 59.90364, 59.87444, 
    59.84494, 59.81516, 59.7851, 59.75474, 59.7241, 59.69318, 59.66196, 
    59.63047, 59.5987, 59.56664, 59.5343, 59.50168, 59.46879, 59.43562, 
    59.40216, 59.36844, 59.33443, 59.30016, 59.26561, 59.23079, 59.1957, 
    59.16034, 59.1247, 59.0888, 59.05264, 59.0162, 58.9795, 58.94254, 
    58.90531, 58.86782, 58.83007, 58.79205, 58.75378, 58.71525, 58.67646, 
    58.63742, 58.59811, 58.55856, 58.51875, 58.47869, 58.43837, 58.39781, 
    58.35699, 58.31593, 58.27462, 58.23306, 58.19126, 58.14921, 58.10692, 
    58.06438, 58.02161, 57.97859, 57.93533, 57.89183, 57.8481, 57.80413, 
    57.75992, 57.71548, 57.67081, 57.6259, 57.58076, 57.53539, 57.48978, 
    57.44396, 57.3979, 57.35162, 57.30511, 57.25837, 57.21141, 57.16423, 
    57.11683, 57.06921, 57.02136, 56.9733, 56.92502, 56.87652, 56.82781, 
    56.77888, 56.72974,
  51.45166, 51.5168, 51.5818, 51.64666, 51.7114, 51.77599, 51.84045, 
    51.90477, 51.96896, 52.033, 52.09691, 52.16068, 52.22431, 52.2878, 
    52.35114, 52.41434, 52.4774, 52.54031, 52.60308, 52.6657, 52.72818, 
    52.79051, 52.85269, 52.91472, 52.9766, 53.03833, 53.09991, 53.16133, 
    53.2226, 53.28372, 53.34469, 53.40549, 53.46615, 53.52664, 53.58698, 
    53.64716, 53.70718, 53.76703, 53.82673, 53.88626, 53.94563, 54.00484, 
    54.06388, 54.12276, 54.18147, 54.24001, 54.29838, 54.35659, 54.41462, 
    54.47248, 54.53018, 54.5877, 54.64504, 54.70221, 54.75921, 54.81603, 
    54.87267, 54.92913, 54.98542, 55.04153, 55.09745, 55.15319, 55.20876, 
    55.26413, 55.31932, 55.37433, 55.42915, 55.48379, 55.53823, 55.59249, 
    55.64655, 55.70043, 55.75411, 55.8076, 55.8609, 55.914, 55.96691, 
    56.01962, 56.07213, 56.12445, 56.17656, 56.22847, 56.28019, 56.3317, 
    56.383, 56.4341, 56.485, 56.53569, 56.58617, 56.63645, 56.68652, 
    56.73637, 56.78601, 56.83545, 56.88467, 56.93367, 56.98246, 57.03103, 
    57.07939, 57.12753, 57.17545, 57.22314, 57.27062, 57.31788, 57.36491, 
    57.41172, 57.4583, 57.50466, 57.55079, 57.59669, 57.64236, 57.68781, 
    57.73302, 57.778, 57.82275, 57.86726, 57.91153, 57.95557, 57.99938, 
    58.04294, 58.08627, 58.12936, 58.1722, 58.2148, 58.25716, 58.29928, 
    58.34114, 58.38277, 58.42414, 58.46527, 58.50615, 58.54678, 58.58716, 
    58.62729, 58.66716, 58.70677, 58.74614, 58.78524, 58.82409, 58.86268, 
    58.90101, 58.93908, 58.97689, 59.01444, 59.05172, 59.08875, 59.1255, 
    59.16199, 59.19821, 59.23417, 59.26985, 59.30526, 59.34041, 59.37528, 
    59.40988, 59.44421, 59.47826, 59.51203, 59.54553, 59.57875, 59.61169, 
    59.64436, 59.67674, 59.70884, 59.74066, 59.7722, 59.80345, 59.83442, 
    59.8651, 59.89549, 59.9256, 59.95542, 59.98495, 60.01419, 60.04313, 
    60.07179, 60.10015, 60.12822, 60.15599, 60.18348, 60.21066, 60.23755, 
    60.26413, 60.29042, 60.31641, 60.3421, 60.36749, 60.39257, 60.41736, 
    60.44184, 60.46601, 60.48989, 60.51345, 60.53671, 60.55966, 60.58231, 
    60.60464, 60.62666, 60.64838, 60.66978, 60.69088, 60.71165, 60.73212, 
    60.75228, 60.77212, 60.79164, 60.81085, 60.82974, 60.84832, 60.86658, 
    60.88452, 60.90214, 60.91944, 60.93642, 60.95309, 60.96943, 60.98545, 
    61.00114, 61.01652, 61.03157, 61.0463, 61.0607, 61.07478, 61.08854, 
    61.10196, 61.11507, 61.12784, 61.14029, 61.15241, 61.16421, 61.17567, 
    61.18681, 61.19762, 61.2081, 61.21824, 61.22806, 61.23755, 61.24671, 
    61.25554, 61.26403, 61.27219, 61.28002, 61.28752, 61.29469, 61.30152, 
    61.30802, 61.31419, 61.32002, 61.32552, 61.33068, 61.33551, 61.34001, 
    61.34417, 61.348, 61.3515, 61.35466, 61.35748, 61.35997, 61.36212, 
    61.36394, 61.36542, 61.36657, 61.36738, 61.36786, 61.368, 61.36781, 
    61.36728, 61.36641, 61.36521, 61.36367, 61.3618, 61.3596, 61.35706, 
    61.35418, 61.35097, 61.34742, 61.34354, 61.33932, 61.33477, 61.32989, 
    61.32467, 61.31912, 61.31323, 61.30701, 61.30046, 61.29358, 61.28636, 
    61.2788, 61.27092, 61.26271, 61.25416, 61.24528, 61.23607, 61.22653, 
    61.21666, 61.20646, 61.19593, 61.18507, 61.17388, 61.16236, 61.15052, 
    61.13834, 61.12584, 61.11301, 61.09986, 61.08638, 61.07257, 61.05844, 
    61.04399, 61.02921, 61.01411, 60.99868, 60.98293, 60.96686, 60.95047, 
    60.93376, 60.91673, 60.89937, 60.8817, 60.86371, 60.8454, 60.82677, 
    60.80783, 60.78857, 60.769, 60.74911, 60.72891, 60.70839, 60.68756, 
    60.66642, 60.64497, 60.6232, 60.60113, 60.57874, 60.55605, 60.53305, 
    60.50974, 60.48613, 60.46221, 60.43799, 60.41346, 60.38863, 60.36349, 
    60.33806, 60.31232, 60.28628, 60.25994, 60.23331, 60.20638, 60.17915, 
    60.15162, 60.1238, 60.09568, 60.06728, 60.03857, 60.00958, 59.98029, 
    59.95072, 59.92086, 59.8907, 59.86026, 59.82954, 59.79852, 59.76723, 
    59.73565, 59.70378, 59.67163, 59.63921, 59.6065, 59.57351, 59.54025, 
    59.50671, 59.47289, 59.43879, 59.40443, 59.36978, 59.33487, 59.29968, 
    59.26422, 59.22849, 59.1925, 59.15623, 59.1197, 59.0829, 59.04584, 
    59.00852, 58.97093, 58.93307, 58.89497, 58.85659, 58.81796, 58.77907, 
    58.73993, 58.70052, 58.66087, 58.62095, 58.58079, 58.54037, 58.4997, 
    58.45879, 58.41762, 58.3762, 58.33454, 58.29263, 58.25048, 58.20808, 
    58.16544, 58.12255, 58.07943, 58.03607, 57.99247, 57.94862, 57.90454, 
    57.86023, 57.81568, 57.7709, 57.72588, 57.68063, 57.63515, 57.58945, 
    57.54351, 57.49734, 57.45095, 57.40433, 57.35749, 57.31042, 57.26313, 
    57.21561, 57.16788, 57.11993, 57.07175, 57.02337, 56.97476, 56.92593, 
    56.87689, 56.82764,
  51.53936, 51.6046, 51.6697, 51.73467, 51.7995, 51.8642, 51.92876, 51.99319, 
    52.05748, 52.12163, 52.18564, 52.24952, 52.31325, 52.37684, 52.44029, 
    52.5036, 52.56676, 52.62978, 52.69265, 52.75538, 52.81796, 52.88039, 
    52.94268, 53.00482, 53.06681, 53.12864, 53.19033, 53.25186, 53.31324, 
    53.37447, 53.43554, 53.49646, 53.55722, 53.61782, 53.67826, 53.73855, 
    53.79868, 53.85865, 53.91845, 53.9781, 54.03757, 54.09689, 54.15604, 
    54.21503, 54.27385, 54.3325, 54.39098, 54.4493, 54.50744, 54.56542, 
    54.62322, 54.68085, 54.73831, 54.79559, 54.8527, 54.90963, 54.96638, 
    55.02296, 55.07935, 55.13557, 55.19161, 55.24746, 55.30313, 55.35862, 
    55.41393, 55.46905, 55.52398, 55.57872, 55.63328, 55.68765, 55.74183, 
    55.79582, 55.84961, 55.90322, 55.95662, 56.00984, 56.06286, 56.11568, 
    56.1683, 56.22073, 56.27296, 56.32498, 56.37681, 56.42843, 56.47985, 
    56.53106, 56.58207, 56.63287, 56.68347, 56.73385, 56.78403, 56.834, 
    56.88375, 56.9333, 56.98263, 57.03174, 57.08065, 57.12933, 57.1778, 
    57.22604, 57.27407, 57.32188, 57.36947, 57.41684, 57.46398, 57.5109, 
    57.55759, 57.60406, 57.6503, 57.69631, 57.74209, 57.78764, 57.83297, 
    57.87805, 57.92291, 57.96753, 58.01191, 58.05606, 58.09997, 58.14364, 
    58.18708, 58.23027, 58.27322, 58.31593, 58.35839, 58.40062, 58.44259, 
    58.48432, 58.5258, 58.56703, 58.60801, 58.64875, 58.68923, 58.72945, 
    58.76943, 58.80915, 58.84861, 58.88782, 58.92677, 58.96546, 59.00389, 
    59.04206, 59.07998, 59.11762, 59.155, 59.19212, 59.22898, 59.26556, 
    59.30188, 59.33793, 59.37371, 59.40923, 59.44446, 59.47943, 59.51412, 
    59.54854, 59.58269, 59.61655, 59.65015, 59.68346, 59.71649, 59.74924, 
    59.78172, 59.81391, 59.84582, 59.87744, 59.90878, 59.93983, 59.9706, 
    60.00108, 60.03128, 60.06118, 60.09079, 60.12011, 60.14914, 60.17788, 
    60.20633, 60.23448, 60.26233, 60.28989, 60.31715, 60.34412, 60.37078, 
    60.39715, 60.42321, 60.44898, 60.47444, 60.4996, 60.52446, 60.54901, 
    60.57326, 60.5972, 60.62083, 60.64416, 60.66718, 60.68989, 60.71229, 
    60.73438, 60.75616, 60.77763, 60.79879, 60.81963, 60.84016, 60.86037, 
    60.88027, 60.89986, 60.91912, 60.93807, 60.95671, 60.97502, 60.99302, 
    61.01069, 61.02805, 61.04508, 61.06179, 61.07818, 61.09425, 61.11, 
    61.12542, 61.14052, 61.15529, 61.16974, 61.18386, 61.19766, 61.21113, 
    61.22427, 61.23709, 61.24958, 61.26174, 61.27357, 61.28507, 61.29624, 
    61.30708, 61.31759, 61.32777, 61.33762, 61.34714, 61.35632, 61.36518, 
    61.3737, 61.38189, 61.38974, 61.39727, 61.40445, 61.41131, 61.41783, 
    61.42402, 61.42987, 61.43538, 61.44057, 61.44541, 61.44992, 61.4541, 
    61.45794, 61.46144, 61.46461, 61.46745, 61.46994, 61.4721, 61.47393, 
    61.47541, 61.47657, 61.47738, 61.47786, 61.478, 61.4778, 61.47727, 
    61.47641, 61.4752, 61.47366, 61.47178, 61.46957, 61.46702, 61.46413, 
    61.46091, 61.45736, 61.45346, 61.44923, 61.44467, 61.43977, 61.43453, 
    61.42896, 61.42306, 61.41682, 61.41025, 61.40334, 61.3961, 61.38852, 
    61.38062, 61.37238, 61.3638, 61.35489, 61.34566, 61.33609, 61.32618, 
    61.31595, 61.30539, 61.29449, 61.28327, 61.27172, 61.25983, 61.24762, 
    61.23508, 61.22222, 61.20902, 61.1955, 61.18165, 61.16748, 61.15298, 
    61.13815, 61.123, 61.10753, 61.09173, 61.07561, 61.05917, 61.04241, 
    61.02532, 61.00792, 60.99019, 60.97215, 60.95378, 60.9351, 60.9161, 
    60.89678, 60.87714, 60.8572, 60.83693, 60.81635, 60.79546, 60.77426, 
    60.75274, 60.73091, 60.70877, 60.68632, 60.66356, 60.64049, 60.61712, 
    60.59343, 60.56944, 60.54515, 60.52055, 60.49564, 60.47043, 60.44492, 
    60.41911, 60.393, 60.36658, 60.33987, 60.31286, 60.28555, 60.25795, 
    60.23005, 60.20185, 60.17336, 60.14457, 60.11549, 60.08613, 60.05647, 
    60.02652, 59.99628, 59.96576, 59.93494, 59.90384, 59.87246, 59.84079, 
    59.80883, 59.7766, 59.74408, 59.71128, 59.67821, 59.64485, 59.61122, 
    59.5773, 59.54312, 59.50866, 59.47392, 59.43891, 59.40363, 59.36807, 
    59.33225, 59.29615, 59.25979, 59.22316, 59.18627, 59.14911, 59.11168, 
    59.07399, 59.03605, 58.99783, 58.95936, 58.92063, 58.88163, 58.84239, 
    58.80288, 58.76312, 58.72311, 58.68284, 58.64232, 58.60155, 58.56052, 
    58.51925, 58.47773, 58.43597, 58.39395, 58.35169, 58.30919, 58.26644, 
    58.22345, 58.18022, 58.13675, 58.09304, 58.04909, 58.00491, 57.96048, 
    57.91583, 57.87094, 57.82581, 57.78046, 57.73487, 57.68905, 57.643, 
    57.59673, 57.55022, 57.50349, 57.45654, 57.40936, 57.36196, 57.31434, 
    57.26649, 57.21843, 57.17014, 57.12164, 57.07293, 57.02399, 56.97484, 
    56.92548,
  51.62696, 51.6923, 51.75751, 51.82258, 51.88752, 51.95232, 52.01698, 
    52.08151, 52.14591, 52.21016, 52.27428, 52.33826, 52.40209, 52.46579, 
    52.52934, 52.59275, 52.65602, 52.71915, 52.78213, 52.84496, 52.90765, 
    52.97019, 53.03259, 53.09483, 53.15692, 53.21887, 53.28066, 53.3423, 
    53.40379, 53.46512, 53.5263, 53.58733, 53.6482, 53.70891, 53.76946, 
    53.82986, 53.89009, 53.95017, 54.01009, 54.06984, 54.12943, 54.18885, 
    54.24812, 54.30721, 54.36614, 54.4249, 54.4835, 54.54192, 54.60018, 
    54.65827, 54.71618, 54.77392, 54.83149, 54.88888, 54.9461, 55.00314, 
    55.06001, 55.1167, 55.17321, 55.22953, 55.28568, 55.34165, 55.39743, 
    55.45303, 55.50845, 55.56368, 55.61873, 55.67358, 55.72826, 55.78274, 
    55.83703, 55.89113, 55.94503, 55.99875, 56.05227, 56.1056, 56.15873, 
    56.21167, 56.2644, 56.31694, 56.36928, 56.42142, 56.47335, 56.52509, 
    56.57662, 56.62795, 56.67907, 56.72998, 56.78069, 56.83119, 56.88148, 
    56.93156, 56.98143, 57.03108, 57.08052, 57.12975, 57.17876, 57.22756, 
    57.27614, 57.3245, 57.37264, 57.42056, 57.46826, 57.51574, 57.56299, 
    57.61002, 57.65682, 57.7034, 57.74975, 57.79587, 57.84176, 57.88742, 
    57.93285, 57.97805, 58.02301, 58.06774, 58.11223, 58.15649, 58.20051, 
    58.24429, 58.28783, 58.33113, 58.37419, 58.417, 58.45958, 58.5019, 
    58.54398, 58.58582, 58.6274, 58.66874, 58.70983, 58.75066, 58.79125, 
    58.83158, 58.87165, 58.91148, 58.95105, 58.99036, 59.02941, 59.0682, 
    59.10673, 59.145, 59.18301, 59.22076, 59.25824, 59.29546, 59.33241, 
    59.36909, 59.40551, 59.44166, 59.47754, 59.51315, 59.54848, 59.58354, 
    59.61833, 59.65284, 59.68708, 59.72104, 59.75473, 59.78813, 59.82125, 
    59.8541, 59.88667, 59.91895, 59.95094, 59.98265, 60.01408, 60.04523, 
    60.07608, 60.10665, 60.13692, 60.16691, 60.19661, 60.22602, 60.25513, 
    60.28395, 60.31248, 60.34071, 60.36864, 60.39628, 60.42362, 60.45066, 
    60.47741, 60.50385, 60.52999, 60.55583, 60.58137, 60.60661, 60.63153, 
    60.65616, 60.68048, 60.70449, 60.7282, 60.75159, 60.77468, 60.79746, 
    60.81993, 60.84209, 60.86393, 60.88546, 60.90668, 60.92759, 60.94818, 
    60.96846, 60.98841, 61.00806, 61.02739, 61.04639, 61.06508, 61.08345, 
    61.1015, 61.11923, 61.13664, 61.15372, 61.17049, 61.18693, 61.20305, 
    61.21885, 61.23431, 61.24946, 61.26428, 61.27877, 61.29294, 61.30678, 
    61.32029, 61.33347, 61.34633, 61.35886, 61.37106, 61.38292, 61.39446, 
    61.40567, 61.41654, 61.42709, 61.4373, 61.44718, 61.45673, 61.46594, 
    61.47482, 61.48337, 61.49158, 61.49947, 61.50701, 61.51422, 61.5211, 
    61.52764, 61.53384, 61.53971, 61.54525, 61.55045, 61.55531, 61.55983, 
    61.56403, 61.56787, 61.57139, 61.57457, 61.57741, 61.57992, 61.58208, 
    61.58391, 61.5854, 61.58656, 61.58738, 61.58786, 61.588, 61.5878, 
    61.58727, 61.5864, 61.58519, 61.58364, 61.58176, 61.57954, 61.57698, 
    61.57409, 61.57086, 61.56729, 61.56339, 61.55914, 61.55456, 61.54965, 
    61.5444, 61.53881, 61.53289, 61.52663, 61.52003, 61.5131, 61.50584, 
    61.49824, 61.49031, 61.48204, 61.47344, 61.4645, 61.45524, 61.44564, 
    61.4357, 61.42544, 61.41484, 61.40392, 61.39265, 61.38107, 61.36915, 
    61.3569, 61.34432, 61.33141, 61.31818, 61.30461, 61.29072, 61.2765, 
    61.26196, 61.24709, 61.23189, 61.21637, 61.20052, 61.18435, 61.16786, 
    61.15104, 61.13391, 61.11645, 61.09867, 61.08057, 61.06215, 61.04341, 
    61.02435, 61.00497, 60.98528, 60.96527, 60.94494, 60.9243, 60.90335, 
    60.88208, 60.8605, 60.8386, 60.81639, 60.79388, 60.77105, 60.74791, 
    60.72447, 60.70071, 60.67665, 60.65228, 60.62761, 60.60263, 60.57735, 
    60.55177, 60.52588, 60.49969, 60.4732, 60.44641, 60.41932, 60.39193, 
    60.36424, 60.33626, 60.30798, 60.27941, 60.25055, 60.22139, 60.19193, 
    60.16219, 60.13216, 60.10183, 60.07122, 60.04032, 60.00913, 59.97766, 
    59.9459, 59.91386, 59.88153, 59.84892, 59.81604, 59.78287, 59.74942, 
    59.71569, 59.68169, 59.6474, 59.61285, 59.57801, 59.54291, 59.50753, 
    59.47188, 59.43596, 59.39977, 59.36331, 59.32658, 59.28959, 59.25233, 
    59.21481, 59.17702, 59.13897, 59.10065, 59.06208, 59.02325, 58.98415, 
    58.94481, 58.9052, 58.86533, 58.82521, 58.78484, 58.74422, 58.70334, 
    58.66222, 58.62084, 58.57922, 58.53734, 58.49522, 58.45286, 58.41025, 
    58.36739, 58.3243, 58.28096, 58.23738, 58.19356, 58.14951, 58.10521, 
    58.06068, 58.01591, 57.97091, 57.92568, 57.88021, 57.83452, 57.78859, 
    57.74243, 57.69604, 57.64943, 57.60259, 57.55553, 57.50824, 57.46073, 
    57.41299, 57.36504, 57.31686, 57.26847, 57.21986, 57.17102, 57.12198, 
    57.07272, 57.02324,
  51.71447, 51.77991, 51.84522, 51.91039, 51.97543, 52.04034, 52.10511, 
    52.16974, 52.23424, 52.2986, 52.36282, 52.4269, 52.49084, 52.55464, 
    52.6183, 52.68182, 52.74519, 52.80843, 52.87151, 52.93445, 52.99725, 
    53.05989, 53.12239, 53.18475, 53.24694, 53.309, 53.3709, 53.43265, 
    53.49424, 53.55569, 53.61697, 53.67811, 53.73909, 53.79991, 53.86057, 
    53.92107, 53.98142, 54.04161, 54.10163, 54.1615, 54.2212, 54.28073, 
    54.3401, 54.39931, 54.45835, 54.51722, 54.57593, 54.63446, 54.69283, 
    54.75103, 54.80905, 54.86691, 54.92458, 54.98209, 55.03942, 55.09658, 
    55.15355, 55.21035, 55.26697, 55.32341, 55.37967, 55.43575, 55.49165, 
    55.54736, 55.60289, 55.65824, 55.71339, 55.76837, 55.82315, 55.87774, 
    55.93215, 55.98636, 56.04038, 56.09421, 56.14784, 56.20128, 56.25453, 
    56.30758, 56.36042, 56.41308, 56.46553, 56.51778, 56.56983, 56.62168, 
    56.67332, 56.72476, 56.77599, 56.82702, 56.87784, 56.92846, 56.97886, 
    57.02905, 57.07903, 57.1288, 57.17835, 57.22769, 57.27681, 57.32572, 
    57.37441, 57.42289, 57.47114, 57.51917, 57.56698, 57.61457, 57.66193, 
    57.70907, 57.75599, 57.80268, 57.84914, 57.89537, 57.94137, 57.98714, 
    58.03268, 58.07798, 58.12306, 58.1679, 58.2125, 58.25686, 58.30099, 
    58.34488, 58.38853, 58.43193, 58.4751, 58.51802, 58.5607, 58.60313, 
    58.64532, 58.68726, 58.72895, 58.7704, 58.81159, 58.85253, 58.89322, 
    58.93365, 58.97383, 59.01376, 59.05343, 59.09284, 59.132, 59.17089, 
    59.20953, 59.2479, 59.28601, 59.32386, 59.36144, 59.39875, 59.43581, 
    59.47259, 59.50911, 59.54535, 59.58133, 59.61703, 59.65246, 59.68762, 
    59.7225, 59.75711, 59.79144, 59.8255, 59.85927, 59.89277, 59.92599, 
    59.95892, 59.99158, 60.02395, 60.05604, 60.08784, 60.11935, 60.15059, 
    60.18153, 60.21218, 60.24255, 60.27262, 60.3024, 60.33189, 60.36109, 
    60.38999, 60.4186, 60.44691, 60.47493, 60.50265, 60.53007, 60.55719, 
    60.58401, 60.61053, 60.63675, 60.66267, 60.68828, 60.71359, 60.73859, 
    60.76329, 60.78768, 60.81177, 60.83554, 60.85901, 60.88217, 60.90501, 
    60.92755, 60.94977, 60.97168, 60.99328, 61.01456, 61.03553, 61.05619, 
    61.07653, 61.09655, 61.11625, 61.13563, 61.1547, 61.17345, 61.19187, 
    61.20998, 61.22776, 61.24522, 61.26236, 61.27918, 61.29567, 61.31184, 
    61.32768, 61.3432, 61.35839, 61.37326, 61.3878, 61.40201, 61.41589, 
    61.42944, 61.44267, 61.45557, 61.46813, 61.48037, 61.49227, 61.50385, 
    61.51509, 61.526, 61.53658, 61.54682, 61.55673, 61.56631, 61.57555, 
    61.58446, 61.59304, 61.60128, 61.60918, 61.61675, 61.62399, 61.63089, 
    61.63745, 61.64367, 61.64956, 61.65511, 61.66033, 61.6652, 61.66975, 
    61.67395, 61.67781, 61.68134, 61.68453, 61.68738, 61.68989, 61.69207, 
    61.6939, 61.6954, 61.69656, 61.69738, 61.69786, 61.698, 61.6978, 
    61.69727, 61.6964, 61.69518, 61.69363, 61.69174, 61.68951, 61.68695, 
    61.68405, 61.68081, 61.67722, 61.67331, 61.66905, 61.66446, 61.65953, 
    61.65426, 61.64865, 61.64271, 61.63643, 61.62981, 61.62286, 61.61558, 
    61.60796, 61.59999, 61.5917, 61.58308, 61.57411, 61.56482, 61.55518, 
    61.54522, 61.53492, 61.52429, 61.51333, 61.50204, 61.49041, 61.47845, 
    61.46617, 61.45355, 61.4406, 61.42732, 61.41372, 61.39978, 61.38552, 
    61.37093, 61.35601, 61.34077, 61.3252, 61.3093, 61.29308, 61.27654, 
    61.25967, 61.24248, 61.22497, 61.20713, 61.18898, 61.1705, 61.1517, 
    61.13259, 61.11315, 61.0934, 61.07333, 61.05294, 61.03224, 61.01122, 
    60.98989, 60.96824, 60.94628, 60.924, 60.90142, 60.87852, 60.85532, 
    60.8318, 60.80798, 60.78384, 60.7594, 60.73466, 60.70961, 60.68425, 
    60.65859, 60.63263, 60.60636, 60.57979, 60.55292, 60.52575, 60.49828, 
    60.47052, 60.44246, 60.4141, 60.38544, 60.35649, 60.32725, 60.29771, 
    60.26788, 60.23776, 60.20735, 60.17665, 60.14566, 60.11439, 60.08283, 
    60.05098, 60.01885, 59.98643, 59.95373, 59.92075, 59.88749, 59.85395, 
    59.82013, 59.78603, 59.75165, 59.717, 59.68208, 59.64687, 59.6114, 
    59.57565, 59.53963, 59.50335, 59.46679, 59.42996, 59.39287, 59.35551, 
    59.31789, 59.28, 59.24185, 59.20343, 59.16476, 59.12582, 59.08662, 
    59.04717, 59.00746, 58.96749, 58.92727, 58.8868, 58.84607, 58.80509, 
    58.76386, 58.72237, 58.68064, 58.63866, 58.59644, 58.55397, 58.51125, 
    58.46829, 58.42508, 58.38164, 58.33795, 58.29403, 58.24986, 58.20546, 
    58.16082, 58.11594, 58.07084, 58.02549, 57.97992, 57.93411, 57.88807, 
    57.8418, 57.79531, 57.74858, 57.70163, 57.65446, 57.60706, 57.55943, 
    57.51159, 57.46352, 57.41523, 57.36673, 57.318, 57.26906, 57.2199, 
    57.17052, 57.12094,
  51.80188, 51.86742, 51.93283, 51.9981, 52.06325, 52.12826, 52.19313, 
    52.25787, 52.32247, 52.38693, 52.45126, 52.51545, 52.57949, 52.6434, 
    52.70716, 52.77079, 52.83427, 52.89761, 52.9608, 53.02385, 53.08675, 
    53.1495, 53.21211, 53.27457, 53.33688, 53.39904, 53.46104, 53.5229, 
    53.58461, 53.64616, 53.70755, 53.7688, 53.82988, 53.89082, 53.95159, 
    54.0122, 54.07265, 54.13295, 54.19308, 54.25306, 54.31287, 54.37252, 
    54.432, 54.49132, 54.55047, 54.60945, 54.66827, 54.72692, 54.7854, 
    54.8437, 54.90184, 54.9598, 55.0176, 55.07521, 55.13266, 55.18992, 
    55.24701, 55.30392, 55.36066, 55.41721, 55.47358, 55.52978, 55.58578, 
    55.64161, 55.69725, 55.75271, 55.80798, 55.86307, 55.91796, 55.97267, 
    56.02719, 56.08151, 56.13565, 56.18959, 56.24334, 56.29689, 56.35025, 
    56.40341, 56.45638, 56.50914, 56.5617, 56.61407, 56.66623, 56.71819, 
    56.76995, 56.8215, 56.87285, 56.92399, 56.97492, 57.02565, 57.07616, 
    57.12647, 57.17656, 57.22644, 57.27611, 57.32556, 57.3748, 57.42382, 
    57.47262, 57.52121, 57.56957, 57.61771, 57.66564, 57.71334, 57.76081, 
    57.80806, 57.85509, 57.90189, 57.94846, 57.9948, 58.04092, 58.0868, 
    58.13245, 58.17786, 58.22305, 58.26799, 58.31271, 58.35718, 58.40142, 
    58.44541, 58.48917, 58.53268, 58.57596, 58.61899, 58.66177, 58.70432, 
    58.74661, 58.78865, 58.83045, 58.872, 58.9133, 58.95435, 58.99514, 
    59.03568, 59.07597, 59.116, 59.15577, 59.19529, 59.23454, 59.27354, 
    59.31227, 59.35075, 59.38896, 59.42691, 59.46459, 59.50201, 59.53916, 
    59.57604, 59.61266, 59.649, 59.68507, 59.72087, 59.7564, 59.79165, 
    59.82663, 59.86134, 59.89576, 59.92991, 59.96378, 59.99738, 60.03069, 
    60.06371, 60.09646, 60.12892, 60.1611, 60.19299, 60.22459, 60.25591, 
    60.28695, 60.31768, 60.34814, 60.3783, 60.40816, 60.43774, 60.46702, 
    60.49601, 60.5247, 60.5531, 60.58119, 60.60899, 60.63649, 60.66369, 
    60.69059, 60.71719, 60.74349, 60.76948, 60.79517, 60.82055, 60.84563, 
    60.8704, 60.89487, 60.91902, 60.94287, 60.96641, 60.98963, 61.01255, 
    61.03515, 61.05745, 61.07942, 61.10109, 61.12243, 61.14347, 61.16418, 
    61.18458, 61.20466, 61.22443, 61.24387, 61.26299, 61.2818, 61.30028, 
    61.31844, 61.33628, 61.3538, 61.37099, 61.38786, 61.4044, 61.42062, 
    61.43651, 61.45208, 61.46732, 61.48223, 61.49681, 61.51107, 61.525, 
    61.53859, 61.55186, 61.5648, 61.5774, 61.58968, 61.60162, 61.61323, 
    61.6245, 61.63545, 61.64606, 61.65634, 61.66628, 61.67589, 61.68516, 
    61.6941, 61.7027, 61.71097, 61.7189, 61.72649, 61.73375, 61.74067, 
    61.74725, 61.7535, 61.75941, 61.76498, 61.77021, 61.7751, 61.77966, 
    61.78387, 61.78775, 61.79129, 61.79448, 61.79734, 61.79987, 61.80204, 
    61.80389, 61.80539, 61.80655, 61.80737, 61.80786, 61.808, 61.8078, 
    61.80727, 61.80639, 61.80517, 61.80362, 61.80172, 61.79949, 61.79691, 
    61.794, 61.79075, 61.78716, 61.78323, 61.77896, 61.77435, 61.7694, 
    61.76412, 61.7585, 61.75253, 61.74623, 61.7396, 61.73262, 61.72532, 
    61.71767, 61.70968, 61.70136, 61.69271, 61.68372, 61.67439, 61.66473, 
    61.65474, 61.64441, 61.63374, 61.62274, 61.61141, 61.59975, 61.58776, 
    61.57543, 61.56277, 61.54978, 61.53646, 61.52282, 61.50884, 61.49453, 
    61.47989, 61.46493, 61.44964, 61.43402, 61.41808, 61.40181, 61.38521, 
    61.36829, 61.35105, 61.33348, 61.31559, 61.29738, 61.27885, 61.25999, 
    61.24081, 61.22132, 61.20151, 61.18138, 61.16093, 61.14016, 61.11908, 
    61.09768, 61.07597, 61.05394, 61.0316, 61.00895, 60.98598, 60.9627, 
    60.93912, 60.91522, 60.89102, 60.8665, 60.84168, 60.81656, 60.79113, 
    60.76539, 60.73935, 60.71301, 60.68636, 60.65941, 60.63216, 60.60461, 
    60.57677, 60.54862, 60.52018, 60.49144, 60.46241, 60.43308, 60.40346, 
    60.37355, 60.34334, 60.31284, 60.28205, 60.25098, 60.21962, 60.18797, 
    60.15602, 60.1238, 60.0913, 60.05851, 60.02543, 59.99208, 59.95844, 
    59.92453, 59.89034, 59.85587, 59.82112, 59.78609, 59.7508, 59.71523, 
    59.67938, 59.64327, 59.60688, 59.57022, 59.5333, 59.49611, 59.45865, 
    59.42093, 59.38293, 59.34468, 59.30616, 59.26739, 59.22835, 59.18905, 
    59.14949, 59.10968, 59.06961, 59.02929, 58.9887, 58.94787, 58.90678, 
    58.86545, 58.82386, 58.78202, 58.73993, 58.6976, 58.65502, 58.6122, 
    58.56913, 58.52582, 58.48227, 58.43847, 58.39443, 58.35016, 58.30565, 
    58.2609, 58.21592, 58.1707, 58.12524, 58.07956, 58.03364, 57.98749, 
    57.94111, 57.8945, 57.84767, 57.80061, 57.75332, 57.70581, 57.65807, 
    57.61012, 57.56194, 57.51353, 57.46492, 57.41608, 57.36702, 57.31775, 
    57.26827, 57.21857,
  51.88918, 51.95483, 52.02034, 52.08572, 52.15097, 52.21608, 52.28106, 
    52.3459, 52.41061, 52.47517, 52.5396, 52.6039, 52.66805, 52.73206, 
    52.79593, 52.85966, 52.92325, 52.98669, 53.04999, 53.11314, 53.17615, 
    53.23901, 53.30173, 53.3643, 53.42671, 53.48898, 53.55109, 53.61306, 
    53.67487, 53.73653, 53.79804, 53.85939, 53.92059, 53.98163, 54.04251, 
    54.10323, 54.1638, 54.22421, 54.28445, 54.34454, 54.40445, 54.46421, 
    54.52381, 54.58324, 54.6425, 54.7016, 54.76052, 54.81928, 54.87787, 
    54.93629, 54.99454, 55.05262, 55.11052, 55.16825, 55.2258, 55.28318, 
    55.34039, 55.39741, 55.45426, 55.51093, 55.56741, 55.62371, 55.67984, 
    55.73578, 55.79153, 55.8471, 55.90249, 55.95769, 56.0127, 56.06752, 
    56.12215, 56.17659, 56.23083, 56.28489, 56.33875, 56.39242, 56.44589, 
    56.49917, 56.55225, 56.60512, 56.6578, 56.71028, 56.76256, 56.81463, 
    56.8665, 56.91817, 56.96963, 57.02089, 57.07193, 57.12277, 57.1734, 
    57.22382, 57.27402, 57.32402, 57.3738, 57.42336, 57.47271, 57.52185, 
    57.57076, 57.61946, 57.66794, 57.71619, 57.76423, 57.81204, 57.85963, 
    57.90699, 57.95413, 58.00104, 58.04772, 58.09418, 58.1404, 58.18639, 
    58.23215, 58.27768, 58.32298, 58.36803, 58.41285, 58.45744, 58.50178, 
    58.54589, 58.58976, 58.63338, 58.67676, 58.7199, 58.76279, 58.80544, 
    58.84784, 58.89, 58.9319, 58.97356, 59.01496, 59.05611, 59.09701, 
    59.13766, 59.17805, 59.21818, 59.25806, 59.29768, 59.33704, 59.37614, 
    59.41498, 59.45356, 59.49187, 59.52992, 59.5677, 59.60522, 59.64247, 
    59.67945, 59.71616, 59.75261, 59.78878, 59.82468, 59.8603, 59.89565, 
    59.93073, 59.96553, 60.00005, 60.03429, 60.06826, 60.10194, 60.13535, 
    60.16847, 60.20131, 60.23386, 60.26613, 60.29811, 60.3298, 60.36121, 
    60.39233, 60.42316, 60.4537, 60.48394, 60.5139, 60.54356, 60.57293, 
    60.602, 60.63077, 60.65925, 60.68743, 60.71531, 60.74289, 60.77017, 
    60.79715, 60.82383, 60.8502, 60.87627, 60.90204, 60.9275, 60.95265, 
    60.97749, 61.00203, 61.02626, 61.05018, 61.07379, 61.09708, 61.12007, 
    61.14274, 61.1651, 61.18714, 61.20887, 61.23029, 61.25138, 61.27216, 
    61.29263, 61.31277, 61.33259, 61.3521, 61.37128, 61.39014, 61.40868, 
    61.4269, 61.44479, 61.46236, 61.47961, 61.49653, 61.51312, 61.52939, 
    61.54533, 61.56095, 61.57624, 61.5912, 61.60583, 61.62012, 61.63409, 
    61.64774, 61.66105, 61.67402, 61.68666, 61.69898, 61.71096, 61.72261, 
    61.73392, 61.7449, 61.75554, 61.76585, 61.77583, 61.78547, 61.79477, 
    61.80373, 61.81236, 61.82066, 61.82861, 61.83623, 61.84351, 61.85045, 
    61.85706, 61.86332, 61.86925, 61.87484, 61.88008, 61.88499, 61.88956, 
    61.89379, 61.89768, 61.90123, 61.90444, 61.90731, 61.90984, 61.91203, 
    61.91387, 61.91538, 61.91655, 61.91737, 61.91785, 61.918, 61.9178, 
    61.91726, 61.91639, 61.91516, 61.9136, 61.9117, 61.90946, 61.90688, 
    61.90396, 61.90069, 61.89709, 61.89315, 61.88886, 61.88424, 61.87928, 
    61.87398, 61.86834, 61.86235, 61.85604, 61.84938, 61.84238, 61.83505, 
    61.82738, 61.81937, 61.81102, 61.80234, 61.79332, 61.78396, 61.77427, 
    61.76424, 61.75388, 61.74318, 61.73215, 61.72079, 61.70909, 61.69705, 
    61.68469, 61.67199, 61.65896, 61.6456, 61.63191, 61.61789, 61.60353, 
    61.58885, 61.57384, 61.5585, 61.54284, 61.52684, 61.51052, 61.49387, 
    61.4769, 61.45961, 61.44198, 61.42404, 61.40577, 61.38718, 61.36826, 
    61.34903, 61.32948, 61.3096, 61.28941, 61.2689, 61.24807, 61.22692, 
    61.20546, 61.18368, 61.16158, 61.13918, 61.11646, 61.09342, 61.07007, 
    61.04642, 61.02245, 60.99817, 60.97358, 60.94869, 60.92349, 60.89798, 
    60.87217, 60.84605, 60.81963, 60.7929, 60.76588, 60.73855, 60.71092, 
    60.68299, 60.65477, 60.62624, 60.59742, 60.5683, 60.53889, 60.50918, 
    60.47918, 60.44889, 60.4183, 60.38743, 60.35626, 60.32481, 60.29307, 
    60.26104, 60.22873, 60.19613, 60.16325, 60.13008, 60.09663, 60.0629, 
    60.0289, 59.99461, 59.96004, 59.9252, 59.89008, 59.85468, 59.81902, 
    59.78307, 59.74686, 59.71038, 59.67362, 59.6366, 59.5993, 59.56174, 
    59.52392, 59.48582, 59.44747, 59.40885, 59.36997, 59.33083, 59.29143, 
    59.25177, 59.21185, 59.17168, 59.13124, 59.09056, 59.04962, 59.00843, 
    58.96698, 58.92529, 58.88335, 58.84115, 58.79871, 58.75602, 58.71309, 
    58.66991, 58.6265, 58.58283, 58.53893, 58.49479, 58.4504, 58.40578, 
    58.36092, 58.31583, 58.2705, 58.22493, 58.17913, 58.13311, 58.08685, 
    58.04036, 57.99364, 57.94669, 57.89952, 57.85212, 57.80449, 57.75665, 
    57.70858, 57.66029, 57.61177, 57.56304, 57.51409, 57.46492, 57.41554, 
    57.36594, 57.31612,
  51.97639, 52.04214, 52.10775, 52.17324, 52.23859, 52.30381, 52.36889, 
    52.43383, 52.49864, 52.56332, 52.62785, 52.69225, 52.75651, 52.82063, 
    52.8846, 52.94844, 53.01213, 53.07568, 53.13908, 53.20235, 53.26546, 
    53.32843, 53.39125, 53.45393, 53.51645, 53.57883, 53.64105, 53.70313, 
    53.76505, 53.82682, 53.88844, 53.94989, 54.0112, 54.07235, 54.13334, 
    54.19418, 54.25485, 54.31537, 54.37572, 54.43592, 54.49595, 54.55582, 
    54.61552, 54.67506, 54.73444, 54.79364, 54.85268, 54.91156, 54.97026, 
    55.02879, 55.08715, 55.14534, 55.20336, 55.2612, 55.31887, 55.37636, 
    55.43367, 55.49081, 55.54777, 55.60455, 55.66115, 55.71757, 55.77381, 
    55.82986, 55.88573, 55.94141, 55.99691, 56.05222, 56.10735, 56.16228, 
    56.21703, 56.27158, 56.32594, 56.38012, 56.43409, 56.48787, 56.54146, 
    56.59485, 56.64804, 56.70103, 56.75383, 56.80642, 56.85881, 56.911, 
    56.96298, 57.01476, 57.06634, 57.11771, 57.16887, 57.21982, 57.27057, 
    57.32109, 57.37141, 57.42152, 57.47142, 57.5211, 57.57056, 57.61981, 
    57.66884, 57.71765, 57.76624, 57.81461, 57.86275, 57.91068, 57.95838, 
    58.00586, 58.05311, 58.10013, 58.14692, 58.19349, 58.23982, 58.28593, 
    58.3318, 58.37744, 58.42284, 58.46801, 58.51294, 58.55764, 58.60209, 
    58.64631, 58.69028, 58.73402, 58.77751, 58.82076, 58.86376, 58.90651, 
    58.94902, 58.99128, 59.03329, 59.07506, 59.11657, 59.15783, 59.19883, 
    59.23959, 59.28008, 59.32032, 59.3603, 59.40002, 59.43949, 59.47869, 
    59.51764, 59.55632, 59.59473, 59.63288, 59.67077, 59.70839, 59.74574, 
    59.78282, 59.81963, 59.85617, 59.89244, 59.92844, 59.96416, 59.99961, 
    60.03479, 60.06968, 60.1043, 60.13864, 60.1727, 60.20648, 60.23997, 
    60.27319, 60.30612, 60.33876, 60.37112, 60.4032, 60.43498, 60.46648, 
    60.49769, 60.52861, 60.55923, 60.58957, 60.61961, 60.64935, 60.6788, 
    60.70796, 60.73682, 60.76538, 60.79364, 60.82161, 60.84927, 60.87663, 
    60.90369, 60.93044, 60.95689, 60.98304, 61.00888, 61.03442, 61.05965, 
    61.08457, 61.10918, 61.13348, 61.15747, 61.18115, 61.20452, 61.22757, 
    61.25031, 61.27274, 61.29485, 61.31664, 61.33812, 61.35928, 61.38013, 
    61.40065, 61.42086, 61.44074, 61.46031, 61.47955, 61.49847, 61.51707, 
    61.53534, 61.55329, 61.57092, 61.58821, 61.60519, 61.62184, 61.63816, 
    61.65415, 61.66982, 61.68515, 61.70015, 61.71483, 61.72918, 61.74319, 
    61.75687, 61.77022, 61.78324, 61.79593, 61.80828, 61.8203, 61.83198, 
    61.84333, 61.85434, 61.86502, 61.87536, 61.88537, 61.89504, 61.90437, 
    61.91337, 61.92202, 61.93034, 61.93832, 61.94597, 61.95327, 61.96024, 
    61.96686, 61.97315, 61.97909, 61.9847, 61.98996, 61.99489, 61.99947, 
    62.00372, 62.00762, 62.01118, 62.0144, 62.01728, 62.01981, 62.02201, 
    62.02386, 62.02537, 62.02654, 62.02737, 62.02785, 62.028, 62.0278, 
    62.02726, 62.02638, 62.02515, 62.02359, 62.02168, 62.01943, 62.01684, 
    62.01391, 62.01064, 62.00702, 62.00307, 61.99877, 61.99413, 61.98915, 
    61.98383, 61.97818, 61.97218, 61.96584, 61.95916, 61.95214, 61.94478, 
    61.93708, 61.92905, 61.92068, 61.91197, 61.90292, 61.89353, 61.88381, 
    61.87375, 61.86335, 61.85262, 61.84156, 61.83015, 61.81842, 61.80635, 
    61.79394, 61.7812, 61.76813, 61.75473, 61.74099, 61.72693, 61.71253, 
    61.6978, 61.68274, 61.66736, 61.65164, 61.6356, 61.61922, 61.60253, 
    61.5855, 61.56815, 61.55047, 61.53247, 61.51415, 61.4955, 61.47653, 
    61.45723, 61.43762, 61.41768, 61.39743, 61.37685, 61.35596, 61.33475, 
    61.31322, 61.29137, 61.26921, 61.24673, 61.22395, 61.20084, 61.17743, 
    61.15369, 61.12965, 61.1053, 61.08065, 61.05568, 61.0304, 61.00481, 
    60.97893, 60.95273, 60.92623, 60.89943, 60.87232, 60.84491, 60.8172, 
    60.78919, 60.76088, 60.73227, 60.70337, 60.67416, 60.64467, 60.61488, 
    60.58479, 60.55441, 60.52374, 60.49277, 60.46152, 60.42997, 60.39814, 
    60.36602, 60.33362, 60.30093, 60.26795, 60.23469, 60.20115, 60.16733, 
    60.13322, 60.09884, 60.06418, 60.02924, 59.99402, 59.95853, 59.92276, 
    59.88673, 59.85041, 59.81383, 59.77697, 59.73985, 59.70245, 59.66479, 
    59.62687, 59.58867, 59.55021, 59.51149, 59.47251, 59.43327, 59.39376, 
    59.354, 59.31397, 59.27369, 59.23315, 59.19236, 59.15132, 59.11002, 
    59.06847, 59.02667, 58.98462, 58.94231, 58.89977, 58.85697, 58.81393, 
    58.77065, 58.72712, 58.68334, 58.63933, 58.59508, 58.55058, 58.50585, 
    58.46088, 58.41568, 58.37024, 58.32456, 58.27865, 58.23251, 58.18614, 
    58.13954, 58.0927, 58.04565, 57.99836, 57.95085, 57.90311, 57.85515, 
    57.80697, 57.75857, 57.70994, 57.66109, 57.61203, 57.56275, 57.51325, 
    57.46354, 57.41361,
  52.0635, 52.12935, 52.19507, 52.26065, 52.32611, 52.39143, 52.45662, 
    52.52167, 52.58658, 52.65136, 52.716, 52.7805, 52.84486, 52.90909, 
    52.97317, 53.03711, 53.10091, 53.16457, 53.22808, 53.29145, 53.35468, 
    53.41775, 53.48068, 53.54346, 53.6061, 53.66858, 53.73092, 53.7931, 
    53.85513, 53.91701, 53.97873, 54.0403, 54.10172, 54.16298, 54.22408, 
    54.28503, 54.34581, 54.40644, 54.4669, 54.52721, 54.58735, 54.64734, 
    54.70715, 54.7668, 54.82629, 54.88561, 54.94476, 55.00374, 55.06256, 
    55.1212, 55.17968, 55.23798, 55.29611, 55.35406, 55.41185, 55.46945, 
    55.52688, 55.58413, 55.6412, 55.6981, 55.75481, 55.81134, 55.86769, 
    55.92386, 55.97984, 56.03564, 56.09126, 56.14668, 56.20192, 56.25697, 
    56.31183, 56.3665, 56.42097, 56.47526, 56.52935, 56.58324, 56.63694, 
    56.69045, 56.74376, 56.79686, 56.84977, 56.90248, 56.95498, 57.00729, 
    57.05939, 57.11128, 57.16297, 57.21445, 57.26573, 57.3168, 57.36766, 
    57.4183, 57.46873, 57.51896, 57.56897, 57.61876, 57.66834, 57.7177, 
    57.76684, 57.81577, 57.86447, 57.91295, 57.96121, 58.00925, 58.05706, 
    58.10466, 58.15202, 58.19915, 58.24606, 58.29274, 58.33918, 58.3854, 
    58.43139, 58.47713, 58.52265, 58.56793, 58.61297, 58.65778, 58.70234, 
    58.74667, 58.79076, 58.8346, 58.8782, 58.92155, 58.96467, 59.00753, 
    59.05015, 59.09252, 59.13464, 59.17651, 59.21813, 59.25949, 59.30061, 
    59.34146, 59.38206, 59.42241, 59.4625, 59.50232, 59.54189, 59.5812, 
    59.62025, 59.65903, 59.69755, 59.7358, 59.77379, 59.81151, 59.84896, 
    59.88615, 59.92306, 59.9597, 59.99607, 60.03217, 60.06799, 60.10353, 
    60.1388, 60.1738, 60.20851, 60.24295, 60.2771, 60.31097, 60.34457, 
    60.37787, 60.4109, 60.44363, 60.47609, 60.50825, 60.54013, 60.57172, 
    60.60301, 60.63402, 60.66473, 60.69516, 60.72528, 60.75512, 60.78465, 
    60.8139, 60.84284, 60.87148, 60.89983, 60.92787, 60.95562, 60.98306, 
    61.0102, 61.03703, 61.06356, 61.08979, 61.11571, 61.14132, 61.16662, 
    61.19162, 61.2163, 61.24068, 61.26474, 61.28849, 61.31193, 61.33506, 
    61.35786, 61.38036, 61.40254, 61.4244, 61.44595, 61.46717, 61.48808, 
    61.50867, 61.52893, 61.54888, 61.56851, 61.58781, 61.60679, 61.62544, 
    61.64378, 61.66178, 61.67946, 61.69682, 61.71384, 61.73054, 61.74691, 
    61.76295, 61.77867, 61.79405, 61.8091, 61.82383, 61.83822, 61.85228, 
    61.866, 61.87939, 61.89246, 61.90518, 61.91757, 61.92963, 61.94135, 
    61.95273, 61.96378, 61.97449, 61.98487, 61.99491, 62.00461, 62.01397, 
    62.02299, 62.03168, 62.04003, 62.04803, 62.0557, 62.06303, 62.07002, 
    62.07666, 62.08297, 62.08894, 62.09456, 62.09984, 62.10478, 62.10938, 
    62.11364, 62.11755, 62.12112, 62.12435, 62.12724, 62.12978, 62.13199, 
    62.13385, 62.13536, 62.13654, 62.13737, 62.13786, 62.138, 62.1378, 
    62.13726, 62.13638, 62.13515, 62.13358, 62.13166, 62.12941, 62.12681, 
    62.12386, 62.12058, 62.11695, 62.11298, 62.10867, 62.10402, 62.09903, 
    62.09369, 62.08801, 62.08199, 62.07563, 62.06894, 62.06189, 62.05451, 
    62.04679, 62.03873, 62.03033, 62.02159, 62.01252, 62.0031, 61.99334, 
    61.98325, 61.97282, 61.96206, 61.95095, 61.93952, 61.92774, 61.91563, 
    61.90319, 61.89041, 61.8773, 61.86385, 61.85007, 61.83596, 61.82152, 
    61.80674, 61.79164, 61.7762, 61.76044, 61.74434, 61.72792, 61.71117, 
    61.69409, 61.67669, 61.65895, 61.6409, 61.62251, 61.60381, 61.58478, 
    61.56542, 61.54575, 61.52575, 61.50543, 61.48479, 61.46384, 61.44256, 
    61.42096, 61.39905, 61.37682, 61.35428, 61.33142, 61.30824, 61.28476, 
    61.26096, 61.23684, 61.21242, 61.18768, 61.16264, 61.13729, 61.11163, 
    61.08566, 61.05939, 61.03281, 61.00592, 60.97874, 60.95125, 60.92346, 
    60.89536, 60.86697, 60.83828, 60.80929, 60.78, 60.75042, 60.72054, 
    60.69036, 60.6599, 60.62914, 60.59808, 60.56674, 60.53511, 60.50318, 
    60.47097, 60.43848, 60.40569, 60.37262, 60.33927, 60.30563, 60.27172, 
    60.23752, 60.20304, 60.16828, 60.13324, 60.09793, 60.06234, 60.02647, 
    59.99033, 59.95392, 59.91724, 59.88028, 59.84306, 59.80556, 59.7678, 
    59.72977, 59.69147, 59.65291, 59.61409, 59.575, 59.53565, 59.49604, 
    59.45617, 59.41605, 59.37566, 59.33501, 59.29412, 59.25297, 59.21156, 
    59.1699, 59.12799, 59.08583, 59.04342, 59.00077, 58.95786, 58.91471, 
    58.87132, 58.82768, 58.7838, 58.73967, 58.69531, 58.6507, 58.60586, 
    58.56078, 58.51546, 58.46991, 58.42413, 58.37811, 58.33185, 58.28537, 
    58.23866, 58.19171, 58.14454, 58.09714, 58.04952, 58.00167, 57.95359, 
    57.9053, 57.85678, 57.80804, 57.75908, 57.7099, 57.66051, 57.6109, 
    57.56107, 57.51103,
  52.1505, 52.21646, 52.28228, 52.34797, 52.41353, 52.47895, 52.54424, 
    52.6094, 52.67442, 52.7393, 52.80405, 52.86866, 52.93312, 52.99746, 
    53.06165, 53.12569, 53.1896, 53.25336, 53.31698, 53.38046, 53.44379, 
    53.50697, 53.57001, 53.6329, 53.69564, 53.75824, 53.82068, 53.88297, 
    53.94511, 54.0071, 54.06894, 54.13062, 54.19214, 54.25351, 54.31473, 
    54.37578, 54.43668, 54.49742, 54.55799, 54.61841, 54.67867, 54.73876, 
    54.79869, 54.85845, 54.91805, 54.97748, 55.03674, 55.09584, 55.15477, 
    55.21353, 55.27211, 55.33053, 55.38877, 55.44684, 55.50473, 55.56245, 
    55.62, 55.67736, 55.73455, 55.79155, 55.84838, 55.90503, 55.96149, 
    56.01778, 56.07388, 56.12979, 56.18551, 56.24105, 56.29641, 56.35157, 
    56.40654, 56.46133, 56.51592, 56.57032, 56.62453, 56.67854, 56.73235, 
    56.78597, 56.83939, 56.89262, 56.94564, 56.99846, 57.05108, 57.1035, 
    57.15572, 57.20773, 57.25953, 57.31113, 57.36252, 57.4137, 57.46467, 
    57.51543, 57.56598, 57.61632, 57.66644, 57.71635, 57.76604, 57.81552, 
    57.86478, 57.91381, 57.96264, 58.01123, 58.0596, 58.10776, 58.15569, 
    58.20339, 58.25086, 58.29811, 58.34513, 58.39192, 58.43848, 58.48481, 
    58.53091, 58.57677, 58.62239, 58.66779, 58.71294, 58.75786, 58.80254, 
    58.84697, 58.89117, 58.93512, 58.97883, 59.0223, 59.06552, 59.10849, 
    59.15122, 59.1937, 59.23593, 59.2779, 59.31963, 59.3611, 59.40232, 
    59.44329, 59.484, 59.52445, 59.56464, 59.60458, 59.64425, 59.68366, 
    59.72281, 59.7617, 59.80032, 59.83868, 59.87677, 59.91459, 59.95214, 
    59.98943, 60.02644, 60.06318, 60.09965, 60.13585, 60.17177, 60.20741, 
    60.24278, 60.27787, 60.31268, 60.34721, 60.38147, 60.41544, 60.44912, 
    60.48252, 60.51564, 60.54847, 60.58102, 60.61327, 60.64524, 60.67692, 
    60.70831, 60.7394, 60.77021, 60.80072, 60.83093, 60.86085, 60.89048, 
    60.9198, 60.94883, 60.97756, 61.00599, 61.03411, 61.06194, 61.08947, 
    61.11668, 61.1436, 61.17021, 61.19651, 61.22251, 61.2482, 61.27358, 
    61.29865, 61.32341, 61.34786, 61.37199, 61.39582, 61.41933, 61.44252, 
    61.4654, 61.48796, 61.51021, 61.53214, 61.55375, 61.57505, 61.59602, 
    61.61667, 61.637, 61.65701, 61.67669, 61.69606, 61.7151, 61.73381, 
    61.7522, 61.77026, 61.78799, 61.8054, 61.82248, 61.83923, 61.85566, 
    61.87175, 61.88752, 61.90295, 61.91805, 61.93282, 61.94725, 61.96136, 
    61.97512, 61.98856, 62.00166, 62.01443, 62.02686, 62.03896, 62.05071, 
    62.06213, 62.07322, 62.08397, 62.09438, 62.10445, 62.11418, 62.12357, 
    62.13263, 62.14134, 62.14971, 62.15775, 62.16544, 62.17279, 62.17979, 
    62.18646, 62.19279, 62.19878, 62.20442, 62.20972, 62.21467, 62.21929, 
    62.22356, 62.22749, 62.23107, 62.23431, 62.23721, 62.23976, 62.24197, 
    62.24383, 62.24535, 62.24653, 62.24736, 62.24785, 62.248, 62.2478, 
    62.24726, 62.24637, 62.24514, 62.24356, 62.24164, 62.23938, 62.23677, 
    62.23382, 62.23053, 62.22689, 62.2229, 62.21858, 62.21391, 62.2089, 
    62.20355, 62.19785, 62.19181, 62.18543, 62.17871, 62.17165, 62.16424, 
    62.15649, 62.14841, 62.13998, 62.13121, 62.12211, 62.11266, 62.10287, 
    62.09275, 62.08229, 62.07149, 62.06035, 62.04887, 62.03706, 62.02491, 
    62.01243, 61.99961, 61.98646, 61.97297, 61.95915, 61.94499, 61.9305, 
    61.91568, 61.90053, 61.88504, 61.86923, 61.85308, 61.83661, 61.8198, 
    61.80267, 61.78521, 61.76742, 61.74931, 61.73087, 61.7121, 61.69302, 
    61.6736, 61.65387, 61.6338, 61.61342, 61.59272, 61.5717, 61.55036, 
    61.52869, 61.50671, 61.48442, 61.4618, 61.43887, 61.41563, 61.39207, 
    61.3682, 61.34401, 61.31952, 61.2947, 61.26958, 61.24416, 61.21842, 
    61.19238, 61.16602, 61.13936, 61.1124, 61.08513, 61.05756, 61.02969, 
    61.00151, 60.97303, 60.94426, 60.91518, 60.88581, 60.85614, 60.82617, 
    60.79591, 60.76535, 60.7345, 60.70336, 60.67193, 60.64021, 60.60819, 
    60.57589, 60.5433, 60.51042, 60.47726, 60.44381, 60.41008, 60.37607, 
    60.34177, 60.3072, 60.27234, 60.23721, 60.20179, 60.16611, 60.13014, 
    60.0939, 60.05739, 60.0206, 59.98355, 59.94622, 59.90862, 59.87076, 
    59.83263, 59.79423, 59.75557, 59.71664, 59.67744, 59.63799, 59.59827, 
    59.5583, 59.51807, 59.47757, 59.43682, 59.39582, 59.35456, 59.31305, 
    59.27128, 59.22926, 59.187, 59.14448, 59.10171, 59.0587, 59.01544, 
    58.97194, 58.92818, 58.88419, 58.83996, 58.79548, 58.75077, 58.70581, 
    58.66062, 58.61519, 58.56953, 58.52363, 58.4775, 58.43113, 58.38454, 
    58.33771, 58.29065, 58.24337, 58.19586, 58.14812, 58.10015, 58.05197, 
    58.00356, 57.95493, 57.90607, 57.857, 57.80771, 57.7582, 57.70847, 
    57.65853, 57.60837,
  52.23741, 52.30346, 52.36939, 52.43518, 52.50085, 52.56638, 52.63177, 
    52.69703, 52.76216, 52.82714, 52.892, 52.95671, 53.02129, 53.08572, 
    53.15002, 53.21417, 53.27819, 53.34206, 53.40578, 53.46937, 53.53281, 
    53.5961, 53.65924, 53.72224, 53.7851, 53.8478, 53.91035, 53.97275, 
    54.035, 54.0971, 54.15905, 54.22084, 54.28247, 54.34395, 54.40528, 
    54.46644, 54.52745, 54.5883, 54.64899, 54.70952, 54.76988, 54.83009, 
    54.89013, 54.95, 55.00972, 55.06926, 55.12864, 55.18785, 55.24689, 
    55.30576, 55.36446, 55.42299, 55.48134, 55.53952, 55.59753, 55.65536, 
    55.71302, 55.7705, 55.8278, 55.88493, 55.94187, 55.99863, 56.05521, 
    56.11161, 56.16782, 56.22385, 56.27969, 56.33534, 56.39081, 56.44609, 
    56.50118, 56.55608, 56.61079, 56.6653, 56.71962, 56.77375, 56.82768, 
    56.88142, 56.93495, 56.98829, 57.04143, 57.09437, 57.1471, 57.19964, 
    57.25197, 57.3041, 57.35601, 57.40773, 57.45923, 57.51053, 57.56162, 
    57.6125, 57.66316, 57.71361, 57.76385, 57.81387, 57.86368, 57.91327, 
    57.96264, 58.0118, 58.06073, 58.10944, 58.15793, 58.2062, 58.25424, 
    58.30205, 58.34964, 58.397, 58.44414, 58.49104, 58.53772, 58.58416, 
    58.63037, 58.67634, 58.72208, 58.76758, 58.81285, 58.85788, 58.90267, 
    58.94722, 58.99152, 59.03559, 59.07941, 59.12299, 59.16632, 59.2094, 
    59.25224, 59.29483, 59.33716, 59.37925, 59.42108, 59.46267, 59.50399, 
    59.54506, 59.58588, 59.62644, 59.66674, 59.70678, 59.74656, 59.78607, 
    59.82533, 59.86432, 59.90305, 59.94151, 59.9797, 60.01762, 60.05528, 
    60.09267, 60.12978, 60.16663, 60.20319, 60.23949, 60.27551, 60.31126, 
    60.34672, 60.38191, 60.41682, 60.45145, 60.48579, 60.51986, 60.55364, 
    60.58714, 60.62035, 60.65327, 60.68591, 60.71826, 60.75032, 60.78209, 
    60.81357, 60.84476, 60.87565, 60.90625, 60.93655, 60.96656, 60.99627, 
    61.02568, 61.05479, 61.08361, 61.11212, 61.14034, 61.16824, 61.19585, 
    61.22315, 61.25014, 61.27683, 61.30322, 61.32929, 61.35506, 61.38052, 
    61.40566, 61.4305, 61.45502, 61.47923, 61.50312, 61.52671, 61.54997, 
    61.57292, 61.59555, 61.61787, 61.63987, 61.66154, 61.6829, 61.70394, 
    61.72466, 61.74505, 61.76512, 61.78487, 61.80429, 61.82339, 61.84216, 
    61.86061, 61.87873, 61.89652, 61.91398, 61.93111, 61.94792, 61.96439, 
    61.98054, 61.99635, 62.01183, 62.02698, 62.0418, 62.05628, 62.07043, 
    62.08424, 62.09772, 62.11087, 62.12367, 62.13614, 62.14828, 62.16007, 
    62.17153, 62.18265, 62.19344, 62.20388, 62.21398, 62.22374, 62.23317, 
    62.24225, 62.25099, 62.25939, 62.26745, 62.27517, 62.28254, 62.28957, 
    62.29626, 62.30261, 62.30861, 62.31427, 62.31959, 62.32456, 62.32919, 
    62.33348, 62.33742, 62.34101, 62.34426, 62.34717, 62.34973, 62.35195, 
    62.35382, 62.35535, 62.35653, 62.35736, 62.35785, 62.358, 62.3578, 
    62.35725, 62.35636, 62.35513, 62.35355, 62.35162, 62.34935, 62.34673, 
    62.34377, 62.34047, 62.33682, 62.33282, 62.32848, 62.3238, 62.31877, 
    62.3134, 62.30769, 62.30163, 62.29523, 62.28848, 62.2814, 62.27397, 
    62.2662, 62.25808, 62.24963, 62.24083, 62.2317, 62.22222, 62.2124, 
    62.20225, 62.19175, 62.18092, 62.16974, 62.15823, 62.14638, 62.13419, 
    62.12167, 62.10881, 62.09561, 62.08208, 62.06821, 62.05401, 62.03948, 
    62.02461, 62.00941, 61.99387, 61.97801, 61.96181, 61.94529, 61.92843, 
    61.91124, 61.89373, 61.87588, 61.85771, 61.83921, 61.82039, 61.80124, 
    61.78176, 61.76197, 61.74184, 61.7214, 61.70063, 61.67955, 61.65814, 
    61.63641, 61.61436, 61.592, 61.56931, 61.54631, 61.52299, 61.49937, 
    61.47542, 61.45116, 61.42659, 61.4017, 61.37651, 61.351, 61.32519, 
    61.29906, 61.27263, 61.2459, 61.21885, 61.1915, 61.16385, 61.13589, 
    61.10763, 61.07907, 61.05021, 61.02105, 60.99159, 60.96183, 60.93178, 
    60.90143, 60.87078, 60.83984, 60.80861, 60.77708, 60.74527, 60.71317, 
    60.68077, 60.64809, 60.61512, 60.58186, 60.54832, 60.51449, 60.48038, 
    60.44599, 60.41132, 60.37636, 60.34113, 60.30562, 60.26983, 60.23377, 
    60.19743, 60.16082, 60.12393, 60.08677, 60.04934, 60.01164, 59.97367, 
    59.93544, 59.89694, 59.85817, 59.81914, 59.77984, 59.74028, 59.70046, 
    59.66038, 59.62004, 59.57944, 59.53858, 59.49747, 59.4561, 59.41448, 
    59.37261, 59.33048, 59.28811, 59.24548, 59.2026, 59.15948, 59.11611, 
    59.07249, 59.02863, 58.98453, 58.94019, 58.8956, 58.85077, 58.80571, 
    58.7604, 58.71486, 58.66908, 58.62307, 58.57683, 58.53035, 58.48364, 
    58.4367, 58.38953, 58.34213, 58.29451, 58.24665, 58.19857, 58.15027, 
    58.10175, 58.053, 58.00404, 57.95485, 57.90544, 57.85582, 57.80597, 
    57.75592, 57.70565,
  52.32421, 52.39037, 52.4564, 52.5223, 52.58806, 52.6537, 52.7192, 52.78456, 
    52.84979, 52.91489, 52.97984, 53.04466, 53.10934, 53.17389, 53.23829, 
    53.30255, 53.36667, 53.43065, 53.49449, 53.55818, 53.62173, 53.68513, 
    53.74838, 53.81149, 53.87445, 53.93726, 53.99992, 54.06244, 54.12479, 
    54.187, 54.24906, 54.31096, 54.3727, 54.4343, 54.49573, 54.55701, 
    54.61813, 54.67909, 54.73989, 54.80053, 54.86101, 54.92133, 54.98148, 
    55.04147, 55.10129, 55.16095, 55.22044, 55.27976, 55.33892, 55.3979, 
    55.45671, 55.51535, 55.57383, 55.63212, 55.69024, 55.74819, 55.80596, 
    55.86356, 55.92097, 55.97821, 56.03527, 56.09214, 56.14884, 56.20535, 
    56.26168, 56.31782, 56.37378, 56.42955, 56.48513, 56.54053, 56.59573, 
    56.65075, 56.70557, 56.7602, 56.81464, 56.86888, 56.92293, 56.97678, 
    57.03043, 57.08389, 57.13714, 57.19019, 57.24305, 57.2957, 57.34814, 
    57.40039, 57.45242, 57.50425, 57.55587, 57.60728, 57.65849, 57.70948, 
    57.76026, 57.81083, 57.86118, 57.91132, 57.96125, 58.01095, 58.06044, 
    58.10971, 58.15875, 58.20758, 58.25618, 58.30457, 58.35272, 58.40065, 
    58.44836, 58.49583, 58.54308, 58.5901, 58.63689, 58.68344, 58.72976, 
    58.77585, 58.8217, 58.86732, 58.9127, 58.95784, 59.00274, 59.0474, 
    59.09182, 59.13599, 59.17993, 59.22361, 59.26706, 59.31025, 59.3532, 
    59.3959, 59.43834, 59.48054, 59.52248, 59.56417, 59.60561, 59.64679, 
    59.68771, 59.72837, 59.76878, 59.80893, 59.84881, 59.88844, 59.9278, 
    59.96689, 60.00572, 60.04429, 60.08258, 60.12061, 60.15837, 60.19586, 
    60.23308, 60.27002, 60.30669, 60.34309, 60.37921, 60.41505, 60.45062, 
    60.48591, 60.52092, 60.55564, 60.59008, 60.62425, 60.65812, 60.69172, 
    60.72503, 60.75804, 60.79078, 60.82322, 60.85537, 60.88723, 60.9188, 
    60.95008, 60.98106, 61.01175, 61.04214, 61.07224, 61.10204, 61.13153, 
    61.16073, 61.18963, 61.21823, 61.24652, 61.27452, 61.3022, 61.32959, 
    61.35667, 61.38343, 61.4099, 61.43605, 61.46189, 61.48743, 61.51265, 
    61.53756, 61.56216, 61.58644, 61.61041, 61.63406, 61.6574, 61.68042, 
    61.70313, 61.72551, 61.74758, 61.76932, 61.79074, 61.81185, 61.83263, 
    61.85308, 61.87322, 61.89303, 61.91251, 61.93167, 61.9505, 61.96901, 
    61.98718, 62.00503, 62.02255, 62.03974, 62.05659, 62.07312, 62.08932, 
    62.10518, 62.12071, 62.13591, 62.15077, 62.1653, 62.1795, 62.19336, 
    62.20687, 62.22006, 62.23291, 62.24542, 62.2576, 62.26943, 62.28093, 
    62.29208, 62.3029, 62.31337, 62.32351, 62.33331, 62.34276, 62.35187, 
    62.36064, 62.36907, 62.37715, 62.3849, 62.3923, 62.39935, 62.40606, 
    62.41243, 62.41845, 62.42413, 62.42947, 62.43445, 62.4391, 62.4434, 
    62.44735, 62.45096, 62.45422, 62.45713, 62.45971, 62.46193, 62.46381, 
    62.46534, 62.46652, 62.46736, 62.46785, 62.468, 62.4678, 62.46725, 
    62.46636, 62.46512, 62.46353, 62.4616, 62.45932, 62.4567, 62.45373, 
    62.45041, 62.44675, 62.44274, 62.43839, 62.43369, 62.42864, 62.42326, 
    62.41752, 62.41145, 62.40502, 62.39826, 62.39115, 62.38369, 62.3759, 
    62.36776, 62.35928, 62.35045, 62.34129, 62.33178, 62.32193, 62.31174, 
    62.30121, 62.29034, 62.27913, 62.26758, 62.25569, 62.24347, 62.2309, 
    62.218, 62.20476, 62.19118, 62.17727, 62.16302, 62.14845, 62.13353, 
    62.11828, 62.1027, 62.08678, 62.07053, 62.05395, 62.03704, 62.0198, 
    62.00223, 61.98433, 61.9661, 61.94754, 61.92866, 61.90945, 61.88992, 
    61.87006, 61.84987, 61.82936, 61.80853, 61.78738, 61.7659, 61.74411, 
    61.72199, 61.69956, 61.6768, 61.65373, 61.63034, 61.60664, 61.58262, 
    61.55829, 61.53364, 61.50868, 61.48341, 61.45783, 61.43193, 61.40573, 
    61.37922, 61.3524, 61.32528, 61.29784, 61.27011, 61.24207, 61.21373, 
    61.18508, 61.15614, 61.12689, 61.09734, 61.0675, 61.03735, 61.00691, 
    60.97618, 60.94515, 60.91383, 60.88221, 60.8503, 60.8181, 60.78562, 
    60.75284, 60.71977, 60.68642, 60.65279, 60.61886, 60.58466, 60.55017, 
    60.5154, 60.48035, 60.44501, 60.4094, 60.37352, 60.33735, 60.30091, 
    60.2642, 60.22721, 60.18995, 60.15242, 60.11462, 60.07655, 60.0382, 
    59.9996, 59.96073, 59.92159, 59.88219, 59.84252, 59.80259, 59.76241, 
    59.72196, 59.68125, 59.64029, 59.59907, 59.55759, 59.51587, 59.47388, 
    59.43164, 59.38916, 59.34642, 59.30344, 59.2602, 59.21672, 59.173, 
    59.12902, 59.08481, 59.04035, 58.99565, 58.95071, 58.90554, 58.86012, 
    58.81446, 58.76857, 58.72245, 58.67609, 58.6295, 58.58268, 58.53562, 
    58.48834, 58.44083, 58.39309, 58.34512, 58.29693, 58.24851, 58.19987, 
    58.15101, 58.10193, 58.05262, 58.0031, 57.95336, 57.9034, 57.85323, 
    57.80285,
  52.4109, 52.47717, 52.5433, 52.60931, 52.67518, 52.74092, 52.80652, 
    52.87199, 52.93733, 53.00253, 53.06759, 53.13251, 53.1973, 53.26196, 
    53.32646, 53.39083, 53.45506, 53.51915, 53.58309, 53.64689, 53.71054, 
    53.77406, 53.83742, 53.90063, 53.9637, 54.02663, 54.0894, 54.15202, 
    54.21449, 54.27681, 54.33897, 54.40099, 54.46284, 54.52454, 54.58609, 
    54.64748, 54.70871, 54.76978, 54.8307, 54.89145, 54.95204, 55.01247, 
    55.07273, 55.13284, 55.19277, 55.25254, 55.31215, 55.37158, 55.43085, 
    55.48995, 55.54888, 55.60764, 55.66622, 55.72463, 55.78287, 55.84093, 
    55.89882, 55.95652, 56.01405, 56.07141, 56.12858, 56.18557, 56.24238, 
    56.29901, 56.35545, 56.41171, 56.46778, 56.52367, 56.57937, 56.63488, 
    56.6902, 56.74533, 56.80027, 56.85502, 56.90957, 56.96393, 57.01809, 
    57.07206, 57.12583, 57.1794, 57.23277, 57.28594, 57.33891, 57.39168, 
    57.44424, 57.4966, 57.54875, 57.6007, 57.65244, 57.70396, 57.75528, 
    57.80639, 57.85729, 57.90797, 57.95844, 58.0087, 58.05874, 58.10856, 
    58.15816, 58.20755, 58.25671, 58.30565, 58.35437, 58.40287, 58.45114, 
    58.49918, 58.547, 58.59459, 58.64196, 58.68909, 58.73599, 58.78266, 
    58.82909, 58.87529, 58.92126, 58.96699, 59.01248, 59.05774, 59.10275, 
    59.14753, 59.19205, 59.23634, 59.28039, 59.32419, 59.36774, 59.41105, 
    59.4541, 59.49691, 59.53947, 59.58177, 59.62383, 59.66563, 59.70717, 
    59.74846, 59.78949, 59.83026, 59.87077, 59.91103, 59.95102, 59.99075, 
    60.03022, 60.06942, 60.10836, 60.14703, 60.18542, 60.22356, 60.26142, 
    60.29902, 60.33633, 60.37338, 60.41015, 60.44665, 60.48287, 60.51881, 
    60.55448, 60.58987, 60.62497, 60.6598, 60.69434, 60.7286, 60.76257, 
    60.79626, 60.82966, 60.86278, 60.8956, 60.92814, 60.96038, 60.99234, 
    61.024, 61.05537, 61.08644, 61.11722, 61.1477, 61.17788, 61.20777, 
    61.23736, 61.26664, 61.29563, 61.32431, 61.35269, 61.38077, 61.40854, 
    61.436, 61.46316, 61.49001, 61.51655, 61.54279, 61.56871, 61.59432, 
    61.61962, 61.64461, 61.66928, 61.69364, 61.71768, 61.74141, 61.76482, 
    61.78791, 61.81068, 61.83314, 61.85527, 61.87708, 61.89857, 61.91974, 
    61.94059, 61.96111, 61.9813, 62.00117, 62.02072, 62.03994, 62.05883, 
    62.07739, 62.09563, 62.11353, 62.13111, 62.14835, 62.16526, 62.18184, 
    62.19809, 62.214, 62.22958, 62.24483, 62.25974, 62.27431, 62.28856, 
    62.30246, 62.31602, 62.32925, 62.34214, 62.35469, 62.36691, 62.37878, 
    62.39031, 62.4015, 62.41236, 62.42287, 62.43304, 62.44286, 62.45235, 
    62.46149, 62.47029, 62.47874, 62.48685, 62.49462, 62.50204, 62.50912, 
    62.51586, 62.52225, 62.52829, 62.53399, 62.53934, 62.54434, 62.549, 
    62.55331, 62.55728, 62.5609, 62.56417, 62.5671, 62.56968, 62.57191, 
    62.57379, 62.57533, 62.57652, 62.57736, 62.57785, 62.578, 62.5778, 
    62.57725, 62.57635, 62.57511, 62.57352, 62.57158, 62.56929, 62.56666, 
    62.56368, 62.56035, 62.55668, 62.55266, 62.54829, 62.54358, 62.53851, 
    62.53311, 62.52736, 62.52126, 62.51482, 62.50803, 62.50089, 62.49342, 
    62.4856, 62.47743, 62.46892, 62.46007, 62.45087, 62.44133, 62.43145, 
    62.42123, 62.41066, 62.39976, 62.38851, 62.37692, 62.365, 62.35273, 
    62.34013, 62.32718, 62.3139, 62.30028, 62.28633, 62.27203, 62.2574, 
    62.24244, 62.22714, 62.21151, 62.19554, 62.17924, 62.16261, 62.14565, 
    62.12835, 62.11072, 62.09277, 62.07448, 62.05587, 62.03692, 62.01765, 
    61.99805, 61.97813, 61.95789, 61.93731, 61.91642, 61.8952, 61.87365, 
    61.85179, 61.82961, 61.8071, 61.78428, 61.76114, 61.73767, 61.7139, 
    61.6898, 61.6654, 61.64067, 61.61564, 61.59029, 61.56463, 61.53866, 
    61.51237, 61.48578, 61.45889, 61.43168, 61.40416, 61.37635, 61.34822, 
    61.31979, 61.29106, 61.26203, 61.2327, 61.20306, 61.17313, 61.1429, 
    61.11237, 61.08155, 61.05043, 61.01901, 60.9873, 60.9553, 60.92301, 
    60.89043, 60.85756, 60.8244, 60.79095, 60.75722, 60.7232, 60.68889, 
    60.65431, 60.61944, 60.58429, 60.54886, 60.51315, 60.47716, 60.4409, 
    60.40435, 60.36754, 60.33045, 60.29308, 60.25545, 60.21754, 60.17937, 
    60.14093, 60.10221, 60.06324, 60.02399, 59.98449, 59.94471, 59.90468, 
    59.86438, 59.82383, 59.78302, 59.74194, 59.70061, 59.65903, 59.61719, 
    59.5751, 59.53275, 59.49015, 59.44731, 59.40421, 59.36087, 59.31728, 
    59.27344, 59.22935, 59.18503, 59.14046, 59.09565, 59.05059, 59.0053, 
    58.95977, 58.91401, 58.868, 58.82177, 58.77529, 58.72858, 58.68165, 
    58.63448, 58.58708, 58.53945, 58.4916, 58.44352, 58.39521, 58.34668, 
    58.29792, 58.24895, 58.19975, 58.15033, 58.10069, 58.05083, 58.00076, 
    57.95047, 57.89997,
  52.4975, 52.56387, 52.6301, 52.69621, 52.76219, 52.82803, 52.89374, 
    52.95932, 53.02476, 53.09007, 53.15524, 53.22027, 53.28516, 53.34992, 
    53.41454, 53.47901, 53.54335, 53.60754, 53.67159, 53.7355, 53.79926, 
    53.86288, 53.92635, 53.98968, 54.05286, 54.11589, 54.17877, 54.2415, 
    54.30408, 54.36651, 54.42879, 54.49091, 54.55288, 54.61469, 54.67635, 
    54.73785, 54.7992, 54.86038, 54.92141, 54.98227, 55.04298, 55.10352, 
    55.16389, 55.22411, 55.28416, 55.34404, 55.40376, 55.46331, 55.52269, 
    55.58191, 55.64095, 55.69982, 55.75852, 55.81704, 55.8754, 55.93357, 
    55.99157, 56.0494, 56.10704, 56.16451, 56.2218, 56.27891, 56.33583, 
    56.39258, 56.44913, 56.50551, 56.5617, 56.6177, 56.67352, 56.72915, 
    56.78458, 56.83983, 56.89489, 56.94975, 57.00442, 57.0589, 57.11318, 
    57.16726, 57.22115, 57.27483, 57.32832, 57.38161, 57.4347, 57.48758, 
    57.54026, 57.59274, 57.645, 57.69707, 57.74892, 57.80057, 57.85201, 
    57.90323, 57.95424, 58.00504, 58.05563, 58.106, 58.15615, 58.20609, 
    58.25581, 58.30531, 58.35459, 58.40365, 58.45249, 58.5011, 58.54948, 
    58.59764, 58.64558, 58.69329, 58.74076, 58.78801, 58.83503, 58.88181, 
    58.92836, 58.97468, 59.02076, 59.0666, 59.11221, 59.15757, 59.2027, 
    59.24759, 59.29223, 59.33663, 59.38079, 59.4247, 59.46836, 59.51178, 
    59.55495, 59.59787, 59.64054, 59.68295, 59.72512, 59.76702, 59.80868, 
    59.85007, 59.89122, 59.93209, 59.97272, 60.01308, 60.05318, 60.09302, 
    60.13259, 60.1719, 60.21094, 60.24971, 60.28822, 60.32646, 60.36443, 
    60.40212, 60.43954, 60.47669, 60.51357, 60.55017, 60.58649, 60.62253, 
    60.6583, 60.69379, 60.72899, 60.76391, 60.79855, 60.83291, 60.86698, 
    60.90076, 60.93427, 60.96747, 61.00039, 61.03302, 61.06536, 61.09741, 
    61.12917, 61.16063, 61.19179, 61.22266, 61.25323, 61.2835, 61.31348, 
    61.34315, 61.37252, 61.4016, 61.43036, 61.45883, 61.48699, 61.51484, 
    61.54239, 61.56963, 61.59657, 61.62319, 61.6495, 61.6755, 61.70119, 
    61.72657, 61.75163, 61.77638, 61.80081, 61.82493, 61.84873, 61.87221, 
    61.89537, 61.91822, 61.94074, 61.96295, 61.98483, 62.00639, 62.02762, 
    62.04853, 62.06912, 62.08938, 62.10931, 62.12892, 62.1482, 62.16715, 
    62.18577, 62.20406, 62.22202, 62.23965, 62.25695, 62.27392, 62.29055, 
    62.30685, 62.32281, 62.33845, 62.35374, 62.3687, 62.38332, 62.39761, 
    62.41156, 62.42517, 62.43844, 62.45137, 62.46396, 62.47621, 62.48812, 
    62.49969, 62.51093, 62.52181, 62.53236, 62.54256, 62.55242, 62.56193, 
    62.57111, 62.57993, 62.58842, 62.59655, 62.60435, 62.61179, 62.6189, 
    62.62565, 62.63206, 62.63813, 62.64384, 62.64921, 62.65423, 62.65891, 
    62.66323, 62.66721, 62.67085, 62.67413, 62.67706, 62.67965, 62.68189, 
    62.68378, 62.68532, 62.68651, 62.68736, 62.68785, 62.688, 62.6878, 
    62.68725, 62.68635, 62.6851, 62.6835, 62.68156, 62.67926, 62.67662, 
    62.67363, 62.67029, 62.66661, 62.66257, 62.65819, 62.65346, 62.64838, 
    62.64296, 62.63719, 62.63107, 62.62461, 62.6178, 62.61064, 62.60314, 
    62.59529, 62.5871, 62.57856, 62.56968, 62.56045, 62.55088, 62.54097, 
    62.53071, 62.52011, 62.50917, 62.49789, 62.48626, 62.4743, 62.46199, 
    62.44934, 62.43636, 62.42303, 62.40937, 62.39537, 62.38103, 62.36636, 
    62.35135, 62.33599, 62.32031, 62.30429, 62.28794, 62.27126, 62.25424, 
    62.23689, 62.2192, 62.20119, 62.18285, 62.16417, 62.14517, 62.12584, 
    62.10618, 62.08619, 62.06588, 62.04525, 62.02428, 62.003, 61.98139, 
    61.95945, 61.9372, 61.91463, 61.89173, 61.86852, 61.84499, 61.82114, 
    61.79697, 61.77248, 61.74769, 61.72257, 61.69715, 61.67141, 61.64536, 
    61.619, 61.59232, 61.56534, 61.53806, 61.51046, 61.48256, 61.45435, 
    61.42583, 61.39702, 61.3679, 61.33848, 61.30875, 61.27873, 61.24841, 
    61.2178, 61.18688, 61.15567, 61.12416, 61.09236, 61.06027, 61.02788, 
    60.9952, 60.96224, 60.92899, 60.89544, 60.86161, 60.8275, 60.79309, 
    60.75841, 60.72344, 60.68819, 60.65266, 60.61685, 60.58076, 60.5444, 
    60.50775, 60.47083, 60.43364, 60.39618, 60.35844, 60.32043, 60.28215, 
    60.2436, 60.20478, 60.1657, 60.12635, 60.08673, 60.04685, 60.00671, 
    59.96631, 59.92565, 59.88472, 59.84354, 59.8021, 59.76041, 59.71846, 
    59.67626, 59.6338, 59.59109, 59.54814, 59.50493, 59.46148, 59.41777, 
    59.37382, 59.32962, 59.28519, 59.2405, 59.19558, 59.15041, 59.10501, 
    59.05936, 59.01348, 58.96737, 58.92101, 58.87443, 58.82761, 58.78055, 
    58.73327, 58.68576, 58.63801, 58.59004, 58.54185, 58.49342, 58.44477, 
    58.3959, 58.34681, 58.2975, 58.24796, 58.19821, 58.14824, 58.09805, 
    58.04764, 57.99702,
  52.58399, 52.65046, 52.7168, 52.78301, 52.84909, 52.91504, 52.98086, 
    53.04654, 53.11209, 53.1775, 53.24277, 53.30791, 53.37291, 53.43778, 
    53.5025, 53.56709, 53.63153, 53.69583, 53.75999, 53.82401, 53.88788, 
    53.95161, 54.01519, 54.07863, 54.14191, 54.20506, 54.26805, 54.33089, 
    54.39358, 54.45612, 54.51851, 54.58074, 54.64282, 54.70475, 54.76652, 
    54.82813, 54.88958, 54.95088, 55.01202, 55.073, 55.13382, 55.19447, 
    55.25496, 55.31529, 55.37545, 55.43545, 55.49529, 55.55495, 55.61444, 
    55.67377, 55.73293, 55.79192, 55.85073, 55.90937, 55.96783, 56.02613, 
    56.08424, 56.14219, 56.19995, 56.25753, 56.31493, 56.37216, 56.4292, 
    56.48606, 56.54274, 56.59923, 56.65553, 56.71165, 56.76759, 56.82333, 
    56.87888, 56.93425, 56.98942, 57.0444, 57.09919, 57.15378, 57.20818, 
    57.26238, 57.31638, 57.37019, 57.42379, 57.4772, 57.5304, 57.5834, 
    57.6362, 57.68879, 57.74118, 57.79336, 57.84533, 57.89709, 57.94865, 
    57.99999, 58.05112, 58.10204, 58.15274, 58.20323, 58.2535, 58.30356, 
    58.35339, 58.40301, 58.4524, 58.50158, 58.55053, 58.59926, 58.64776, 
    58.69604, 58.74409, 58.79191, 58.8395, 58.88687, 58.934, 58.9809, 
    59.02757, 59.07399, 59.12019, 59.16615, 59.21187, 59.25735, 59.30259, 
    59.34759, 59.39235, 59.43686, 59.48113, 59.52515, 59.56893, 59.61246, 
    59.65574, 59.69877, 59.74155, 59.78408, 59.82635, 59.86837, 59.91013, 
    59.95164, 59.99289, 60.03388, 60.07461, 60.11508, 60.15528, 60.19523, 
    60.23491, 60.27433, 60.31347, 60.35236, 60.39097, 60.42931, 60.46738, 
    60.50518, 60.54271, 60.57996, 60.61694, 60.65364, 60.69006, 60.72621, 
    60.76208, 60.79766, 60.83297, 60.86799, 60.90273, 60.93718, 60.97135, 
    61.00523, 61.03883, 61.07214, 61.10515, 61.13787, 61.17031, 61.20245, 
    61.2343, 61.26585, 61.2971, 61.32806, 61.35873, 61.38909, 61.41916, 
    61.44892, 61.47838, 61.50753, 61.53639, 61.56494, 61.59319, 61.62112, 
    61.64875, 61.67608, 61.70309, 61.7298, 61.75619, 61.78227, 61.80804, 
    61.83349, 61.85863, 61.88346, 61.90797, 61.93216, 61.95603, 61.97959, 
    62.00282, 62.02574, 62.04833, 62.07061, 62.09256, 62.11418, 62.13548, 
    62.15646, 62.17711, 62.19744, 62.21743, 62.2371, 62.25644, 62.27545, 
    62.29414, 62.31248, 62.33051, 62.34819, 62.36554, 62.38256, 62.39925, 
    62.4156, 62.43162, 62.4473, 62.46265, 62.47765, 62.49232, 62.50665, 
    62.52065, 62.5343, 62.54762, 62.56059, 62.57322, 62.58551, 62.59747, 
    62.60907, 62.62034, 62.63126, 62.64184, 62.65208, 62.66197, 62.67152, 
    62.68072, 62.68958, 62.69809, 62.70625, 62.71407, 62.72154, 62.72867, 
    62.73545, 62.74187, 62.74796, 62.75369, 62.75908, 62.76412, 62.76881, 
    62.77315, 62.77715, 62.78079, 62.78408, 62.78703, 62.78962, 62.79187, 
    62.79377, 62.79531, 62.79651, 62.79736, 62.79785, 62.798, 62.7978, 
    62.79725, 62.79634, 62.79509, 62.79349, 62.79153, 62.78923, 62.78658, 
    62.78358, 62.78024, 62.77654, 62.77249, 62.76809, 62.76335, 62.75825, 
    62.75281, 62.74702, 62.74088, 62.7344, 62.72756, 62.72038, 62.71286, 
    62.70498, 62.69676, 62.6882, 62.67929, 62.67003, 62.66043, 62.65048, 
    62.64019, 62.62956, 62.61858, 62.60726, 62.5956, 62.5836, 62.57125, 
    62.55856, 62.54553, 62.53217, 62.51846, 62.50441, 62.49002, 62.4753, 
    62.46024, 62.44484, 62.42911, 62.41304, 62.39663, 62.37989, 62.36282, 
    62.34541, 62.32767, 62.3096, 62.2912, 62.27247, 62.25341, 62.23401, 
    62.21429, 62.19424, 62.17387, 62.15316, 62.13213, 62.11078, 62.0891, 
    62.0671, 62.04478, 62.02214, 61.99917, 61.97588, 61.95228, 61.92835, 
    61.90411, 61.87955, 61.85468, 61.82949, 61.80398, 61.77816, 61.75203, 
    61.72559, 61.69884, 61.67178, 61.64441, 61.61673, 61.58874, 61.56044, 
    61.53185, 61.50294, 61.47374, 61.44423, 61.41442, 61.38431, 61.3539, 
    61.32319, 61.29218, 61.26088, 61.22928, 61.19739, 61.1652, 61.13272, 
    61.09995, 61.06689, 61.03354, 60.99989, 60.96597, 60.93175, 60.89725, 
    60.86247, 60.8274, 60.79205, 60.75642, 60.72051, 60.68432, 60.64785, 
    60.61111, 60.57409, 60.53679, 60.49922, 60.46138, 60.42326, 60.38488, 
    60.34622, 60.3073, 60.26811, 60.22865, 60.18893, 60.14894, 60.1087, 
    60.06818, 60.02741, 59.98638, 59.94509, 59.90354, 59.86174, 59.81968, 
    59.77737, 59.7348, 59.69198, 59.64891, 59.60559, 59.56202, 59.51821, 
    59.47414, 59.42984, 59.38528, 59.34049, 59.29545, 59.25017, 59.20465, 
    59.15889, 59.1129, 59.06667, 59.0202, 58.9735, 58.92656, 58.87939, 
    58.83199, 58.78436, 58.7365, 58.68842, 58.64011, 58.59157, 58.5428, 
    58.49382, 58.44461, 58.39518, 58.34552, 58.29565, 58.24556, 58.19526, 
    58.14474, 58.094,
  52.67037, 52.73695, 52.80339, 52.86971, 52.93589, 53.00195, 53.06787, 
    53.13366, 53.19931, 53.26483, 53.33021, 53.39546, 53.46056, 53.52554, 
    53.59037, 53.65506, 53.71961, 53.78402, 53.84829, 53.91241, 53.9764, 
    54.04023, 54.10392, 54.16747, 54.23087, 54.29412, 54.35722, 54.42017, 
    54.48298, 54.54563, 54.60813, 54.67047, 54.73266, 54.7947, 54.85658, 
    54.91831, 54.97988, 55.04129, 55.10254, 55.16363, 55.22456, 55.28533, 
    55.34593, 55.40638, 55.46665, 55.52676, 55.58671, 55.64649, 55.7061, 
    55.76554, 55.82481, 55.88391, 55.94284, 56.0016, 56.06018, 56.11859, 
    56.17682, 56.23488, 56.29276, 56.35046, 56.40798, 56.46532, 56.52248, 
    56.57945, 56.63625, 56.69285, 56.74928, 56.80551, 56.86156, 56.91742, 
    56.97309, 57.02858, 57.08387, 57.13897, 57.19387, 57.24858, 57.3031, 
    57.35741, 57.41154, 57.46546, 57.51918, 57.5727, 57.62603, 57.67914, 
    57.73206, 57.78477, 57.83727, 57.88957, 57.94166, 57.99354, 58.04522, 
    58.09668, 58.14792, 58.19896, 58.24978, 58.30038, 58.35077, 58.40094, 
    58.4509, 58.50063, 58.55014, 58.59944, 58.64851, 58.69735, 58.74597, 
    58.79436, 58.84253, 58.89047, 58.93818, 58.98566, 59.03291, 59.07992, 
    59.1267, 59.17324, 59.21955, 59.26563, 59.31146, 59.35706, 59.40242, 
    59.44753, 59.4924, 59.53703, 59.58141, 59.62555, 59.66944, 59.71308, 
    59.75647, 59.79961, 59.84251, 59.88514, 59.92753, 59.96966, 60.01153, 
    60.05315, 60.09451, 60.13561, 60.17645, 60.21703, 60.25734, 60.29739, 
    60.33718, 60.37671, 60.41596, 60.45495, 60.49367, 60.53211, 60.57029, 
    60.6082, 60.64583, 60.68318, 60.72026, 60.75707, 60.79359, 60.82985, 
    60.86581, 60.9015, 60.9369, 60.97203, 61.00687, 61.04142, 61.07569, 
    61.10966, 61.14336, 61.17676, 61.20987, 61.24269, 61.27522, 61.30746, 
    61.3394, 61.37104, 61.40239, 61.43344, 61.4642, 61.49465, 61.5248, 
    61.55465, 61.5842, 61.61345, 61.64239, 61.67102, 61.69936, 61.72738, 
    61.75509, 61.7825, 61.8096, 61.83638, 61.86285, 61.88902, 61.91486, 
    61.9404, 61.96561, 61.99052, 62.0151, 62.03937, 62.06332, 62.08694, 
    62.11026, 62.13324, 62.15591, 62.17825, 62.20027, 62.22196, 62.24333, 
    62.26437, 62.28509, 62.30548, 62.32554, 62.34527, 62.36467, 62.38375, 
    62.40249, 62.42089, 62.43897, 62.45671, 62.47412, 62.4912, 62.50794, 
    62.52435, 62.54042, 62.55615, 62.57154, 62.5866, 62.60131, 62.61569, 
    62.62973, 62.64343, 62.65679, 62.6698, 62.68248, 62.69481, 62.7068, 
    62.71845, 62.72975, 62.74071, 62.75132, 62.76159, 62.77152, 62.7811, 
    62.79033, 62.79921, 62.80775, 62.81594, 62.82379, 62.83129, 62.83844, 
    62.84524, 62.85169, 62.85779, 62.86355, 62.86895, 62.87401, 62.87871, 
    62.88307, 62.88707, 62.89073, 62.89404, 62.89699, 62.89959, 62.90185, 
    62.90375, 62.9053, 62.9065, 62.90735, 62.90785, 62.908, 62.90779, 
    62.90724, 62.90634, 62.90508, 62.90347, 62.90152, 62.8992, 62.89655, 
    62.89354, 62.89017, 62.88646, 62.8824, 62.87799, 62.87323, 62.86812, 
    62.86266, 62.85685, 62.85069, 62.84418, 62.83733, 62.83012, 62.82257, 
    62.81467, 62.80643, 62.79783, 62.78889, 62.77961, 62.76997, 62.75999, 
    62.74967, 62.739, 62.72799, 62.71663, 62.70493, 62.69288, 62.6805, 
    62.66777, 62.6547, 62.64128, 62.62753, 62.61344, 62.59901, 62.58424, 
    62.56913, 62.55368, 62.5379, 62.52177, 62.50532, 62.48852, 62.47139, 
    62.45393, 62.43613, 62.41801, 62.39954, 62.38075, 62.36163, 62.34217, 
    62.32239, 62.30228, 62.28183, 62.26107, 62.23997, 62.21855, 62.19681, 
    62.17474, 62.15234, 62.12963, 62.10659, 62.08323, 62.05955, 62.03555, 
    62.01123, 61.9866, 61.96165, 61.93638, 61.9108, 61.8849, 61.85869, 
    61.83216, 61.80533, 61.77819, 61.75073, 61.72297, 61.6949, 61.66652, 
    61.63783, 61.60884, 61.57955, 61.54995, 61.52005, 61.48985, 61.45935, 
    61.42855, 61.39745, 61.36605, 61.33436, 61.30238, 61.2701, 61.23752, 
    61.20465, 61.1715, 61.13805, 61.10431, 61.07029, 61.03597, 61.00137, 
    60.96649, 60.93132, 60.89587, 60.86014, 60.82413, 60.78784, 60.75127, 
    60.71442, 60.67729, 60.63989, 60.60222, 60.56427, 60.52605, 60.48756, 
    60.4488, 60.40977, 60.37047, 60.33091, 60.29108, 60.25098, 60.21062, 
    60.17001, 60.12912, 60.08798, 60.04659, 60.00492, 59.96301, 59.92084, 
    59.87841, 59.83574, 59.7928, 59.74962, 59.70619, 59.66251, 59.61858, 
    59.57441, 59.52998, 59.48532, 59.44041, 59.39526, 59.34986, 59.30423, 
    59.25836, 59.21225, 59.1659, 59.11932, 59.0725, 59.02545, 58.97816, 
    58.93065, 58.8829, 58.83493, 58.78672, 58.7383, 58.68964, 58.64076, 
    58.59166, 58.54233, 58.49278, 58.44301, 58.39302, 58.34282, 58.29239, 
    58.24175, 58.1909,
  52.75665, 52.82333, 52.88988, 52.9563, 53.02259, 53.08875, 53.15478, 
    53.22067, 53.28643, 53.35205, 53.41754, 53.48289, 53.54811, 53.61319, 
    53.67813, 53.74293, 53.80759, 53.87211, 53.93649, 54.00072, 54.06481, 
    54.12876, 54.19256, 54.25621, 54.31972, 54.38308, 54.4463, 54.50936, 
    54.57227, 54.63504, 54.69764, 54.7601, 54.82241, 54.88456, 54.94655, 
    55.00839, 55.07007, 55.13159, 55.19296, 55.25416, 55.3152, 55.37609, 
    55.43681, 55.49736, 55.55775, 55.61798, 55.67804, 55.73793, 55.79766, 
    55.85722, 55.91661, 55.97582, 56.03487, 56.09374, 56.15244, 56.21096, 
    56.26931, 56.32748, 56.38548, 56.44329, 56.50093, 56.55839, 56.61566, 
    56.67276, 56.72966, 56.78639, 56.84293, 56.89928, 56.95545, 57.01143, 
    57.06722, 57.12282, 57.17823, 57.23344, 57.28847, 57.3433, 57.39793, 
    57.45237, 57.5066, 57.56065, 57.61449, 57.66813, 57.72157, 57.7748, 
    57.82784, 57.88066, 57.93329, 57.98571, 58.03791, 58.08991, 58.1417, 
    58.19328, 58.24465, 58.2958, 58.34674, 58.39746, 58.44797, 58.49826, 
    58.54833, 58.59818, 58.64781, 58.69722, 58.74641, 58.79537, 58.84411, 
    58.89262, 58.9409, 58.98896, 59.03679, 59.08438, 59.13174, 59.17887, 
    59.22577, 59.27243, 59.31886, 59.36505, 59.411, 59.45671, 59.50218, 
    59.54741, 59.59239, 59.63713, 59.68163, 59.72588, 59.76988, 59.81364, 
    59.85714, 59.9004, 59.9434, 59.98615, 60.02865, 60.07089, 60.11288, 
    60.15461, 60.19608, 60.23729, 60.27824, 60.31892, 60.35935, 60.39951, 
    60.4394, 60.47903, 60.5184, 60.55749, 60.59632, 60.63487, 60.67315, 
    60.71116, 60.7489, 60.78636, 60.82355, 60.86045, 60.89708, 60.93344, 
    60.96951, 61.00529, 61.0408, 61.07602, 61.11096, 61.14561, 61.17998, 
    61.21406, 61.24785, 61.28135, 61.31456, 61.34747, 61.3801, 61.41243, 
    61.44446, 61.4762, 61.50764, 61.53878, 61.56963, 61.60017, 61.63042, 
    61.66036, 61.68999, 61.71933, 61.74836, 61.77708, 61.8055, 61.83361, 
    61.86141, 61.8889, 61.91608, 61.94294, 61.9695, 61.99574, 62.02167, 
    62.04728, 62.07257, 62.09756, 62.12222, 62.14656, 62.17058, 62.19429, 
    62.21767, 62.24073, 62.26346, 62.28587, 62.30796, 62.32973, 62.35116, 
    62.37227, 62.39305, 62.41351, 62.43364, 62.45343, 62.47289, 62.49203, 
    62.51083, 62.5293, 62.54743, 62.56523, 62.5827, 62.59983, 62.61662, 
    62.63308, 62.6492, 62.66499, 62.68043, 62.69553, 62.7103, 62.72472, 
    62.73881, 62.75255, 62.76596, 62.77901, 62.79173, 62.8041, 62.81613, 
    62.82782, 62.83916, 62.85015, 62.8608, 62.87111, 62.88106, 62.89067, 
    62.89994, 62.90885, 62.91742, 62.92564, 62.93351, 62.94103, 62.9482, 
    62.95503, 62.9615, 62.96762, 62.9734, 62.97882, 62.98389, 62.98861, 
    62.99298, 62.99701, 63.00067, 63.00399, 63.00695, 63.00957, 63.01183, 
    63.01374, 63.01529, 63.0165, 63.01735, 63.01785, 63.018, 63.0178, 
    63.01724, 63.01633, 63.01507, 63.01346, 63.01149, 63.00917, 63.00651, 
    63.00349, 63.00011, 62.99639, 62.99232, 62.98789, 62.98312, 62.97799, 
    62.97251, 62.96668, 62.9605, 62.95397, 62.94709, 62.93987, 62.93229, 
    62.92436, 62.91609, 62.90746, 62.89849, 62.88918, 62.87951, 62.8695, 
    62.85914, 62.84844, 62.83739, 62.82599, 62.81425, 62.80217, 62.78974, 
    62.77697, 62.76386, 62.7504, 62.73661, 62.72247, 62.70799, 62.69317, 
    62.67801, 62.66251, 62.64668, 62.6305, 62.61399, 62.59714, 62.57996, 
    62.56244, 62.54458, 62.5264, 62.50788, 62.48902, 62.46984, 62.45032, 
    62.43047, 62.4103, 62.38979, 62.36895, 62.34779, 62.32631, 62.30449, 
    62.28235, 62.25989, 62.2371, 62.21399, 62.19056, 62.16681, 62.14273, 
    62.11834, 62.09362, 62.0686, 62.04325, 62.01759, 61.99161, 61.96532, 
    61.93871, 61.9118, 61.88457, 61.85703, 61.82918, 61.80103, 61.77256, 
    61.74379, 61.71471, 61.68533, 61.65564, 61.62565, 61.59536, 61.56477, 
    61.53388, 61.50269, 61.4712, 61.43941, 61.40733, 61.37496, 61.34229, 
    61.30932, 61.27607, 61.24252, 61.20869, 61.17456, 61.14015, 61.10546, 
    61.07047, 61.03521, 60.99965, 60.96382, 60.9277, 60.89131, 60.85464, 
    60.81768, 60.78045, 60.74295, 60.70517, 60.66712, 60.62879, 60.59019, 
    60.55133, 60.51219, 60.47279, 60.43311, 60.39317, 60.35297, 60.3125, 
    60.27177, 60.23079, 60.18953, 60.14802, 60.10625, 60.06423, 60.02195, 
    59.97941, 59.93662, 59.89357, 59.85028, 59.80674, 59.76294, 59.7189, 
    59.67461, 59.63007, 59.58529, 59.54027, 59.495, 59.44949, 59.40374, 
    59.35775, 59.31153, 59.26507, 59.21837, 59.17143, 59.12427, 59.07687, 
    59.02923, 58.98137, 58.93328, 58.88496, 58.83641, 58.78764, 58.73864, 
    58.68942, 58.63998, 58.59031, 58.54042, 58.49032, 58.43999, 58.38945, 
    58.3387, 58.28772,
  52.84282, 52.9096, 52.97626, 53.04278, 53.10918, 53.17545, 53.24158, 
    53.30758, 53.37344, 53.43917, 53.50477, 53.57023, 53.63555, 53.70074, 
    53.76579, 53.8307, 53.89546, 53.96009, 54.02458, 54.08892, 54.15312, 
    54.21717, 54.28109, 54.34485, 54.40847, 54.47194, 54.53527, 54.59844, 
    54.66147, 54.72434, 54.78706, 54.84963, 54.91205, 54.97431, 55.03642, 
    55.09837, 55.16016, 55.2218, 55.28328, 55.34459, 55.40575, 55.46675, 
    55.52758, 55.58825, 55.64876, 55.7091, 55.76928, 55.82928, 55.88913, 
    55.9488, 56.0083, 56.06763, 56.1268, 56.18578, 56.2446, 56.30324, 
    56.3617, 56.41999, 56.4781, 56.53604, 56.59379, 56.65137, 56.70876, 
    56.76597, 56.823, 56.87984, 56.9365, 56.99297, 57.04926, 57.10535, 
    57.16126, 57.21698, 57.2725, 57.32784, 57.38298, 57.43793, 57.49268, 
    57.54723, 57.60159, 57.65575, 57.70971, 57.76347, 57.81703, 57.87038, 
    57.92353, 57.97648, 58.02922, 58.08176, 58.13409, 58.1862, 58.23811, 
    58.28981, 58.34129, 58.39257, 58.44362, 58.49446, 58.54509, 58.5955, 
    58.64569, 58.69566, 58.74541, 58.79493, 58.84424, 58.89332, 58.94217, 
    58.9908, 59.0392, 59.08738, 59.13532, 59.18303, 59.23051, 59.27776, 
    59.32477, 59.37155, 59.41809, 59.4644, 59.51046, 59.55629, 59.60188, 
    59.64722, 59.69232, 59.73717, 59.78179, 59.82615, 59.87027, 59.91414, 
    59.95776, 60.00113, 60.04424, 60.0871, 60.12971, 60.17207, 60.21416, 
    60.256, 60.29759, 60.33891, 60.37997, 60.42076, 60.4613, 60.50157, 
    60.54158, 60.58131, 60.62078, 60.65999, 60.69892, 60.73758, 60.77597, 
    60.81409, 60.85193, 60.8895, 60.92678, 60.9638, 61.00053, 61.03698, 
    61.07316, 61.10905, 61.14466, 61.17998, 61.21502, 61.24977, 61.28424, 
    61.31842, 61.3523, 61.3859, 61.4192, 61.45222, 61.48494, 61.51736, 
    61.54949, 61.58133, 61.61286, 61.6441, 61.67503, 61.70567, 61.736, 
    61.76603, 61.79576, 61.82518, 61.8543, 61.88311, 61.91161, 61.93981, 
    61.96769, 61.99527, 62.02253, 62.04948, 62.07612, 62.10244, 62.12845, 
    62.15414, 62.17952, 62.20457, 62.22931, 62.25373, 62.27783, 62.30161, 
    62.32506, 62.34819, 62.371, 62.39348, 62.41564, 62.43747, 62.45898, 
    62.48016, 62.501, 62.52152, 62.54171, 62.56157, 62.5811, 62.60029, 
    62.61916, 62.63768, 62.65588, 62.67374, 62.69126, 62.70845, 62.7253, 
    62.74181, 62.75798, 62.77382, 62.78931, 62.80446, 62.81928, 62.83375, 
    62.84788, 62.86167, 62.87511, 62.88822, 62.90098, 62.91339, 62.92546, 
    62.93718, 62.94856, 62.95959, 62.97028, 62.98061, 62.9906, 63.00025, 
    63.00954, 63.01849, 63.02708, 63.03533, 63.04322, 63.05077, 63.05797, 
    63.06482, 63.07131, 63.07746, 63.08325, 63.08869, 63.09378, 63.09851, 
    63.1029, 63.10693, 63.11061, 63.11394, 63.11692, 63.11954, 63.12181, 
    63.12372, 63.12528, 63.12649, 63.12735, 63.12785, 63.128, 63.12779, 
    63.12724, 63.12632, 63.12506, 63.12344, 63.12147, 63.11914, 63.11647, 
    63.11344, 63.11005, 63.10632, 63.10223, 63.09779, 63.093, 63.08785, 
    63.08236, 63.07651, 63.07031, 63.06376, 63.05685, 63.0496, 63.042, 
    63.03405, 63.02575, 63.01709, 63.00809, 62.99874, 62.98905, 62.979, 
    62.96861, 62.95787, 62.94678, 62.93535, 62.92357, 62.91145, 62.89898, 
    62.88617, 62.87301, 62.85951, 62.84567, 62.83148, 62.81696, 62.80209, 
    62.78688, 62.77133, 62.75544, 62.73922, 62.72265, 62.70575, 62.68851, 
    62.67093, 62.65302, 62.63477, 62.6162, 62.59728, 62.57803, 62.55845, 
    62.53854, 62.5183, 62.49773, 62.47683, 62.4556, 62.43404, 62.41216, 
    62.38995, 62.36741, 62.34455, 62.32137, 62.29786, 62.27404, 62.24989, 
    62.22542, 62.20063, 62.17552, 62.1501, 62.12436, 62.0983, 62.07193, 
    62.04524, 62.01824, 61.99092, 61.9633, 61.93537, 61.90713, 61.87857, 
    61.84972, 61.82055, 61.79108, 61.7613, 61.73122, 61.70084, 61.67016, 
    61.63918, 61.60789, 61.57631, 61.54443, 61.51225, 61.47978, 61.44702, 
    61.41396, 61.3806, 61.34696, 61.31303, 61.2788, 61.24429, 61.2095, 
    61.17441, 61.13904, 61.10339, 61.06746, 61.03124, 60.99474, 60.95796, 
    60.92091, 60.88357, 60.84596, 60.80807, 60.76992, 60.73148, 60.69278, 
    60.6538, 60.61456, 60.57505, 60.53527, 60.49522, 60.45491, 60.41433, 
    60.37349, 60.33239, 60.29103, 60.2494, 60.20752, 60.16539, 60.12299, 
    60.08034, 60.03744, 59.99428, 59.95087, 59.90722, 59.86331, 59.81915, 
    59.77475, 59.7301, 59.6852, 59.64006, 59.59468, 59.54906, 59.50319, 
    59.45709, 59.41075, 59.36417, 59.31735, 59.2703, 59.22301, 59.1755, 
    59.12775, 59.07977, 59.03156, 58.98312, 58.93446, 58.88557, 58.83646, 
    58.78712, 58.73755, 58.68777, 58.63776, 58.58754, 58.5371, 58.48644, 
    58.43556, 58.38447,
  52.92888, 52.99577, 53.06253, 53.12916, 53.19566, 53.26203, 53.32827, 
    53.39437, 53.46035, 53.52619, 53.59189, 53.65746, 53.72289, 53.78818, 
    53.85334, 53.91835, 53.98323, 54.04797, 54.11256, 54.17702, 54.24133, 
    54.30549, 54.36951, 54.43339, 54.49712, 54.5607, 54.62414, 54.68742, 
    54.75056, 54.81355, 54.87638, 54.93906, 55.00159, 55.06396, 55.12618, 
    55.18825, 55.25016, 55.3119, 55.3735, 55.43493, 55.4962, 55.55731, 
    55.61826, 55.67904, 55.73967, 55.80012, 55.86041, 55.92054, 55.9805, 
    56.04028, 56.0999, 56.15935, 56.21863, 56.27773, 56.33667, 56.39542, 
    56.454, 56.51241, 56.57064, 56.62869, 56.68656, 56.74425, 56.80176, 
    56.85909, 56.91624, 56.9732, 57.02998, 57.08656, 57.14297, 57.19918, 
    57.25521, 57.31105, 57.36669, 57.42214, 57.4774, 57.53247, 57.58734, 
    57.64201, 57.69649, 57.75077, 57.80485, 57.85873, 57.9124, 57.96588, 
    58.01915, 58.07222, 58.12508, 58.17773, 58.23018, 58.28242, 58.33444, 
    58.38626, 58.43786, 58.48925, 58.54043, 58.59139, 58.64214, 58.69266, 
    58.74297, 58.79306, 58.84293, 58.89257, 58.942, 58.9912, 59.04017, 
    59.08891, 59.13743, 59.18572, 59.23378, 59.28161, 59.32921, 59.37658, 
    59.42371, 59.4706, 59.51726, 59.56368, 59.60986, 59.65581, 59.70151, 
    59.74697, 59.79219, 59.83716, 59.88189, 59.92636, 59.9706, 60.01458, 
    60.05831, 60.1018, 60.14502, 60.188, 60.23072, 60.27319, 60.3154, 
    60.35735, 60.39904, 60.44048, 60.48165, 60.52256, 60.5632, 60.60358, 
    60.6437, 60.68354, 60.72312, 60.76243, 60.80147, 60.84024, 60.87874, 
    60.91696, 60.95491, 60.99258, 61.02998, 61.06709, 61.10393, 61.14049, 
    61.17677, 61.21276, 61.24847, 61.2839, 61.31903, 61.35389, 61.38845, 
    61.42273, 61.45672, 61.49041, 61.52382, 61.55693, 61.58974, 61.62226, 
    61.65449, 61.68642, 61.71804, 61.74937, 61.7804, 61.81113, 61.84156, 
    61.87168, 61.9015, 61.93101, 61.96022, 61.98911, 62.0177, 62.04598, 
    62.07395, 62.10161, 62.12896, 62.15599, 62.18271, 62.20912, 62.23521, 
    62.26098, 62.28643, 62.31157, 62.33638, 62.36088, 62.38505, 62.40891, 
    62.43243, 62.45564, 62.47852, 62.50108, 62.5233, 62.5452, 62.56678, 
    62.58802, 62.60894, 62.62952, 62.64978, 62.6697, 62.68929, 62.70855, 
    62.72747, 62.74606, 62.76431, 62.78223, 62.79981, 62.81705, 62.83395, 
    62.85052, 62.86675, 62.88263, 62.89818, 62.91338, 62.92825, 62.94277, 
    62.95695, 62.97078, 62.98427, 62.99741, 63.01022, 63.02267, 63.03478, 
    63.04654, 63.05796, 63.06903, 63.07975, 63.09012, 63.10014, 63.10982, 
    63.11914, 63.12812, 63.13674, 63.14502, 63.15294, 63.16051, 63.16773, 
    63.1746, 63.18112, 63.18729, 63.1931, 63.19855, 63.20366, 63.20842, 
    63.21282, 63.21686, 63.22055, 63.22389, 63.22688, 63.22951, 63.23178, 
    63.23371, 63.23528, 63.23649, 63.23735, 63.23785, 63.238, 63.23779, 
    63.23723, 63.23632, 63.23505, 63.23343, 63.23145, 63.22911, 63.22643, 
    63.22339, 63.21999, 63.21625, 63.21214, 63.20769, 63.20288, 63.19772, 
    63.1922, 63.18633, 63.18011, 63.17354, 63.16661, 63.15934, 63.15171, 
    63.14373, 63.1354, 63.12672, 63.11769, 63.10831, 63.09858, 63.0885, 
    63.07808, 63.0673, 63.05618, 63.0447, 63.03289, 63.02073, 63.00821, 
    62.99536, 62.98216, 62.96861, 62.95473, 62.94049, 62.92592, 62.911, 
    62.89574, 62.88014, 62.8642, 62.84792, 62.8313, 62.81435, 62.79705, 
    62.77942, 62.76145, 62.74314, 62.7245, 62.70552, 62.68621, 62.66657, 
    62.6466, 62.62629, 62.60565, 62.58469, 62.56339, 62.54176, 62.51981, 
    62.49753, 62.47492, 62.45199, 62.42873, 62.40515, 62.38125, 62.35703, 
    62.33248, 62.30761, 62.28242, 62.25692, 62.2311, 62.20496, 62.1785, 
    62.15174, 62.12465, 62.09726, 62.06955, 62.04153, 62.0132, 61.98456, 
    61.95562, 61.92636, 61.8968, 61.86694, 61.83677, 61.80629, 61.77552, 
    61.74444, 61.71306, 61.68139, 61.64941, 61.61714, 61.58457, 61.55171, 
    61.51855, 61.4851, 61.45136, 61.41733, 61.38301, 61.3484, 61.3135, 
    61.27831, 61.24284, 61.20708, 61.17105, 61.13472, 61.09812, 61.06124, 
    61.02408, 60.98664, 60.94893, 60.91093, 60.87267, 60.83413, 60.79531, 
    60.75623, 60.71688, 60.67726, 60.63737, 60.59721, 60.55679, 60.5161, 
    60.47515, 60.43394, 60.39246, 60.35073, 60.30874, 60.26649, 60.22398, 
    60.18122, 60.1382, 60.09493, 60.05141, 60.00764, 59.96362, 59.91935, 
    59.87482, 59.83006, 59.78505, 59.7398, 59.6943, 59.64856, 59.60258, 
    59.55635, 59.5099, 59.4632, 59.41627, 59.3691, 59.3217, 59.27406, 
    59.2262, 59.1781, 59.12977, 59.08122, 59.03244, 58.98343, 58.93419, 
    58.88474, 58.83505, 58.78515, 58.73503, 58.68468, 58.63412, 58.58334, 
    58.53235, 58.48114,
  53.01483, 53.08183, 53.14869, 53.21543, 53.28204, 53.34851, 53.41486, 
    53.48107, 53.54715, 53.61309, 53.6789, 53.74458, 53.81012, 53.87552, 
    53.94078, 54.00591, 54.07089, 54.13574, 54.20044, 54.26501, 54.32943, 
    54.3937, 54.45784, 54.52182, 54.58566, 54.64936, 54.7129, 54.7763, 
    54.83955, 54.90265, 54.96559, 55.02839, 55.09103, 55.15351, 55.21585, 
    55.27803, 55.34005, 55.40191, 55.46362, 55.52516, 55.58655, 55.64777, 
    55.70884, 55.76974, 55.83047, 55.89105, 55.95145, 56.0117, 56.07177, 
    56.13167, 56.19141, 56.25097, 56.31036, 56.36959, 56.42863, 56.48751, 
    56.54621, 56.60473, 56.66308, 56.72125, 56.77924, 56.83705, 56.89468, 
    56.95212, 57.00938, 57.06646, 57.12336, 57.18007, 57.23659, 57.29293, 
    57.34907, 57.40503, 57.46079, 57.51636, 57.57174, 57.62693, 57.68192, 
    57.73671, 57.79131, 57.8457, 57.8999, 57.9539, 58.0077, 58.06129, 
    58.11468, 58.16787, 58.22085, 58.27362, 58.32619, 58.37855, 58.43069, 
    58.48263, 58.53435, 58.58586, 58.63716, 58.68824, 58.73911, 58.78975, 
    58.84018, 58.89038, 58.94037, 58.99014, 59.03968, 59.089, 59.13809, 
    59.18695, 59.23559, 59.284, 59.33218, 59.38013, 59.42784, 59.47533, 
    59.52258, 59.56959, 59.61636, 59.6629, 59.7092, 59.75526, 59.80108, 
    59.84665, 59.89199, 59.93708, 59.98192, 60.02651, 60.07086, 60.11496, 
    60.15881, 60.2024, 60.24575, 60.28884, 60.33167, 60.37425, 60.41658, 
    60.45864, 60.50044, 60.54199, 60.58327, 60.62429, 60.66505, 60.70554, 
    60.74576, 60.78572, 60.82541, 60.86483, 60.90398, 60.94286, 60.98146, 
    61.01979, 61.05784, 61.09562, 61.13312, 61.17035, 61.20729, 61.24395, 
    61.28033, 61.31643, 61.35224, 61.38777, 61.42301, 61.45797, 61.49263, 
    61.52701, 61.5611, 61.59489, 61.62839, 61.6616, 61.69452, 61.72713, 
    61.75945, 61.79147, 61.8232, 61.85462, 61.88574, 61.91656, 61.94708, 
    61.97729, 62.0072, 62.0368, 62.0661, 62.09509, 62.12376, 62.15213, 
    62.18019, 62.20793, 62.23536, 62.26248, 62.28928, 62.31577, 62.34194, 
    62.36779, 62.39333, 62.41854, 62.44344, 62.46801, 62.49226, 62.51619, 
    62.53979, 62.56307, 62.58602, 62.60865, 62.63095, 62.65292, 62.67456, 
    62.69588, 62.71686, 62.73751, 62.75783, 62.77782, 62.79747, 62.81679, 
    62.83577, 62.85442, 62.87273, 62.89071, 62.90835, 62.92565, 62.94261, 
    62.95923, 62.97551, 62.99144, 63.00704, 63.0223, 63.03721, 63.05178, 
    63.066, 63.07988, 63.09342, 63.10661, 63.11945, 63.13195, 63.1441, 
    63.1559, 63.16735, 63.17846, 63.18921, 63.19962, 63.20968, 63.21938, 
    63.22874, 63.23775, 63.2464, 63.2547, 63.26265, 63.27025, 63.2775, 
    63.28439, 63.29093, 63.29711, 63.30294, 63.30842, 63.31355, 63.31832, 
    63.32273, 63.32679, 63.3305, 63.33385, 63.33684, 63.33948, 63.34176, 
    63.34369, 63.34526, 63.34648, 63.34734, 63.34785, 63.348, 63.34779, 
    63.34723, 63.34631, 63.34504, 63.34341, 63.34143, 63.33908, 63.33639, 
    63.33334, 63.32993, 63.32617, 63.32206, 63.31758, 63.31276, 63.30758, 
    63.30205, 63.29616, 63.28992, 63.28332, 63.27637, 63.26907, 63.26142, 
    63.25341, 63.24506, 63.23634, 63.22728, 63.21787, 63.20811, 63.198, 
    63.18753, 63.17672, 63.16556, 63.15405, 63.1422, 63.12999, 63.11744, 
    63.10455, 63.0913, 63.07771, 63.06377, 63.0495, 63.03487, 63.01991, 
    63.0046, 62.98895, 62.97295, 62.95662, 62.93995, 62.92293, 62.90558, 
    62.88789, 62.86986, 62.8515, 62.83279, 62.81376, 62.79438, 62.77468, 
    62.75464, 62.73427, 62.71356, 62.69253, 62.67116, 62.64947, 62.62744, 
    62.60509, 62.58241, 62.55941, 62.53608, 62.51242, 62.48844, 62.46414, 
    62.43952, 62.41457, 62.38931, 62.36372, 62.33782, 62.3116, 62.28506, 
    62.25821, 62.23104, 62.20356, 62.17577, 62.14766, 62.11925, 62.09052, 
    62.06149, 62.03214, 62.00249, 61.97253, 61.94228, 61.91171, 61.88084, 
    61.84967, 61.8182, 61.78643, 61.75436, 61.72199, 61.68933, 61.65637, 
    61.62311, 61.58957, 61.55572, 61.52159, 61.48717, 61.45246, 61.41746, 
    61.38217, 61.3466, 61.31074, 61.27459, 61.23817, 61.20146, 61.16447, 
    61.12721, 61.08966, 61.05184, 61.01374, 60.97537, 60.93672, 60.8978, 
    60.85861, 60.81915, 60.77942, 60.73942, 60.69915, 60.65862, 60.61782, 
    60.57676, 60.53543, 60.49385, 60.452, 60.4099, 60.36753, 60.32491, 
    60.28204, 60.23891, 60.19552, 60.15189, 60.108, 60.06386, 60.01947, 
    59.97484, 59.92996, 59.88483, 59.83946, 59.79385, 59.74799, 59.70189, 
    59.65556, 59.60898, 59.56216, 59.51511, 59.46783, 59.42031, 59.37256, 
    59.32457, 59.27636, 59.22791, 59.17924, 59.13034, 59.08121, 59.03186, 
    58.98228, 58.93248, 58.88246, 58.83221, 58.78175, 58.73107, 58.68018, 
    58.62906, 58.57773,
  53.10067, 53.16777, 53.23475, 53.30159, 53.3683, 53.43488, 53.50133, 
    53.56765, 53.63384, 53.69989, 53.76581, 53.83159, 53.89724, 53.96275, 
    54.02812, 54.09336, 54.15845, 54.2234, 54.28822, 54.35289, 54.41742, 
    54.48181, 54.54605, 54.61015, 54.6741, 54.73791, 54.80156, 54.86507, 
    54.92843, 54.99164, 55.0547, 55.11761, 55.18036, 55.24297, 55.30541, 
    55.3677, 55.42984, 55.49181, 55.55363, 55.6153, 55.6768, 55.73814, 
    55.79932, 55.86033, 55.92118, 55.98187, 56.0424, 56.10275, 56.16294, 
    56.22296, 56.28281, 56.34249, 56.40201, 56.46135, 56.52051, 56.5795, 
    56.63832, 56.69696, 56.75542, 56.81371, 56.87182, 56.92975, 56.9875, 
    57.04506, 57.10244, 57.15964, 57.21666, 57.27348, 57.33012, 57.38658, 
    57.44284, 57.49892, 57.5548, 57.61049, 57.66599, 57.72129, 57.77641, 
    57.83132, 57.88603, 57.94055, 57.99487, 58.04899, 58.10291, 58.15662, 
    58.21013, 58.26344, 58.31654, 58.36943, 58.42212, 58.47459, 58.52686, 
    58.57892, 58.63076, 58.68239, 58.73381, 58.78501, 58.83599, 58.88676, 
    58.93731, 58.98764, 59.03774, 59.08763, 59.13729, 59.18672, 59.23594, 
    59.28492, 59.33368, 59.3822, 59.4305, 59.47857, 59.5264, 59.57401, 
    59.62137, 59.6685, 59.7154, 59.76205, 59.80847, 59.85464, 59.90058, 
    59.94627, 59.99172, 60.03693, 60.08189, 60.1266, 60.17106, 60.21527, 
    60.25924, 60.30295, 60.34641, 60.38961, 60.43256, 60.47526, 60.51769, 
    60.55987, 60.60179, 60.64344, 60.68484, 60.72597, 60.76684, 60.80744, 
    60.84778, 60.88784, 60.92764, 60.96717, 61.00643, 61.04542, 61.08413, 
    61.12257, 61.16073, 61.19862, 61.23622, 61.27355, 61.3106, 61.34737, 
    61.38385, 61.42005, 61.45597, 61.4916, 61.52695, 61.562, 61.59677, 
    61.63125, 61.66543, 61.69933, 61.73293, 61.76624, 61.79925, 61.83196, 
    61.86438, 61.8965, 61.92831, 61.95984, 61.99105, 62.02197, 62.05257, 
    62.08288, 62.11288, 62.14257, 62.17196, 62.20103, 62.22979, 62.25825, 
    62.28639, 62.31422, 62.34174, 62.36894, 62.39583, 62.4224, 62.44865, 
    62.47458, 62.5002, 62.52549, 62.55046, 62.57512, 62.59944, 62.62345, 
    62.64713, 62.67048, 62.6935, 62.71621, 62.73857, 62.76062, 62.78233, 
    62.80371, 62.82476, 62.84548, 62.86587, 62.88592, 62.90564, 62.92502, 
    62.94407, 62.96278, 62.98115, 62.99918, 63.01688, 63.03423, 63.05125, 
    63.06792, 63.08426, 63.10025, 63.1159, 63.1312, 63.14616, 63.16078, 
    63.17505, 63.18898, 63.20256, 63.21579, 63.22868, 63.24122, 63.25341, 
    63.26525, 63.27674, 63.28788, 63.29868, 63.30912, 63.31921, 63.32895, 
    63.33834, 63.34737, 63.35606, 63.36439, 63.37236, 63.37999, 63.38726, 
    63.39417, 63.40073, 63.40694, 63.41279, 63.41829, 63.42343, 63.42822, 
    63.43264, 63.43672, 63.44044, 63.4438, 63.4468, 63.44945, 63.45174, 
    63.45368, 63.45526, 63.45648, 63.45734, 63.45785, 63.458, 63.45779, 
    63.45723, 63.45631, 63.45503, 63.4534, 63.4514, 63.44905, 63.44635, 
    63.44329, 63.43987, 63.4361, 63.43197, 63.42748, 63.42264, 63.41744, 
    63.41189, 63.40598, 63.39972, 63.3931, 63.38613, 63.3788, 63.37112, 
    63.36309, 63.35471, 63.34597, 63.33688, 63.32743, 63.31763, 63.30749, 
    63.29699, 63.28614, 63.27495, 63.2634, 63.2515, 63.23926, 63.22666, 
    63.21372, 63.20044, 63.1868, 63.17282, 63.15849, 63.14382, 63.1288, 
    63.11345, 63.09774, 63.0817, 63.06531, 63.04858, 63.03151, 63.0141, 
    62.99635, 62.97826, 62.95984, 62.94107, 62.92197, 62.90254, 62.88277, 
    62.86267, 62.84223, 62.82146, 62.80035, 62.77892, 62.75715, 62.73506, 
    62.71264, 62.68988, 62.66681, 62.6434, 62.61967, 62.59562, 62.57124, 
    62.54654, 62.52151, 62.49617, 62.4705, 62.44452, 62.41822, 62.3916, 
    62.36466, 62.33741, 62.30984, 62.28196, 62.25377, 62.22527, 62.19645, 
    62.16733, 62.13789, 62.10815, 62.07811, 62.04775, 62.01709, 61.98613, 
    61.95487, 61.9233, 61.89144, 61.85927, 61.82681, 61.79404, 61.76099, 
    61.72763, 61.69398, 61.66005, 61.62581, 61.59129, 61.55648, 61.52137, 
    61.48598, 61.45031, 61.41434, 61.3781, 61.34157, 61.30476, 61.26767, 
    61.23029, 61.19264, 61.15471, 61.1165, 61.07803, 61.03927, 61.00024, 
    60.96094, 60.92137, 60.88153, 60.84142, 60.80104, 60.76039, 60.71948, 
    60.67831, 60.63688, 60.59518, 60.55322, 60.511, 60.46852, 60.42579, 
    60.3828, 60.33955, 60.29605, 60.2523, 60.2083, 60.16404, 60.11954, 
    60.07479, 60.02979, 59.98455, 59.93906, 59.89333, 59.84736, 59.80114, 
    59.75469, 59.70799, 59.66106, 59.6139, 59.56649, 59.51885, 59.47098, 
    59.42288, 59.37454, 59.32598, 59.27719, 59.22816, 59.17892, 59.12945, 
    59.07975, 59.02983, 58.97969, 58.92933, 58.87875, 58.82794, 58.77692, 
    58.72569, 58.67424,
  53.18641, 53.25361, 53.32069, 53.38764, 53.45446, 53.52114, 53.5877, 
    53.65413, 53.72042, 53.78658, 53.8526, 53.9185, 53.98425, 54.04987, 
    54.11535, 54.18069, 54.2459, 54.31096, 54.37589, 54.44067, 54.50531, 
    54.56981, 54.63416, 54.69837, 54.76243, 54.82635, 54.89012, 54.95374, 
    55.01722, 55.08054, 55.14371, 55.20673, 55.2696, 55.33231, 55.39487, 
    55.45728, 55.51953, 55.58162, 55.64355, 55.70533, 55.76694, 55.8284, 
    55.88969, 55.95082, 56.0118, 56.0726, 56.13324, 56.19371, 56.25402, 
    56.31415, 56.37412, 56.43392, 56.49355, 56.55301, 56.61229, 56.6714, 
    56.73034, 56.78909, 56.84768, 56.90608, 56.96431, 57.02235, 57.08022, 
    57.13791, 57.1954, 57.25272, 57.30986, 57.3668, 57.42356, 57.48014, 
    57.53652, 57.59272, 57.64872, 57.70453, 57.76015, 57.81557, 57.8708, 
    57.92584, 57.98067, 58.03531, 58.08975, 58.14399, 58.19803, 58.25187, 
    58.3055, 58.35892, 58.41214, 58.46516, 58.51797, 58.57056, 58.62295, 
    58.67513, 58.72709, 58.77884, 58.83038, 58.8817, 58.9328, 58.98369, 
    59.03436, 59.08481, 59.13503, 59.18504, 59.23482, 59.28438, 59.33371, 
    59.38281, 59.43169, 59.48034, 59.52875, 59.57694, 59.62489, 59.67261, 
    59.7201, 59.76735, 59.81436, 59.86113, 59.90767, 59.95396, 60.00002, 
    60.04583, 60.0914, 60.13672, 60.18179, 60.22662, 60.2712, 60.31553, 
    60.35961, 60.40344, 60.44701, 60.49033, 60.53339, 60.5762, 60.61876, 
    60.66105, 60.70308, 60.74485, 60.78635, 60.8276, 60.86858, 60.90929, 
    60.94974, 60.98992, 61.02983, 61.06947, 61.10883, 61.14793, 61.18675, 
    61.2253, 61.26357, 61.30156, 61.33928, 61.37671, 61.41386, 61.45074, 
    61.48733, 61.52364, 61.55965, 61.59539, 61.63084, 61.666, 61.70087, 
    61.73544, 61.76973, 61.80373, 61.83743, 61.87083, 61.90394, 61.93676, 
    61.96927, 62.00148, 62.0334, 62.06501, 62.09632, 62.12733, 62.15803, 
    62.18843, 62.21852, 62.24831, 62.27778, 62.30695, 62.3358, 62.36434, 
    62.39257, 62.42049, 62.44809, 62.47538, 62.50235, 62.529, 62.55534, 
    62.58135, 62.60705, 62.63242, 62.65747, 62.6822, 62.7066, 62.73069, 
    62.75444, 62.77787, 62.80097, 62.82374, 62.84618, 62.8683, 62.89008, 
    62.91153, 62.93265, 62.95344, 62.97389, 62.99401, 63.01379, 63.03323, 
    63.05234, 63.07111, 63.08955, 63.10764, 63.12539, 63.14281, 63.15988, 
    63.17661, 63.193, 63.20904, 63.22474, 63.2401, 63.25511, 63.26978, 
    63.2841, 63.29807, 63.3117, 63.32497, 63.3379, 63.35048, 63.36271, 
    63.3746, 63.38612, 63.3973, 63.40813, 63.41861, 63.42874, 63.43851, 
    63.44793, 63.457, 63.46571, 63.47407, 63.48207, 63.48972, 63.49702, 
    63.50396, 63.51054, 63.51677, 63.52264, 63.52815, 63.53331, 63.53811, 
    63.54256, 63.54665, 63.55038, 63.55375, 63.55676, 63.55942, 63.56172, 
    63.56366, 63.56525, 63.56647, 63.56734, 63.56785, 63.568, 63.56779, 
    63.56723, 63.5663, 63.56502, 63.56338, 63.56138, 63.55902, 63.55631, 
    63.55324, 63.54981, 63.54602, 63.54188, 63.53738, 63.53252, 63.52731, 
    63.52173, 63.5158, 63.50952, 63.50288, 63.49588, 63.48853, 63.48083, 
    63.47277, 63.46435, 63.45559, 63.44646, 63.43699, 63.42716, 63.41698, 
    63.40644, 63.39556, 63.38432, 63.37274, 63.3608, 63.34851, 63.33588, 
    63.3229, 63.30956, 63.29588, 63.28185, 63.26748, 63.25276, 63.23769, 
    63.22228, 63.20653, 63.19043, 63.17398, 63.1572, 63.14008, 63.12261, 
    63.1048, 63.08665, 63.06817, 63.04934, 63.03018, 63.01068, 62.99085, 
    62.97068, 62.95017, 62.92933, 62.90816, 62.88666, 62.86482, 62.84266, 
    62.82016, 62.79734, 62.77419, 62.75071, 62.7269, 62.70277, 62.67831, 
    62.65353, 62.62843, 62.603, 62.57726, 62.55119, 62.52481, 62.4981, 
    62.47108, 62.44374, 62.4161, 62.38813, 62.35985, 62.33126, 62.30235, 
    62.27314, 62.24361, 62.21378, 62.18364, 62.1532, 62.12244, 62.09139, 
    62.06003, 62.02837, 61.99641, 61.96415, 61.93158, 61.89872, 61.86557, 
    61.83212, 61.79837, 61.76433, 61.73, 61.69537, 61.66045, 61.62525, 
    61.58976, 61.55398, 61.51791, 61.48156, 61.44492, 61.408, 61.37081, 
    61.33333, 61.29557, 61.25753, 61.21922, 61.18063, 61.14177, 61.10263, 
    61.06321, 61.02353, 60.98358, 60.94336, 60.90287, 60.86211, 60.82109, 
    60.77981, 60.73826, 60.69645, 60.65437, 60.61204, 60.56945, 60.5266, 
    60.48349, 60.44014, 60.39652, 60.35265, 60.30854, 60.26416, 60.21955, 
    60.17468, 60.12957, 60.08421, 60.0386, 59.99275, 59.94666, 59.90033, 
    59.85375, 59.80694, 59.75989, 59.7126, 59.66508, 59.61732, 59.56933, 
    59.52111, 59.47266, 59.42397, 59.37506, 59.32592, 59.27655, 59.22696, 
    59.17714, 59.12711, 59.07684, 59.02636, 58.97566, 58.92474, 58.8736, 
    58.82224, 58.77067,
  53.27203, 53.33934, 53.40652, 53.47358, 53.5405, 53.6073, 53.67396, 
    53.74049, 53.80689, 53.87316, 53.93929, 54.00529, 54.07116, 54.13688, 
    54.20247, 54.26793, 54.33324, 54.39841, 54.46345, 54.52834, 54.59309, 
    54.6577, 54.72216, 54.78648, 54.85066, 54.91469, 54.97857, 55.0423, 
    55.10589, 55.16932, 55.23261, 55.29574, 55.35873, 55.42155, 55.48423, 
    55.54675, 55.60911, 55.67132, 55.73337, 55.79526, 55.85699, 55.91856, 
    55.97997, 56.04122, 56.1023, 56.16322, 56.22398, 56.28457, 56.34499, 
    56.40525, 56.46533, 56.52525, 56.585, 56.64457, 56.70397, 56.7632, 
    56.82225, 56.88113, 56.93983, 56.99835, 57.0567, 57.11486, 57.17285, 
    57.23065, 57.28827, 57.34571, 57.40297, 57.46003, 57.51691, 57.5736, 
    57.63011, 57.68642, 57.74255, 57.79848, 57.85422, 57.90977, 57.96512, 
    58.02027, 58.07523, 58.12999, 58.18455, 58.23891, 58.29307, 58.34702, 
    58.40078, 58.45432, 58.50767, 58.5608, 58.61373, 58.66645, 58.71896, 
    58.77126, 58.82334, 58.87521, 58.92687, 58.97831, 59.02954, 59.08054, 
    59.13133, 59.1819, 59.23225, 59.28238, 59.33228, 59.38195, 59.4314, 
    59.48063, 59.52962, 59.5784, 59.62693, 59.67524, 59.72331, 59.77115, 
    59.81876, 59.86612, 59.91326, 59.96015, 60.0068, 60.05322, 60.09939, 
    60.14532, 60.191, 60.23644, 60.28164, 60.32658, 60.37128, 60.41572, 
    60.45992, 60.50386, 60.54755, 60.59099, 60.63417, 60.67709, 60.71976, 
    60.76216, 60.80431, 60.84619, 60.88781, 60.92917, 60.97026, 61.01109, 
    61.05165, 61.09194, 61.13196, 61.17171, 61.21119, 61.25039, 61.28932, 
    61.32798, 61.36636, 61.40446, 61.44228, 61.47982, 61.51709, 61.55406, 
    61.59076, 61.62717, 61.6633, 61.69913, 61.73469, 61.76995, 61.80492, 
    61.8396, 61.87399, 61.90808, 61.94189, 61.97539, 62.0086, 62.04151, 
    62.07412, 62.10643, 62.13845, 62.17015, 62.20156, 62.23266, 62.26346, 
    62.29395, 62.32413, 62.35401, 62.38358, 62.41283, 62.44177, 62.47041, 
    62.49872, 62.52673, 62.55442, 62.58179, 62.60884, 62.63558, 62.662, 
    62.6881, 62.71387, 62.73933, 62.76446, 62.78926, 62.81375, 62.83791, 
    62.86174, 62.88524, 62.90842, 62.93126, 62.95378, 62.97596, 62.99782, 
    63.01934, 63.04052, 63.06138, 63.0819, 63.10208, 63.12193, 63.14144, 
    63.16061, 63.17944, 63.19793, 63.21609, 63.2339, 63.25137, 63.2685, 
    63.28529, 63.30173, 63.31783, 63.33358, 63.34899, 63.36405, 63.37876, 
    63.39313, 63.40715, 63.42082, 63.43414, 63.44712, 63.45974, 63.47201, 
    63.48394, 63.49551, 63.50672, 63.51759, 63.5281, 63.53826, 63.54807, 
    63.55752, 63.56662, 63.57536, 63.58374, 63.59178, 63.59945, 63.60677, 
    63.61374, 63.62034, 63.62659, 63.63248, 63.63802, 63.64319, 63.64801, 
    63.65247, 63.65657, 63.66032, 63.6637, 63.66673, 63.66939, 63.6717, 
    63.67365, 63.67524, 63.67647, 63.67734, 63.67785, 63.678, 63.67779, 
    63.67722, 63.6763, 63.67501, 63.67336, 63.67136, 63.66899, 63.66627, 
    63.66319, 63.65975, 63.65595, 63.65179, 63.64727, 63.6424, 63.63717, 
    63.63157, 63.62563, 63.61932, 63.61266, 63.60564, 63.59826, 63.59053, 
    63.58244, 63.574, 63.5652, 63.55605, 63.54654, 63.53668, 63.52646, 
    63.51589, 63.50497, 63.4937, 63.48207, 63.4701, 63.45777, 63.44509, 
    63.43206, 63.41868, 63.40496, 63.39088, 63.37646, 63.36169, 63.34657, 
    63.33111, 63.3153, 63.29915, 63.28265, 63.26581, 63.24863, 63.23111, 
    63.21324, 63.19503, 63.17648, 63.1576, 63.13837, 63.11881, 63.09891, 
    63.07867, 63.0581, 63.0372, 63.01596, 62.99438, 62.97248, 62.95024, 
    62.92767, 62.90477, 62.88155, 62.85799, 62.83411, 62.8099, 62.78536, 
    62.76051, 62.73532, 62.70982, 62.68399, 62.65784, 62.63137, 62.60458, 
    62.57748, 62.55006, 62.52232, 62.49427, 62.4659, 62.43722, 62.40822, 
    62.37892, 62.3493, 62.31938, 62.28915, 62.25861, 62.22776, 62.19661, 
    62.16516, 62.1334, 62.10135, 62.06898, 62.03632, 62.00337, 61.97011, 
    61.93656, 61.90271, 61.86857, 61.83414, 61.79941, 61.76439, 61.72908, 
    61.69349, 61.6576, 61.62143, 61.58497, 61.54823, 61.51121, 61.4739, 
    61.43632, 61.39845, 61.36031, 61.32188, 61.28318, 61.24421, 61.20496, 
    61.16544, 61.12564, 61.08558, 61.04525, 61.00465, 60.96378, 60.92265, 
    60.88124, 60.83958, 60.79766, 60.75547, 60.71302, 60.67032, 60.62735, 
    60.58413, 60.54066, 60.49693, 60.45295, 60.40871, 60.36422, 60.31948, 
    60.2745, 60.22927, 60.18379, 60.13807, 60.0921, 60.04589, 59.99944, 
    59.95275, 59.90582, 59.85865, 59.81124, 59.7636, 59.71572, 59.66761, 
    59.61927, 59.57069, 59.52189, 59.47286, 59.4236, 59.37411, 59.3244, 
    59.27446, 59.2243, 59.17392, 59.12331, 59.07249, 59.02145, 58.97019, 
    58.91871, 58.86702,
  53.35754, 53.42495, 53.49224, 53.5594, 53.62643, 53.69334, 53.76011, 
    53.82675, 53.89325, 53.95963, 54.02587, 54.09198, 54.15795, 54.22379, 
    54.28949, 54.35505, 54.42047, 54.48576, 54.5509, 54.6159, 54.68077, 
    54.74548, 54.81006, 54.87449, 54.93878, 55.00292, 55.06691, 55.13076, 
    55.19446, 55.25801, 55.3214, 55.38465, 55.44775, 55.51069, 55.57348, 
    55.63611, 55.69859, 55.76091, 55.82308, 55.88508, 55.94693, 56.00862, 
    56.07014, 56.13151, 56.19271, 56.25375, 56.31462, 56.37532, 56.43587, 
    56.49624, 56.55644, 56.61648, 56.67634, 56.73603, 56.79555, 56.8549, 
    56.91407, 56.97307, 57.03189, 57.09053, 57.14899, 57.20728, 57.26538, 
    57.32331, 57.38105, 57.43861, 57.49598, 57.55317, 57.61017, 57.66698, 
    57.72361, 57.78004, 57.83629, 57.89234, 57.9482, 58.00387, 58.05934, 
    58.11461, 58.16969, 58.22458, 58.27925, 58.33374, 58.38802, 58.44209, 
    58.49597, 58.54964, 58.6031, 58.65636, 58.70941, 58.76225, 58.81488, 
    58.8673, 58.91951, 58.9715, 59.02328, 59.07484, 59.12619, 59.17732, 
    59.22823, 59.27892, 59.32939, 59.37963, 59.42966, 59.47945, 59.52903, 
    59.57837, 59.62749, 59.67638, 59.72504, 59.77346, 59.82166, 59.86962, 
    59.91734, 59.96483, 60.01208, 60.05909, 60.10587, 60.1524, 60.19869, 
    60.24474, 60.29054, 60.3361, 60.38141, 60.42647, 60.47129, 60.51585, 
    60.56017, 60.60423, 60.64803, 60.69158, 60.73488, 60.77792, 60.8207, 
    60.86322, 60.90548, 60.94748, 60.98921, 61.03069, 61.07189, 61.11283, 
    61.1535, 61.1939, 61.23404, 61.2739, 61.31349, 61.3528, 61.39185, 
    61.43061, 61.4691, 61.50731, 61.54524, 61.58289, 61.62026, 61.65734, 
    61.69415, 61.73066, 61.7669, 61.80284, 61.83849, 61.87386, 61.90894, 
    61.94372, 61.97821, 62.01241, 62.04631, 62.07991, 62.11322, 62.14623, 
    62.17894, 62.21135, 62.24346, 62.27526, 62.30677, 62.33796, 62.36885, 
    62.39944, 62.42971, 62.45968, 62.48934, 62.51868, 62.54772, 62.57644, 
    62.60485, 62.63294, 62.66071, 62.68817, 62.71531, 62.74213, 62.76863, 
    62.79482, 62.82067, 62.84621, 62.87142, 62.89631, 62.92087, 62.94511, 
    62.96901, 62.99259, 63.01584, 63.03876, 63.06135, 63.08361, 63.10553, 
    63.12712, 63.14838, 63.1693, 63.18989, 63.21014, 63.23005, 63.24963, 
    63.26886, 63.28775, 63.30631, 63.32452, 63.3424, 63.35992, 63.37711, 
    63.39395, 63.41045, 63.4266, 63.44241, 63.45787, 63.47298, 63.48774, 
    63.50216, 63.51622, 63.52994, 63.54331, 63.55633, 63.56899, 63.58131, 
    63.59327, 63.60488, 63.61613, 63.62704, 63.63759, 63.64778, 63.65762, 
    63.6671, 63.67623, 63.68501, 63.69342, 63.70148, 63.70918, 63.71653, 
    63.72351, 63.73014, 63.73641, 63.74232, 63.74788, 63.75307, 63.75791, 
    63.76238, 63.7665, 63.77026, 63.77365, 63.77669, 63.77936, 63.78168, 
    63.78363, 63.78523, 63.78646, 63.78733, 63.78785, 63.788, 63.78779, 
    63.78722, 63.78629, 63.785, 63.78335, 63.78133, 63.77896, 63.77623, 
    63.77314, 63.76968, 63.76587, 63.7617, 63.75717, 63.75227, 63.74702, 
    63.74141, 63.73544, 63.72912, 63.72243, 63.71539, 63.70799, 63.70023, 
    63.69211, 63.68364, 63.67481, 63.66563, 63.65609, 63.64619, 63.63594, 
    63.62534, 63.61438, 63.60307, 63.5914, 63.57938, 63.56701, 63.55429, 
    63.54122, 63.5278, 63.51402, 63.4999, 63.48543, 63.47061, 63.45544, 
    63.43993, 63.42407, 63.40786, 63.39131, 63.37441, 63.35717, 63.33959, 
    63.32167, 63.3034, 63.28479, 63.26584, 63.24655, 63.22692, 63.20696, 
    63.18666, 63.16602, 63.14504, 63.12373, 63.10209, 63.08011, 63.0578, 
    63.03516, 63.01219, 62.98888, 62.96525, 62.9413, 62.91701, 62.8924, 
    62.86745, 62.84219, 62.8166, 62.7907, 62.76447, 62.73791, 62.71104, 
    62.68385, 62.65634, 62.62852, 62.60038, 62.57192, 62.54315, 62.51406, 
    62.48467, 62.45496, 62.42495, 62.39462, 62.36399, 62.33305, 62.3018, 
    62.27026, 62.2384, 62.20625, 62.17379, 62.14103, 62.10797, 62.07462, 
    62.04097, 62.00702, 61.97277, 61.93824, 61.9034, 61.86829, 61.83287, 
    61.79717, 61.76118, 61.72491, 61.68834, 61.6515, 61.61436, 61.57695, 
    61.53926, 61.50128, 61.46303, 61.4245, 61.38568, 61.3466, 61.30724, 
    61.26761, 61.22771, 61.18753, 61.14709, 61.10637, 61.06539, 61.02414, 
    60.98263, 60.94085, 60.89881, 60.85651, 60.81395, 60.77113, 60.72805, 
    60.68471, 60.64112, 60.59727, 60.55317, 60.50882, 60.46421, 60.41936, 
    60.37426, 60.32891, 60.28331, 60.23747, 60.19138, 60.14505, 60.09848, 
    60.05167, 60.00462, 59.95733, 59.90981, 59.86205, 59.81405, 59.76582, 
    59.71735, 59.66866, 59.61974, 59.57058, 59.5212, 59.47159, 59.42176, 
    59.3717, 59.32142, 59.27092, 59.22019, 59.16925, 59.11808, 59.0667, 
    59.0151, 58.96329,
  53.44294, 53.51046, 53.57785, 53.64512, 53.71226, 53.77926, 53.84614, 
    53.91289, 53.9795, 54.04599, 54.11234, 54.17855, 54.24463, 54.31058, 
    54.37639, 54.44206, 54.5076, 54.57299, 54.63824, 54.70336, 54.76833, 
    54.83316, 54.89785, 54.96239, 55.02679, 55.09104, 55.15515, 55.21911, 
    55.28292, 55.34658, 55.4101, 55.47345, 55.53666, 55.59972, 55.66262, 
    55.72537, 55.78797, 55.8504, 55.91269, 55.97481, 56.03677, 56.09857, 
    56.16021, 56.22169, 56.28301, 56.34417, 56.40516, 56.46598, 56.52664, 
    56.58713, 56.64745, 56.7076, 56.76759, 56.8274, 56.88704, 56.9465, 
    57.00579, 57.06491, 57.12385, 57.18261, 57.2412, 57.2996, 57.35782, 
    57.41587, 57.47373, 57.53141, 57.5889, 57.64621, 57.70333, 57.76027, 
    57.81701, 57.87357, 57.92993, 57.98611, 58.04209, 58.09788, 58.15347, 
    58.20887, 58.26407, 58.31907, 58.37387, 58.42848, 58.48288, 58.53708, 
    58.59108, 58.64487, 58.69845, 58.75183, 58.805, 58.85797, 58.91072, 
    58.96326, 59.01559, 59.0677, 59.11961, 59.17129, 59.22276, 59.27401, 
    59.32504, 59.37585, 59.42645, 59.47681, 59.52696, 59.57688, 59.62657, 
    59.67604, 59.72528, 59.77429, 59.82307, 59.87161, 59.91993, 59.96801, 
    60.01585, 60.06347, 60.11084, 60.15797, 60.20486, 60.25151, 60.29792, 
    60.34409, 60.39001, 60.43569, 60.48112, 60.5263, 60.57123, 60.61592, 
    60.66035, 60.70452, 60.74845, 60.79212, 60.83553, 60.87868, 60.92158, 
    60.96422, 61.00659, 61.04871, 61.09056, 61.13214, 61.17346, 61.21452, 
    61.2553, 61.29581, 61.33606, 61.37603, 61.41573, 61.45516, 61.49431, 
    61.53319, 61.57179, 61.61011, 61.64815, 61.68591, 61.72338, 61.76058, 
    61.79749, 61.83411, 61.87045, 61.9065, 61.94226, 61.97773, 62.01291, 
    62.04779, 62.08239, 62.11668, 62.15069, 62.18439, 62.2178, 62.25091, 
    62.28372, 62.31623, 62.34844, 62.38034, 62.41194, 62.44323, 62.47422, 
    62.50489, 62.53526, 62.56532, 62.59507, 62.62451, 62.65364, 62.68245, 
    62.71094, 62.73912, 62.76699, 62.79453, 62.82176, 62.84866, 62.87525, 
    62.90151, 62.92745, 62.95307, 62.97836, 63.00333, 63.02797, 63.05228, 
    63.07627, 63.09993, 63.12325, 63.14624, 63.16891, 63.19124, 63.21323, 
    63.2349, 63.25622, 63.27721, 63.29787, 63.31818, 63.33816, 63.3578, 
    63.3771, 63.39606, 63.41467, 63.43295, 63.45088, 63.46847, 63.48571, 
    63.50261, 63.51916, 63.53537, 63.55122, 63.56674, 63.5819, 63.59671, 
    63.61118, 63.62529, 63.63906, 63.65247, 63.66553, 63.67824, 63.6906, 
    63.7026, 63.71425, 63.72554, 63.73648, 63.74707, 63.7573, 63.76717, 
    63.77669, 63.78585, 63.79465, 63.80309, 63.81118, 63.81891, 63.82628, 
    63.83329, 63.83994, 63.84623, 63.85217, 63.85774, 63.86295, 63.8678, 
    63.8723, 63.87642, 63.88019, 63.8836, 63.88665, 63.88933, 63.89165, 
    63.89362, 63.89522, 63.89646, 63.89733, 63.89785, 63.898, 63.89779, 
    63.89722, 63.89629, 63.89499, 63.89333, 63.89131, 63.88893, 63.88619, 
    63.88309, 63.87962, 63.87579, 63.87161, 63.86706, 63.86215, 63.85688, 
    63.85125, 63.84526, 63.83891, 63.83221, 63.82514, 63.81771, 63.80993, 
    63.80178, 63.79328, 63.78442, 63.7752, 63.76563, 63.7557, 63.74542, 
    63.73478, 63.72378, 63.71243, 63.70073, 63.68867, 63.67625, 63.66349, 
    63.65037, 63.63691, 63.62309, 63.60891, 63.59439, 63.57952, 63.56431, 
    63.54874, 63.53283, 63.51656, 63.49996, 63.48301, 63.46571, 63.44807, 
    63.43008, 63.41175, 63.39308, 63.37407, 63.35472, 63.33503, 63.31499, 
    63.29462, 63.27391, 63.25287, 63.23149, 63.20978, 63.18773, 63.16534, 
    63.14263, 63.11958, 63.09621, 63.0725, 63.04846, 63.02409, 62.9994, 
    62.97438, 62.94904, 62.92337, 62.89738, 62.87106, 62.84443, 62.81747, 
    62.7902, 62.7626, 62.73468, 62.70646, 62.67791, 62.64905, 62.61988, 
    62.59039, 62.56059, 62.53048, 62.50006, 62.46933, 62.4383, 62.40696, 
    62.37531, 62.34336, 62.31111, 62.27855, 62.2457, 62.21254, 62.17908, 
    62.14533, 62.11128, 62.07693, 62.04229, 62.00736, 61.97214, 61.93662, 
    61.90081, 61.86472, 61.82833, 61.79167, 61.75471, 61.71747, 61.67995, 
    61.64215, 61.60406, 61.5657, 61.52706, 61.48814, 61.44894, 61.40947, 
    61.36973, 61.32971, 61.28942, 61.24887, 61.20804, 61.16694, 61.12558, 
    61.08395, 61.04206, 60.99991, 60.95749, 60.91481, 60.87188, 60.82868, 
    60.78522, 60.74152, 60.69755, 60.65334, 60.60886, 60.56414, 60.51917, 
    60.47395, 60.42848, 60.38277, 60.3368, 60.2906, 60.24415, 60.19746, 
    60.15053, 60.10336, 60.05595, 60.0083, 59.96042, 59.9123, 59.86395, 
    59.81536, 59.76655, 59.71751, 59.66823, 59.61873, 59.569, 59.51904, 
    59.46886, 59.41846, 59.36783, 59.31699, 59.26592, 59.21463, 59.16313, 
    59.11141, 59.05947,
  53.52822, 53.59585, 53.66335, 53.73072, 53.79797, 53.86508, 53.93206, 
    53.99892, 54.06564, 54.13223, 54.19869, 54.26502, 54.33121, 54.39726, 
    54.46318, 54.52896, 54.5946, 54.66011, 54.72548, 54.7907, 54.85579, 
    54.92073, 54.98553, 55.05018, 55.11469, 55.17906, 55.24328, 55.30735, 
    55.37127, 55.43505, 55.49868, 55.56215, 55.62547, 55.68864, 55.75166, 
    55.81453, 55.87724, 55.93979, 56.00219, 56.06442, 56.1265, 56.18842, 
    56.25018, 56.31178, 56.37321, 56.43449, 56.49559, 56.55653, 56.61731, 
    56.67792, 56.73836, 56.79863, 56.85873, 56.91866, 56.97842, 57.038, 
    57.09741, 57.15665, 57.21571, 57.27459, 57.33329, 57.39182, 57.45016, 
    57.50833, 57.56631, 57.62411, 57.68172, 57.73915, 57.7964, 57.85345, 
    57.91032, 57.967, 58.02349, 58.07978, 58.13589, 58.1918, 58.24751, 
    58.30303, 58.35835, 58.41348, 58.4684, 58.52313, 58.57765, 58.63197, 
    58.68609, 58.74001, 58.79372, 58.84722, 58.90051, 58.9536, 59.00647, 
    59.05914, 59.11159, 59.16383, 59.21585, 59.26766, 59.31925, 59.37062, 
    59.42178, 59.47271, 59.52343, 59.57392, 59.62418, 59.67422, 59.72404, 
    59.77363, 59.82299, 59.87212, 59.92102, 59.96969, 60.01813, 60.06633, 
    60.1143, 60.16203, 60.20952, 60.25677, 60.30378, 60.35056, 60.39709, 
    60.44337, 60.48942, 60.53521, 60.58076, 60.62606, 60.67111, 60.71592, 
    60.76046, 60.80476, 60.8488, 60.89259, 60.93612, 60.97939, 61.0224, 
    61.06516, 61.10765, 61.14988, 61.19184, 61.23354, 61.27498, 61.31614, 
    61.35704, 61.39767, 61.43803, 61.47812, 61.51793, 61.55747, 61.59673, 
    61.63572, 61.67443, 61.71286, 61.75101, 61.78888, 61.82646, 61.86376, 
    61.90078, 61.93751, 61.97395, 62.01011, 62.04597, 62.08155, 62.11684, 
    62.15182, 62.18652, 62.22092, 62.25503, 62.28884, 62.32235, 62.35556, 
    62.38847, 62.42107, 62.45338, 62.48538, 62.51707, 62.54846, 62.57954, 
    62.61032, 62.64078, 62.67094, 62.70078, 62.7303, 62.75952, 62.78842, 
    62.81701, 62.84528, 62.87323, 62.90086, 62.92817, 62.95517, 62.98183, 
    63.00818, 63.03421, 63.05991, 63.08528, 63.11033, 63.13505, 63.15944, 
    63.18351, 63.20724, 63.23064, 63.25371, 63.27644, 63.29885, 63.32092, 
    63.34265, 63.36405, 63.38511, 63.40583, 63.42621, 63.44626, 63.46596, 
    63.48532, 63.50434, 63.52302, 63.54136, 63.55935, 63.577, 63.5943, 
    63.61125, 63.62786, 63.64412, 63.66003, 63.6756, 63.69081, 63.70568, 
    63.72019, 63.73436, 63.74817, 63.76162, 63.77473, 63.78748, 63.79988, 
    63.81192, 63.82361, 63.83495, 63.84592, 63.85654, 63.86681, 63.87672, 
    63.88626, 63.89546, 63.90429, 63.91277, 63.92088, 63.92863, 63.93603, 
    63.94307, 63.94974, 63.95605, 63.96201, 63.9676, 63.97283, 63.9777, 
    63.9822, 63.98635, 63.99013, 63.99355, 63.99661, 63.9993, 64.00163, 
    64.0036, 64.00521, 64.00645, 64.00733, 64.00784, 64.008, 64.00779, 
    64.00722, 64.00628, 64.00498, 64.00332, 64.00129, 63.9989, 63.99615, 
    63.99303, 63.98956, 63.98572, 63.98151, 63.97695, 63.97203, 63.96674, 
    63.96109, 63.95508, 63.94871, 63.94198, 63.93488, 63.92743, 63.91962, 
    63.91145, 63.90292, 63.89403, 63.88478, 63.87518, 63.86521, 63.85489, 
    63.84421, 63.83318, 63.82179, 63.81004, 63.79794, 63.78549, 63.77268, 
    63.75952, 63.74601, 63.73214, 63.71792, 63.70335, 63.68843, 63.67316, 
    63.65754, 63.64157, 63.62526, 63.60859, 63.59158, 63.57423, 63.55653, 
    63.53848, 63.52009, 63.50136, 63.48228, 63.46287, 63.44311, 63.42301, 
    63.40257, 63.3818, 63.36068, 63.33923, 63.31745, 63.29533, 63.27287, 
    63.25008, 63.22696, 63.20351, 63.17972, 63.15561, 63.13116, 63.10639, 
    63.08129, 63.05586, 63.03011, 63.00404, 62.97764, 62.95092, 62.92387, 
    62.89651, 62.86883, 62.84083, 62.81251, 62.78387, 62.75492, 62.72565, 
    62.69608, 62.66619, 62.63598, 62.60547, 62.57465, 62.54352, 62.51208, 
    62.48034, 62.44829, 62.41594, 62.38328, 62.35032, 62.31707, 62.28351, 
    62.24966, 62.2155, 62.18105, 62.14631, 62.11127, 62.07594, 62.04032, 
    62.00441, 61.96821, 61.93172, 61.89494, 61.85788, 61.82053, 61.78291, 
    61.74499, 61.7068, 61.66832, 61.62957, 61.59054, 61.55123, 61.51165, 
    61.47179, 61.43166, 61.39126, 61.35059, 61.30965, 61.26844, 61.22696, 
    61.18522, 61.14322, 61.10094, 61.05841, 61.01562, 60.97256, 60.92925, 
    60.88568, 60.84185, 60.79777, 60.75343, 60.70884, 60.66401, 60.61891, 
    60.57357, 60.52798, 60.48215, 60.43607, 60.38974, 60.34317, 60.29636, 
    60.24931, 60.20202, 60.15449, 60.10672, 60.05872, 60.01048, 59.96201, 
    59.9133, 59.86436, 59.8152, 59.7658, 59.71618, 59.66632, 59.61625, 
    59.56594, 59.51542, 59.46467, 59.4137, 59.36251, 59.3111, 59.25948, 
    59.20764, 59.15558,
  53.61339, 53.68113, 53.74873, 53.81621, 53.88356, 53.95078, 54.01788, 
    54.08484, 54.15167, 54.21837, 54.28493, 54.35137, 54.41767, 54.48383, 
    54.54986, 54.61575, 54.6815, 54.74712, 54.8126, 54.87793, 54.94313, 
    55.00818, 55.07309, 55.13786, 55.20248, 55.26696, 55.3313, 55.39548, 
    55.45952, 55.52341, 55.58715, 55.65074, 55.71418, 55.77746, 55.8406, 
    55.90358, 55.9664, 56.02907, 56.09158, 56.15393, 56.21613, 56.27817, 
    56.34004, 56.40176, 56.46331, 56.5247, 56.58593, 56.64698, 56.70788, 
    56.7686, 56.82916, 56.88955, 56.94978, 57.00982, 57.0697, 57.12941, 
    57.18893, 57.24829, 57.30747, 57.36647, 57.4253, 57.48394, 57.54241, 
    57.60069, 57.6588, 57.71672, 57.77445, 57.832, 57.88937, 57.94654, 
    58.00354, 58.06034, 58.11695, 58.17336, 58.22959, 58.28562, 58.34146, 
    58.3971, 58.45255, 58.50779, 58.56284, 58.61769, 58.67234, 58.72678, 
    58.78102, 58.83506, 58.88889, 58.94252, 58.99593, 59.04914, 59.10214, 
    59.15493, 59.2075, 59.25986, 59.31201, 59.36395, 59.41566, 59.46716, 
    59.51843, 59.56949, 59.62033, 59.67094, 59.72133, 59.77149, 59.82143, 
    59.87114, 59.92063, 59.96988, 60.0189, 60.06769, 60.11625, 60.16457, 
    60.21266, 60.26051, 60.30813, 60.3555, 60.40264, 60.44953, 60.49618, 
    60.54259, 60.58875, 60.63467, 60.68034, 60.72576, 60.77093, 60.81585, 
    60.86052, 60.90493, 60.94909, 60.993, 61.03664, 61.08003, 61.12317, 
    61.16603, 61.20864, 61.25099, 61.29307, 61.33488, 61.37643, 61.41772, 
    61.45873, 61.49947, 61.53995, 61.58015, 61.62007, 61.65973, 61.6991, 
    61.7382, 61.77702, 61.81556, 61.85382, 61.8918, 61.92949, 61.9669, 
    62.00403, 62.04087, 62.07742, 62.11368, 62.14965, 62.18533, 62.22072, 
    62.25582, 62.29062, 62.32512, 62.35933, 62.39324, 62.42685, 62.46016, 
    62.49317, 62.52588, 62.55828, 62.59038, 62.62217, 62.65366, 62.68484, 
    62.71571, 62.74627, 62.77651, 62.80645, 62.83607, 62.86538, 62.89437, 
    62.92305, 62.9514, 62.97944, 63.00716, 63.03456, 63.06164, 63.0884, 
    63.11483, 63.14094, 63.16672, 63.19218, 63.2173, 63.24211, 63.26658, 
    63.29072, 63.31453, 63.33801, 63.36115, 63.38396, 63.40644, 63.42858, 
    63.45039, 63.47186, 63.49298, 63.51377, 63.53423, 63.55434, 63.57411, 
    63.59354, 63.61262, 63.63136, 63.64976, 63.66781, 63.68552, 63.70288, 
    63.71989, 63.73655, 63.75287, 63.76884, 63.78445, 63.79972, 63.81463, 
    63.8292, 63.84341, 63.85727, 63.87077, 63.88392, 63.89672, 63.90916, 
    63.92125, 63.93297, 63.94435, 63.95536, 63.96602, 63.97632, 63.98626, 
    63.99584, 64.00507, 64.01393, 64.02243, 64.03058, 64.03836, 64.04578, 
    64.05284, 64.05954, 64.06587, 64.07185, 64.07746, 64.08271, 64.08759, 
    64.09212, 64.09628, 64.10007, 64.1035, 64.10657, 64.10928, 64.11161, 
    64.11359, 64.1152, 64.11645, 64.11732, 64.11784, 64.118, 64.11779, 
    64.11721, 64.11627, 64.11497, 64.1133, 64.11127, 64.10887, 64.10611, 
    64.10298, 64.09949, 64.09564, 64.09142, 64.08685, 64.0819, 64.07659, 
    64.07092, 64.0649, 64.0585, 64.05174, 64.04463, 64.03715, 64.02931, 
    64.02111, 64.01255, 64.00363, 63.99435, 63.98471, 63.97471, 63.96436, 
    63.95364, 63.94257, 63.93114, 63.91936, 63.90722, 63.89472, 63.88187, 
    63.86866, 63.8551, 63.84118, 63.82692, 63.8123, 63.79733, 63.78201, 
    63.76633, 63.75031, 63.73394, 63.71722, 63.70015, 63.68274, 63.66498, 
    63.64687, 63.62842, 63.60962, 63.59048, 63.571, 63.55118, 63.53101, 
    63.51051, 63.48967, 63.46848, 63.44696, 63.4251, 63.40291, 63.38038, 
    63.35751, 63.33432, 63.31078, 63.28692, 63.26273, 63.2382, 63.21335, 
    63.18817, 63.16267, 63.13683, 63.11067, 63.08419, 63.05738, 63.03025, 
    63.0028, 62.97503, 62.94694, 62.91853, 62.8898, 62.86076, 62.83141, 
    62.80173, 62.77175, 62.74145, 62.71085, 62.67993, 62.6487, 62.61716, 
    62.58532, 62.55318, 62.52073, 62.48797, 62.45491, 62.42155, 62.3879, 
    62.35394, 62.31968, 62.28513, 62.25029, 62.21515, 62.17971, 62.14398, 
    62.10796, 62.07166, 62.03506, 61.99817, 61.961, 61.92355, 61.88581, 
    61.84779, 61.80948, 61.7709, 61.73203, 61.69289, 61.65347, 61.61377, 
    61.57381, 61.53356, 61.49305, 61.45226, 61.41121, 61.36988, 61.32829, 
    61.28643, 61.24431, 61.20192, 61.15927, 61.11636, 61.07319, 61.02975, 
    60.98607, 60.94212, 60.89792, 60.85347, 60.80876, 60.7638, 60.71859, 
    60.67313, 60.62742, 60.58147, 60.53527, 60.48882, 60.44213, 60.3952, 
    60.34803, 60.30061, 60.25296, 60.20507, 60.15695, 60.10859, 60.05999, 
    60.01116, 59.9621, 59.91282, 59.8633, 59.81355, 59.76357, 59.71337, 
    59.66295, 59.6123, 59.56143, 59.51034, 59.45902, 59.40749, 59.35574, 
    59.30378, 59.2516,
  53.69845, 53.76628, 53.834, 53.90158, 53.96904, 54.03637, 54.10357, 
    54.17064, 54.23758, 54.30439, 54.37106, 54.43761, 54.50401, 54.57029, 
    54.63643, 54.70243, 54.76829, 54.83402, 54.8996, 54.96505, 55.03036, 
    55.09553, 55.16055, 55.22543, 55.29016, 55.35476, 55.4192, 55.4835, 
    55.54765, 55.61166, 55.67551, 55.73922, 55.80277, 55.86617, 55.92942, 
    55.99252, 56.05545, 56.11824, 56.18087, 56.24334, 56.30565, 56.36781, 
    56.4298, 56.49163, 56.5533, 56.61481, 56.67615, 56.73733, 56.79834, 
    56.85919, 56.91986, 56.98038, 57.04071, 57.10088, 57.16088, 57.2207, 
    57.28036, 57.33983, 57.39913, 57.45826, 57.5172, 57.57597, 57.63456, 
    57.69296, 57.75119, 57.80923, 57.86708, 57.92476, 57.98224, 58.03954, 
    58.09666, 58.15358, 58.21031, 58.26685, 58.3232, 58.37935, 58.43531, 
    58.49108, 58.54665, 58.60202, 58.65719, 58.71216, 58.76693, 58.8215, 
    58.87587, 58.93003, 58.98398, 59.03773, 59.09127, 59.1446, 59.19772, 
    59.25064, 59.30333, 59.35582, 59.40809, 59.46014, 59.51198, 59.5636, 
    59.61501, 59.66618, 59.71714, 59.76788, 59.81839, 59.86868, 59.91874, 
    59.96858, 60.01818, 60.06756, 60.11671, 60.16562, 60.2143, 60.26274, 
    60.31096, 60.35893, 60.40667, 60.45416, 60.50142, 60.54844, 60.59521, 
    60.64174, 60.68802, 60.73405, 60.77985, 60.82539, 60.87068, 60.91571, 
    60.9605, 61.00504, 61.04932, 61.09334, 61.13711, 61.18061, 61.22386, 
    61.26685, 61.30957, 61.35204, 61.39424, 61.43617, 61.47783, 61.51923, 
    61.56036, 61.60122, 61.64181, 61.68212, 61.72216, 61.76192, 61.80141, 
    61.84062, 61.87955, 61.91821, 61.95658, 61.99467, 62.03247, 62.06999, 
    62.10723, 62.14417, 62.18083, 62.2172, 62.25328, 62.28907, 62.32457, 
    62.35976, 62.39467, 62.42928, 62.46359, 62.4976, 62.53132, 62.56473, 
    62.59784, 62.63065, 62.66315, 62.69535, 62.72724, 62.75882, 62.7901, 
    62.82106, 62.85172, 62.88206, 62.91209, 62.9418, 62.9712, 63.00029, 
    63.02905, 63.0575, 63.08563, 63.11344, 63.14093, 63.16809, 63.19493, 
    63.22145, 63.24765, 63.27351, 63.29905, 63.32426, 63.34914, 63.37369, 
    63.39791, 63.4218, 63.44535, 63.46858, 63.49146, 63.51402, 63.53623, 
    63.55811, 63.57965, 63.60085, 63.62171, 63.64223, 63.6624, 63.68224, 
    63.70173, 63.72088, 63.73969, 63.75814, 63.77626, 63.79403, 63.81144, 
    63.82851, 63.84523, 63.86161, 63.87763, 63.8933, 63.90862, 63.92358, 
    63.93819, 63.95245, 63.96636, 63.97991, 63.99311, 64.00595, 64.01843, 
    64.03056, 64.04233, 64.05374, 64.0648, 64.07549, 64.08582, 64.0958, 
    64.10542, 64.11467, 64.12357, 64.1321, 64.14027, 64.14808, 64.15553, 
    64.16261, 64.16933, 64.17569, 64.18169, 64.18732, 64.19258, 64.19749, 
    64.20203, 64.2062, 64.21001, 64.21345, 64.21653, 64.21924, 64.22159, 
    64.22357, 64.22519, 64.22644, 64.22733, 64.22784, 64.228, 64.22779, 
    64.22721, 64.22626, 64.22496, 64.22328, 64.22124, 64.21883, 64.21606, 
    64.21293, 64.20943, 64.20556, 64.20133, 64.19673, 64.19177, 64.18645, 
    64.18076, 64.17471, 64.16829, 64.16151, 64.15437, 64.14687, 64.139, 
    64.13078, 64.12218, 64.11323, 64.10392, 64.09425, 64.08421, 64.07382, 
    64.06307, 64.05196, 64.04049, 64.02866, 64.01648, 64.00394, 63.99104, 
    63.97779, 63.96418, 63.95022, 63.93591, 63.92124, 63.90622, 63.89084, 
    63.87511, 63.85904, 63.84261, 63.82584, 63.80871, 63.79124, 63.77341, 
    63.75525, 63.73674, 63.71788, 63.69867, 63.67913, 63.65924, 63.639, 
    63.61843, 63.59752, 63.57626, 63.55467, 63.53274, 63.51047, 63.48787, 
    63.46493, 63.44165, 63.41805, 63.3941, 63.36983, 63.34523, 63.32029, 
    63.29503, 63.26944, 63.24352, 63.21728, 63.19071, 63.16382, 63.1366, 
    63.10906, 63.0812, 63.05302, 63.02452, 62.99571, 62.96658, 62.93712, 
    62.90736, 62.87728, 62.84689, 62.81618, 62.78517, 62.75385, 62.72221, 
    62.69027, 62.65803, 62.62548, 62.59262, 62.55946, 62.526, 62.49224, 
    62.45818, 62.42382, 62.38917, 62.35422, 62.31897, 62.28343, 62.24759, 
    62.21147, 62.17505, 62.13835, 62.10136, 62.06408, 62.02651, 61.98866, 
    61.95053, 61.91211, 61.87342, 61.83444, 61.79519, 61.75565, 61.71584, 
    61.67576, 61.6354, 61.59478, 61.55387, 61.5127, 61.47126, 61.42955, 
    61.38758, 61.34534, 61.30283, 61.26007, 61.21704, 61.17375, 61.1302, 
    61.0864, 61.04233, 60.99801, 60.95343, 60.90861, 60.86353, 60.8182, 
    60.77262, 60.72679, 60.68071, 60.63439, 60.58783, 60.54101, 60.49396, 
    60.44667, 60.39913, 60.35136, 60.30334, 60.2551, 60.20662, 60.1579, 
    60.10895, 60.05976, 60.01035, 59.96071, 59.91084, 59.86074, 59.81042, 
    59.75987, 59.7091, 59.6581, 59.60689, 59.55545, 59.5038, 59.45192, 
    59.39984, 59.34753,
  53.78339, 53.85133, 53.91915, 53.98684, 54.05441, 54.12185, 54.18915, 
    54.25633, 54.32338, 54.39029, 54.45708, 54.52373, 54.59025, 54.65663, 
    54.72288, 54.78899, 54.85497, 54.9208, 54.9865, 55.05206, 55.11748, 
    55.18276, 55.24789, 55.31289, 55.37774, 55.44244, 55.507, 55.57141, 
    55.63568, 55.6998, 55.76377, 55.82759, 55.89125, 55.95477, 56.01814, 
    56.08134, 56.1444, 56.2073, 56.27005, 56.33264, 56.39507, 56.45734, 
    56.51945, 56.5814, 56.64318, 56.70481, 56.76627, 56.82757, 56.8887, 
    56.94967, 57.01046, 57.07109, 57.13155, 57.19184, 57.25196, 57.3119, 
    57.37167, 57.43127, 57.49069, 57.54993, 57.609, 57.66789, 57.7266, 
    57.78513, 57.84348, 57.90164, 57.95962, 58.01741, 58.07502, 58.13244, 
    58.18968, 58.24672, 58.30358, 58.36024, 58.41671, 58.47299, 58.52908, 
    58.58496, 58.64066, 58.69615, 58.75145, 58.80654, 58.86143, 58.91613, 
    58.97062, 59.0249, 59.07898, 59.13285, 59.18652, 59.23997, 59.29322, 
    59.34626, 59.39908, 59.45169, 59.50408, 59.55626, 59.60822, 59.65997, 
    59.71149, 59.7628, 59.81388, 59.86474, 59.91538, 59.96579, 60.01598, 
    60.06593, 60.11566, 60.16516, 60.21443, 60.26347, 60.31227, 60.36084, 
    60.40918, 60.45727, 60.50513, 60.55275, 60.60013, 60.64727, 60.69416, 
    60.74081, 60.78721, 60.83337, 60.87928, 60.92495, 60.97036, 61.01552, 
    61.06042, 61.10508, 61.14948, 61.19362, 61.23751, 61.28113, 61.3245, 
    61.3676, 61.41045, 61.45303, 61.49534, 61.53739, 61.57917, 61.62069, 
    61.66193, 61.70291, 61.74361, 61.78404, 61.82419, 61.86407, 61.90367, 
    61.943, 61.98204, 62.02081, 62.05929, 62.09749, 62.1354, 62.17303, 
    62.21038, 62.24744, 62.2842, 62.32068, 62.35687, 62.39276, 62.42836, 
    62.46367, 62.49868, 62.53339, 62.56781, 62.60192, 62.63574, 62.66926, 
    62.70247, 62.73538, 62.76798, 62.80028, 62.83227, 62.86395, 62.89532, 
    62.92638, 62.95713, 62.98757, 63.0177, 63.0475, 63.077, 63.10617, 
    63.13503, 63.16357, 63.19179, 63.21969, 63.24726, 63.27452, 63.30145, 
    63.32805, 63.35433, 63.38028, 63.4059, 63.43119, 63.45615, 63.48079, 
    63.50508, 63.52905, 63.55268, 63.57598, 63.59895, 63.62157, 63.64386, 
    63.66581, 63.68742, 63.70869, 63.72962, 63.75021, 63.77045, 63.79036, 
    63.80992, 63.82913, 63.848, 63.86652, 63.88469, 63.90252, 63.92, 
    63.93713, 63.9539, 63.97033, 63.98641, 64.00213, 64.0175, 64.03252, 
    64.04719, 64.06149, 64.07545, 64.08904, 64.10229, 64.11517, 64.1277, 
    64.13987, 64.15168, 64.16313, 64.17422, 64.18495, 64.19533, 64.20534, 
    64.21499, 64.22427, 64.2332, 64.24176, 64.24996, 64.2578, 64.26527, 
    64.27238, 64.27913, 64.28551, 64.29152, 64.29717, 64.30246, 64.30738, 
    64.31194, 64.31612, 64.31994, 64.32339, 64.32648, 64.32921, 64.33157, 
    64.33356, 64.33518, 64.33643, 64.33733, 64.33784, 64.338, 64.33778, 
    64.3372, 64.33626, 64.33495, 64.33327, 64.33121, 64.3288, 64.32603, 
    64.32288, 64.31936, 64.31548, 64.31123, 64.30663, 64.30164, 64.2963, 
    64.2906, 64.28452, 64.27808, 64.27128, 64.26411, 64.25658, 64.24869, 
    64.24043, 64.23181, 64.22282, 64.21349, 64.20377, 64.19371, 64.18328, 
    64.17249, 64.16134, 64.14983, 64.13797, 64.12574, 64.11316, 64.10022, 
    64.08692, 64.07327, 64.05926, 64.04489, 64.03017, 64.0151, 63.99967, 
    63.98389, 63.96776, 63.95127, 63.93444, 63.91726, 63.89972, 63.88184, 
    63.86361, 63.84504, 63.82611, 63.80685, 63.78723, 63.76728, 63.74697, 
    63.72633, 63.70535, 63.68402, 63.66236, 63.64035, 63.61802, 63.59533, 
    63.57232, 63.54897, 63.52528, 63.50126, 63.47691, 63.45223, 63.42721, 
    63.40187, 63.37619, 63.35019, 63.32386, 63.29721, 63.27023, 63.24292, 
    63.2153, 63.18735, 63.15908, 63.13049, 63.10158, 63.07235, 63.04281, 
    63.01295, 62.98278, 62.95229, 62.92149, 62.89038, 62.85896, 62.82723, 
    62.79519, 62.76284, 62.73019, 62.69724, 62.66397, 62.63041, 62.59655, 
    62.56239, 62.52792, 62.49316, 62.4581, 62.42275, 62.3871, 62.35116, 
    62.31493, 62.2784, 62.24159, 62.20449, 62.1671, 62.12943, 62.09146, 
    62.05322, 62.01469, 61.97588, 61.93679, 61.89743, 61.85778, 61.81786, 
    61.77766, 61.73719, 61.69645, 61.65543, 61.61414, 61.57259, 61.53076, 
    61.48867, 61.44631, 61.40369, 61.36081, 61.31766, 61.27425, 61.23058, 
    61.18665, 61.14247, 61.09803, 61.05334, 61.00839, 60.96319, 60.91774, 
    60.87204, 60.82609, 60.77989, 60.73345, 60.68676, 60.63982, 60.59265, 
    60.54523, 60.49757, 60.44968, 60.40155, 60.35318, 60.30457, 60.25573, 
    60.20665, 60.15735, 60.10781, 60.05804, 60.00805, 59.95783, 59.90738, 
    59.85671, 59.80582, 59.7547, 59.70336, 59.6518, 59.60002, 59.54802, 
    59.49581, 59.44338,
  53.86821, 53.93626, 54.00418, 54.07198, 54.13966, 54.2072, 54.27462, 
    54.3419, 54.40906, 54.47609, 54.54298, 54.60974, 54.67636, 54.74286, 
    54.80922, 54.87544, 54.94153, 55.00748, 55.07328, 55.13896, 55.20449, 
    55.26988, 55.33512, 55.40023, 55.46519, 55.53001, 55.59468, 55.65921, 
    55.72359, 55.78783, 55.85191, 55.91584, 55.97963, 56.04326, 56.10674, 
    56.17007, 56.23324, 56.29626, 56.35912, 56.42183, 56.48437, 56.54676, 
    56.60899, 56.67106, 56.73296, 56.79471, 56.85629, 56.91771, 56.97896, 
    57.04004, 57.10096, 57.16171, 57.22229, 57.2827, 57.34293, 57.403, 
    57.46289, 57.52261, 57.58215, 57.64151, 57.7007, 57.75972, 57.81855, 
    57.87719, 57.93567, 57.99395, 58.05205, 58.10997, 58.1677, 58.22525, 
    58.2826, 58.33977, 58.39675, 58.45354, 58.51014, 58.56654, 58.62274, 
    58.67876, 58.73457, 58.79019, 58.84561, 58.90083, 58.95585, 59.01067, 
    59.06528, 59.11969, 59.17389, 59.22789, 59.28168, 59.33526, 59.38863, 
    59.44179, 59.49474, 59.54747, 59.59999, 59.65229, 59.70438, 59.75625, 
    59.8079, 59.85933, 59.91053, 59.96152, 60.01228, 60.06282, 60.11313, 
    60.16321, 60.21306, 60.26269, 60.31208, 60.36124, 60.41017, 60.45886, 
    60.50732, 60.55554, 60.60352, 60.65126, 60.69876, 60.74602, 60.79304, 
    60.83981, 60.88634, 60.93262, 60.97865, 61.02444, 61.06997, 61.11525, 
    61.16028, 61.20505, 61.24957, 61.29383, 61.33784, 61.38159, 61.42507, 
    61.4683, 61.51126, 61.55396, 61.59639, 61.63856, 61.68046, 61.72209, 
    61.76345, 61.80454, 61.84536, 61.8859, 61.92617, 61.96616, 62.00588, 
    62.04532, 62.08448, 62.12335, 62.16195, 62.20026, 62.23829, 62.27603, 
    62.31348, 62.35065, 62.38752, 62.42411, 62.46041, 62.49641, 62.53212, 
    62.56753, 62.60265, 62.63747, 62.67199, 62.70621, 62.74013, 62.77375, 
    62.80706, 62.84007, 62.87277, 62.90517, 62.93726, 62.96904, 63.00051, 
    63.03167, 63.06252, 63.09305, 63.12327, 63.15318, 63.18276, 63.21203, 
    63.24098, 63.26961, 63.29792, 63.32591, 63.35357, 63.38091, 63.40793, 
    63.43462, 63.46098, 63.48702, 63.51272, 63.5381, 63.56314, 63.58786, 
    63.61224, 63.63628, 63.65999, 63.68337, 63.70641, 63.72911, 63.75147, 
    63.77349, 63.79518, 63.81652, 63.83752, 63.85818, 63.87849, 63.89846, 
    63.91809, 63.93737, 63.9563, 63.97488, 63.99312, 64.011, 64.02854, 
    64.04573, 64.06257, 64.07905, 64.09518, 64.11096, 64.12638, 64.14145, 
    64.15617, 64.17052, 64.18452, 64.19817, 64.21146, 64.22439, 64.23696, 
    64.24917, 64.26102, 64.27251, 64.28365, 64.29442, 64.30482, 64.31487, 
    64.32455, 64.33387, 64.34283, 64.35142, 64.35965, 64.36752, 64.37502, 
    64.38215, 64.38892, 64.39532, 64.40136, 64.40703, 64.41233, 64.41727, 
    64.42184, 64.42604, 64.42988, 64.43335, 64.43645, 64.43918, 64.44154, 
    64.44354, 64.44517, 64.44643, 64.44732, 64.44785, 64.448, 64.44778, 
    64.4472, 64.44625, 64.44494, 64.44325, 64.44119, 64.43877, 64.43598, 
    64.43282, 64.4293, 64.4254, 64.42114, 64.41651, 64.41151, 64.40616, 
    64.40043, 64.39433, 64.38787, 64.38104, 64.37386, 64.36629, 64.35838, 
    64.35009, 64.34144, 64.33242, 64.32304, 64.3133, 64.3032, 64.29273, 
    64.28191, 64.27072, 64.25917, 64.24726, 64.23499, 64.22237, 64.20938, 
    64.19604, 64.18233, 64.16827, 64.15386, 64.13909, 64.12396, 64.10848, 
    64.09265, 64.07646, 64.05993, 64.04304, 64.02579, 64.0082, 63.99026, 
    63.97197, 63.95333, 63.93434, 63.915, 63.89532, 63.8753, 63.85493, 
    63.83422, 63.81317, 63.79177, 63.77003, 63.74796, 63.72554, 63.70279, 
    63.67969, 63.65627, 63.6325, 63.6084, 63.58397, 63.5592, 63.53411, 
    63.50868, 63.48292, 63.45683, 63.43042, 63.40368, 63.37661, 63.34922, 
    63.3215, 63.29346, 63.2651, 63.23642, 63.20742, 63.1781, 63.14846, 
    63.11851, 63.08824, 63.05766, 63.02676, 62.99556, 62.96404, 62.93221, 
    62.90007, 62.86762, 62.83487, 62.80181, 62.76845, 62.73478, 62.70081, 
    62.66655, 62.63198, 62.59711, 62.56195, 62.52649, 62.49073, 62.45469, 
    62.41834, 62.38171, 62.34479, 62.30758, 62.27008, 62.23229, 62.19422, 
    62.15586, 62.11722, 62.0783, 62.0391, 61.99961, 61.95985, 61.91982, 
    61.87951, 61.83892, 61.79806, 61.75692, 61.71552, 61.67385, 61.6319, 
    61.58969, 61.54722, 61.50448, 61.46148, 61.41821, 61.37468, 61.3309, 
    61.28685, 61.24255, 61.19799, 61.15317, 61.1081, 61.06278, 61.01721, 
    60.97139, 60.92532, 60.879, 60.83243, 60.78562, 60.73856, 60.69127, 
    60.64373, 60.59595, 60.54793, 60.49967, 60.45118, 60.40244, 60.35348, 
    60.30428, 60.25485, 60.20519, 60.1553, 60.10518, 60.05484, 60.00427, 
    59.95347, 59.90245, 59.85121, 59.79974, 59.74806, 59.69616, 59.64404, 
    59.5917, 59.53914,
  53.95292, 54.02107, 54.0891, 54.15701, 54.22479, 54.29244, 54.35997, 
    54.42736, 54.49463, 54.56176, 54.62876, 54.69563, 54.76237, 54.82897, 
    54.89544, 54.96178, 55.02797, 55.09403, 55.15995, 55.22574, 55.29138, 
    55.35688, 55.42225, 55.48746, 55.55254, 55.61747, 55.68226, 55.7469, 
    55.81139, 55.87574, 55.93994, 56.00399, 56.06789, 56.13164, 56.19524, 
    56.25868, 56.32197, 56.3851, 56.44808, 56.51091, 56.57357, 56.63608, 
    56.69843, 56.76061, 56.82264, 56.8845, 56.9462, 57.00773, 57.0691, 
    57.13031, 57.19135, 57.25222, 57.31292, 57.37344, 57.4338, 57.49399, 
    57.554, 57.61384, 57.6735, 57.73299, 57.7923, 57.85144, 57.91039, 
    57.96916, 58.02775, 58.08616, 58.14439, 58.20243, 58.26028, 58.31795, 
    58.37543, 58.43272, 58.48983, 58.54674, 58.60346, 58.65998, 58.71632, 
    58.77245, 58.82839, 58.88414, 58.93968, 58.99502, 59.05017, 59.10511, 
    59.15985, 59.21438, 59.26871, 59.32283, 59.37675, 59.43045, 59.48395, 
    59.53723, 59.59031, 59.64317, 59.69581, 59.74824, 59.80045, 59.85244, 
    59.90422, 59.95577, 60.00711, 60.05822, 60.1091, 60.15976, 60.2102, 
    60.26041, 60.31038, 60.36013, 60.40965, 60.45893, 60.50799, 60.5568, 
    60.60538, 60.65373, 60.70183, 60.7497, 60.79733, 60.84471, 60.89185, 
    60.93874, 60.98539, 61.0318, 61.07795, 61.12386, 61.16951, 61.21492, 
    61.26006, 61.30496, 61.3496, 61.39399, 61.43811, 61.48198, 61.52558, 
    61.56893, 61.61201, 61.65483, 61.69738, 61.73966, 61.78168, 61.82343, 
    61.86491, 61.90611, 61.94705, 61.98771, 62.02809, 62.0682, 62.10803, 
    62.14758, 62.18686, 62.22585, 62.26455, 62.30298, 62.34112, 62.37897, 
    62.41653, 62.45381, 62.4908, 62.5275, 62.5639, 62.60001, 62.63583, 
    62.67135, 62.70657, 62.7415, 62.77612, 62.81045, 62.84447, 62.87819, 
    62.91161, 62.94472, 62.97753, 63.01003, 63.04222, 63.0741, 63.10567, 
    63.13692, 63.16787, 63.1985, 63.22881, 63.25881, 63.28849, 63.31786, 
    63.3469, 63.37562, 63.40402, 63.4321, 63.45985, 63.48729, 63.51439, 
    63.54116, 63.56761, 63.59373, 63.61952, 63.64498, 63.67011, 63.6949, 
    63.71936, 63.74349, 63.76728, 63.79073, 63.81385, 63.83662, 63.85906, 
    63.88116, 63.90292, 63.92433, 63.9454, 63.96613, 63.98651, 64.00655, 
    64.02625, 64.04559, 64.06458, 64.08323, 64.10153, 64.11948, 64.13708, 
    64.15432, 64.17122, 64.18776, 64.20394, 64.21977, 64.23525, 64.25037, 
    64.26514, 64.27955, 64.2936, 64.30729, 64.32063, 64.3336, 64.34621, 
    64.35847, 64.37036, 64.3819, 64.39307, 64.40387, 64.41431, 64.4244, 
    64.43411, 64.44347, 64.45245, 64.46108, 64.46934, 64.47723, 64.48476, 
    64.49191, 64.49871, 64.50513, 64.51119, 64.51688, 64.5222, 64.52716, 
    64.53175, 64.53596, 64.53981, 64.5433, 64.5464, 64.54915, 64.55152, 
    64.55353, 64.55516, 64.55642, 64.55732, 64.55785, 64.558, 64.55779, 
    64.5572, 64.55624, 64.55492, 64.55323, 64.55117, 64.54874, 64.54594, 
    64.54277, 64.53923, 64.53532, 64.53104, 64.5264, 64.52139, 64.51601, 
    64.51025, 64.50414, 64.49766, 64.49081, 64.48359, 64.47601, 64.46806, 
    64.45974, 64.45106, 64.44201, 64.4326, 64.42283, 64.41269, 64.40218, 
    64.39132, 64.3801, 64.36851, 64.35655, 64.34425, 64.33157, 64.31854, 
    64.30515, 64.2914, 64.27729, 64.26283, 64.24801, 64.23283, 64.21729, 
    64.20141, 64.18517, 64.16856, 64.15162, 64.13432, 64.11666, 64.09866, 
    64.08031, 64.0616, 64.04255, 64.02315, 64.0034, 63.98331, 63.96288, 
    63.94209, 63.92097, 63.8995, 63.87769, 63.85554, 63.83305, 63.81021, 
    63.78704, 63.76354, 63.7397, 63.71552, 63.691, 63.66616, 63.64098, 
    63.61547, 63.58962, 63.56345, 63.53695, 63.51012, 63.48297, 63.45549, 
    63.42768, 63.39955, 63.3711, 63.34233, 63.31323, 63.28382, 63.25409, 
    63.22404, 63.19367, 63.16299, 63.132, 63.10069, 63.06907, 63.03714, 
    63.00491, 62.97236, 62.9395, 62.90635, 62.87288, 62.83911, 62.80504, 
    62.77066, 62.73599, 62.70102, 62.66575, 62.63018, 62.59432, 62.55816, 
    62.52171, 62.48497, 62.44793, 62.41061, 62.373, 62.3351, 62.29692, 
    62.25845, 62.2197, 62.18066, 62.14135, 62.10175, 62.06187, 62.02172, 
    61.98129, 61.94059, 61.89961, 61.85836, 61.81684, 61.77505, 61.73299, 
    61.69066, 61.64807, 61.60521, 61.56209, 61.5187, 61.47506, 61.43115, 
    61.38698, 61.34256, 61.29787, 61.25294, 61.20775, 61.16231, 61.11661, 
    61.07067, 61.02447, 60.97803, 60.93134, 60.88441, 60.83723, 60.78981, 
    60.74215, 60.69424, 60.6461, 60.59772, 60.5491, 60.50024, 60.45115, 
    60.40183, 60.35228, 60.30249, 60.25248, 60.20224, 60.15176, 60.10107, 
    60.05015, 59.999, 59.94763, 59.89605, 59.84423, 59.79221, 59.73996, 
    59.6875, 59.63482,
  54.0375, 54.10577, 54.1739, 54.24192, 54.30981, 54.37756, 54.4452, 54.5127, 
    54.58007, 54.64732, 54.71443, 54.78141, 54.84826, 54.91497, 54.98155, 
    55.04799, 55.1143, 55.18047, 55.24651, 55.3124, 55.37816, 55.44378, 
    55.50925, 55.57458, 55.63977, 55.70481, 55.76972, 55.83447, 55.89908, 
    55.96355, 56.02786, 56.09203, 56.15604, 56.21991, 56.28362, 56.34718, 
    56.41058, 56.47384, 56.53693, 56.59987, 56.66266, 56.72528, 56.78775, 
    56.85005, 56.9122, 56.97418, 57.036, 57.09766, 57.15915, 57.22047, 
    57.28163, 57.34262, 57.40343, 57.46409, 57.52457, 57.58487, 57.64501, 
    57.70497, 57.76476, 57.82437, 57.8838, 57.94305, 58.00213, 58.06102, 
    58.11974, 58.17827, 58.23662, 58.29478, 58.35276, 58.41056, 58.46816, 
    58.52558, 58.5828, 58.63984, 58.69668, 58.75333, 58.80979, 58.86605, 
    58.92212, 58.97799, 59.03365, 59.08912, 59.14439, 59.19946, 59.25432, 
    59.30898, 59.36344, 59.41768, 59.47173, 59.52555, 59.57918, 59.63259, 
    59.68579, 59.73877, 59.79154, 59.8441, 59.89643, 59.94855, 60.00045, 
    60.05214, 60.10359, 60.15483, 60.20584, 60.25663, 60.30719, 60.35752, 
    60.40762, 60.4575, 60.50714, 60.55655, 60.60573, 60.65467, 60.70337, 
    60.75184, 60.80007, 60.84806, 60.89581, 60.94332, 60.99058, 61.0376, 
    61.08437, 61.1309, 61.17718, 61.22321, 61.26899, 61.31451, 61.35978, 
    61.4048, 61.44956, 61.49407, 61.53831, 61.5823, 61.62603, 61.66949, 
    61.71269, 61.75563, 61.7983, 61.84071, 61.88284, 61.92471, 61.9663, 
    62.00763, 62.04868, 62.08946, 62.12996, 62.17018, 62.21013, 62.24979, 
    62.28918, 62.32829, 62.36711, 62.40564, 62.4439, 62.48186, 62.51954, 
    62.55693, 62.59402, 62.63083, 62.66735, 62.70357, 62.73949, 62.77512, 
    62.81045, 62.84548, 62.88021, 62.91465, 62.94877, 62.9826, 63.01612, 
    63.04934, 63.08224, 63.11484, 63.14713, 63.17912, 63.21078, 63.24214, 
    63.27318, 63.30391, 63.33432, 63.36441, 63.39419, 63.42365, 63.45279, 
    63.4816, 63.51009, 63.53827, 63.56611, 63.59363, 63.62082, 63.64768, 
    63.67422, 63.70042, 63.7263, 63.75184, 63.77705, 63.80193, 63.82647, 
    63.85068, 63.87455, 63.89808, 63.92127, 63.94412, 63.96664, 63.98881, 
    64.01064, 64.03213, 64.05327, 64.07407, 64.09452, 64.11462, 64.13438, 
    64.15379, 64.17285, 64.19157, 64.20993, 64.22794, 64.2456, 64.2629, 
    64.27985, 64.29646, 64.3127, 64.32858, 64.34412, 64.35929, 64.37411, 
    64.38857, 64.40266, 64.4164, 64.42979, 64.4428, 64.45547, 64.46776, 
    64.4797, 64.49127, 64.50248, 64.51332, 64.5238, 64.53392, 64.54367, 
    64.55306, 64.56208, 64.57073, 64.57902, 64.58694, 64.59449, 64.60168, 
    64.6085, 64.61494, 64.62103, 64.62673, 64.63208, 64.63705, 64.64165, 
    64.64589, 64.64975, 64.65324, 64.65636, 64.65912, 64.6615, 64.66351, 
    64.66515, 64.66642, 64.66731, 64.66784, 64.668, 64.66779, 64.6672, 
    64.66624, 64.66492, 64.66322, 64.66115, 64.65871, 64.65589, 64.65272, 
    64.64916, 64.64524, 64.64095, 64.63629, 64.63126, 64.62585, 64.62009, 
    64.61395, 64.60744, 64.60056, 64.59332, 64.58571, 64.57774, 64.56939, 
    64.56068, 64.5516, 64.54215, 64.53235, 64.52217, 64.51163, 64.50073, 
    64.48946, 64.47783, 64.46584, 64.45348, 64.44077, 64.4277, 64.41425, 
    64.40046, 64.3863, 64.37179, 64.35691, 64.34168, 64.3261, 64.31015, 
    64.29385, 64.2772, 64.26019, 64.24283, 64.22511, 64.20705, 64.18863, 
    64.16986, 64.15075, 64.13128, 64.11147, 64.09131, 64.0708, 64.04995, 
    64.02875, 64.00721, 63.98532, 63.9631, 63.94053, 63.91763, 63.89438, 
    63.87079, 63.84687, 63.82261, 63.79802, 63.77309, 63.74782, 63.72223, 
    63.6963, 63.67004, 63.64346, 63.61654, 63.58929, 63.56173, 63.53383, 
    63.50561, 63.47707, 63.4482, 63.41901, 63.3895, 63.35968, 63.32953, 
    63.29907, 63.26829, 63.2372, 63.2058, 63.17408, 63.14205, 63.10971, 
    63.07706, 63.0441, 63.01084, 62.97727, 62.94339, 62.90922, 62.87474, 
    62.83996, 62.80488, 62.7695, 62.73383, 62.69786, 62.66159, 62.62503, 
    62.58818, 62.55103, 62.5136, 62.47588, 62.43787, 62.39957, 62.36098, 
    62.32212, 62.28297, 62.24354, 62.20383, 62.16384, 62.12357, 62.08302, 
    62.04221, 62.00111, 61.95974, 61.9181, 61.87619, 61.83401, 61.79157, 
    61.74886, 61.70588, 61.66264, 61.61913, 61.57536, 61.53133, 61.48705, 
    61.4425, 61.3977, 61.35264, 61.30733, 61.26176, 61.21594, 61.16988, 
    61.12356, 61.07699, 61.03018, 60.98312, 60.93582, 60.88828, 60.84049, 
    60.79246, 60.74419, 60.69569, 60.64694, 60.59796, 60.54875, 60.4993, 
    60.44962, 60.39971, 60.34957, 60.29921, 60.24861, 60.19778, 60.14674, 
    60.09547, 60.04398, 59.99226, 59.94032, 59.88817, 59.8358, 59.78321, 
    59.7304,
  54.12197, 54.19034, 54.25859, 54.32671, 54.3947, 54.46257, 54.53031, 
    54.59792, 54.66541, 54.73276, 54.79998, 54.86707, 54.93402, 55.00085, 
    55.06754, 55.13409, 55.20052, 55.2668, 55.33294, 55.39895, 55.46482, 
    55.53055, 55.59614, 55.66158, 55.72689, 55.79205, 55.85706, 55.92193, 
    55.98666, 56.05124, 56.11567, 56.17995, 56.24408, 56.30806, 56.37189, 
    56.43557, 56.49909, 56.56246, 56.62568, 56.68873, 56.75163, 56.81438, 
    56.87696, 56.93939, 57.00165, 57.06375, 57.12569, 57.18747, 57.24908, 
    57.31052, 57.3718, 57.43291, 57.49385, 57.55462, 57.61523, 57.67566, 
    57.73591, 57.79599, 57.8559, 57.91563, 57.97519, 58.03457, 58.09377, 
    58.15279, 58.21162, 58.27028, 58.32875, 58.38704, 58.44514, 58.50306, 
    58.56079, 58.61833, 58.67568, 58.73284, 58.78981, 58.84659, 58.90317, 
    58.95956, 59.01575, 59.07174, 59.12753, 59.18313, 59.23852, 59.29372, 
    59.34871, 59.40349, 59.45807, 59.51244, 59.56661, 59.62057, 59.67432, 
    59.72786, 59.78118, 59.83429, 59.88719, 59.93987, 59.99233, 60.04458, 
    60.0966, 60.14841, 60.2, 60.25136, 60.30249, 60.35341, 60.40409, 
    60.45455, 60.50478, 60.55478, 60.60455, 60.65408, 60.70339, 60.75245, 
    60.80128, 60.84988, 60.89824, 60.94635, 60.99422, 61.04185, 61.08924, 
    61.13639, 61.18328, 61.22993, 61.27634, 61.32249, 61.36839, 61.41404, 
    61.45943, 61.50457, 61.54945, 61.59408, 61.63845, 61.68256, 61.72641, 
    61.76999, 61.81332, 61.85637, 61.89916, 61.94169, 61.98394, 62.02593, 
    62.06764, 62.10909, 62.15025, 62.19115, 62.23177, 62.27211, 62.31217, 
    62.35195, 62.39145, 62.43067, 62.46961, 62.50826, 62.54663, 62.58471, 
    62.62249, 62.66, 62.6972, 62.73412, 62.77074, 62.80708, 62.84311, 
    62.87885, 62.91428, 62.94942, 62.98426, 63.0188, 63.05304, 63.08696, 
    63.12059, 63.15391, 63.18692, 63.21962, 63.25201, 63.2841, 63.31586, 
    63.34732, 63.37846, 63.40929, 63.4398, 63.46999, 63.49986, 63.52941, 
    63.55864, 63.58755, 63.61613, 63.6444, 63.67233, 63.69994, 63.72722, 
    63.75417, 63.7808, 63.80709, 63.83305, 63.85868, 63.88397, 63.90893, 
    63.93356, 63.95784, 63.98179, 64.0054, 64.02867, 64.05161, 64.0742, 
    64.09644, 64.11834, 64.1399, 64.16112, 64.18198, 64.20251, 64.22269, 
    64.24251, 64.26199, 64.28111, 64.29989, 64.31831, 64.33639, 64.3541, 
    64.37148, 64.38848, 64.40514, 64.42144, 64.43738, 64.45296, 64.46819, 
    64.48306, 64.49757, 64.51172, 64.52551, 64.53894, 64.552, 64.5647, 
    64.57705, 64.58903, 64.60064, 64.61189, 64.62277, 64.63329, 64.64344, 
    64.65323, 64.66265, 64.6717, 64.68038, 64.68871, 64.69665, 64.70423, 
    64.71144, 64.71828, 64.72475, 64.73086, 64.73659, 64.74195, 64.74694, 
    64.75156, 64.75581, 64.75968, 64.76319, 64.76632, 64.76908, 64.77148, 
    64.77349, 64.77514, 64.77641, 64.77731, 64.77784, 64.778, 64.77779, 
    64.7772, 64.77624, 64.7749, 64.7732, 64.77112, 64.76867, 64.76585, 
    64.76266, 64.75909, 64.75516, 64.75085, 64.74618, 64.74113, 64.7357, 
    64.72991, 64.72375, 64.71722, 64.71033, 64.70306, 64.69542, 64.68741, 
    64.67904, 64.6703, 64.66119, 64.6517, 64.64186, 64.63165, 64.62107, 
    64.61013, 64.59882, 64.58716, 64.57512, 64.56272, 64.54996, 64.53683, 
    64.52335, 64.50951, 64.4953, 64.48074, 64.46581, 64.45052, 64.43488, 
    64.41888, 64.40253, 64.38582, 64.36875, 64.35133, 64.33355, 64.31542, 
    64.29694, 64.27811, 64.25893, 64.2394, 64.21951, 64.19929, 64.17871, 
    64.15778, 64.13651, 64.1149, 64.09294, 64.07064, 64.048, 64.02502, 
    64.00169, 63.97802, 63.95402, 63.92968, 63.90501, 63.87999, 63.85464, 
    63.82896, 63.80295, 63.77661, 63.74993, 63.72293, 63.69559, 63.66793, 
    63.63995, 63.61164, 63.583, 63.55404, 63.52476, 63.49516, 63.46523, 
    63.43499, 63.40443, 63.37356, 63.34237, 63.31086, 63.27904, 63.24691, 
    63.21447, 63.18172, 63.14866, 63.11529, 63.08162, 63.04764, 63.01336, 
    62.97877, 62.94389, 62.9087, 62.87321, 62.83743, 62.80135, 62.76497, 
    62.7283, 62.69134, 62.65408, 62.61654, 62.5787, 62.54058, 62.50217, 
    62.46347, 62.42449, 62.38522, 62.34568, 62.30585, 62.26574, 62.22536, 
    62.1847, 62.14376, 62.10255, 62.06106, 62.01931, 61.97728, 61.93498, 
    61.89241, 61.84958, 61.80648, 61.76311, 61.71949, 61.6756, 61.63145, 
    61.58704, 61.54237, 61.49745, 61.45227, 61.40683, 61.36115, 61.3152, 
    61.26901, 61.22257, 61.17588, 61.12894, 61.08176, 61.03434, 60.98667, 
    60.93876, 60.8906, 60.84221, 60.79358, 60.74471, 60.6956, 60.64626, 
    60.59669, 60.54689, 60.49685, 60.44659, 60.39609, 60.34537, 60.29442, 
    60.24325, 60.19185, 60.14023, 60.08839, 60.03633, 59.98405, 59.93155, 
    59.87883, 59.8259,
  54.20632, 54.2748, 54.34315, 54.41138, 54.47948, 54.54745, 54.6153, 
    54.68302, 54.75061, 54.81808, 54.88541, 54.95261, 55.01968, 55.08661, 
    55.15341, 55.22008, 55.28661, 55.35301, 55.41927, 55.48539, 55.55136, 
    55.61721, 55.68291, 55.74847, 55.81389, 55.87916, 55.94429, 56.00928, 
    56.07412, 56.13881, 56.20336, 56.26775, 56.332, 56.3961, 56.46005, 
    56.52384, 56.58748, 56.65097, 56.7143, 56.77748, 56.8405, 56.90336, 
    56.96606, 57.02861, 57.09099, 57.15321, 57.21527, 57.27717, 57.3389, 
    57.40047, 57.46186, 57.5231, 57.58416, 57.64505, 57.70578, 57.76633, 
    57.82671, 57.88691, 57.94695, 58.0068, 58.06648, 58.12598, 58.1853, 
    58.24445, 58.30341, 58.36219, 58.42078, 58.47919, 58.53742, 58.59546, 
    58.65332, 58.71098, 58.76846, 58.82574, 58.88284, 58.93974, 58.99645, 
    59.05296, 59.10928, 59.1654, 59.22132, 59.27704, 59.33256, 59.38788, 
    59.44299, 59.49791, 59.55261, 59.60711, 59.66141, 59.71549, 59.76937, 
    59.82303, 59.87648, 59.92972, 59.98274, 60.03555, 60.08814, 60.14051, 
    60.19267, 60.2446, 60.29631, 60.3478, 60.39906, 60.4501, 60.50092, 
    60.5515, 60.60186, 60.65198, 60.70188, 60.75154, 60.80097, 60.85016, 
    60.89912, 60.94784, 60.99632, 61.04456, 61.09256, 61.14032, 61.18783, 
    61.2351, 61.28212, 61.32889, 61.37542, 61.4217, 61.46772, 61.51349, 
    61.55901, 61.60427, 61.64928, 61.69403, 61.73852, 61.78275, 61.82672, 
    61.87043, 61.91387, 61.95705, 61.99996, 62.04261, 62.08498, 62.12709, 
    62.16892, 62.21048, 62.25177, 62.29278, 62.33352, 62.37397, 62.41415, 
    62.45405, 62.49367, 62.533, 62.57206, 62.61082, 62.6493, 62.6875, 
    62.7254, 62.76301, 62.80033, 62.83736, 62.8741, 62.91053, 62.94668, 
    62.98252, 63.01807, 63.05332, 63.08827, 63.12291, 63.15725, 63.19129, 
    63.22502, 63.25844, 63.29156, 63.32436, 63.35686, 63.38904, 63.42091, 
    63.45247, 63.48371, 63.51463, 63.54524, 63.57552, 63.6055, 63.63514, 
    63.66447, 63.69347, 63.72215, 63.7505, 63.77853, 63.80623, 63.8336, 
    63.86064, 63.88735, 63.91373, 63.93978, 63.96549, 63.99087, 64.01591, 
    64.04062, 64.06499, 64.08901, 64.1127, 64.13605, 64.15907, 64.18172, 
    64.20405, 64.22603, 64.24767, 64.26895, 64.28989, 64.31049, 64.33073, 
    64.35062, 64.37016, 64.38936, 64.4082, 64.42669, 64.44482, 64.4626, 
    64.48003, 64.4971, 64.51382, 64.53017, 64.54617, 64.56181, 64.57709, 
    64.59201, 64.60658, 64.62077, 64.63461, 64.64809, 64.66119, 64.67394, 
    64.68633, 64.69835, 64.71001, 64.72129, 64.73222, 64.74277, 64.75296, 
    64.76278, 64.77223, 64.78132, 64.79003, 64.79838, 64.80636, 64.81396, 
    64.8212, 64.82806, 64.83456, 64.84068, 64.84644, 64.85182, 64.85683, 
    64.86147, 64.86572, 64.86961, 64.87314, 64.87628, 64.87905, 64.88145, 
    64.88348, 64.88512, 64.88641, 64.88731, 64.88784, 64.888, 64.88778, 
    64.88719, 64.88623, 64.88489, 64.88318, 64.8811, 64.87864, 64.87581, 
    64.8726, 64.86903, 64.86507, 64.86076, 64.85606, 64.85099, 64.84555, 
    64.83974, 64.83356, 64.827, 64.82008, 64.81278, 64.80512, 64.79709, 
    64.78868, 64.77991, 64.77076, 64.76125, 64.75137, 64.74113, 64.73051, 
    64.71953, 64.70818, 64.69647, 64.68439, 64.67195, 64.65915, 64.64597, 
    64.63245, 64.61855, 64.60429, 64.58968, 64.5747, 64.55936, 64.54366, 
    64.52761, 64.51119, 64.49442, 64.47729, 64.45982, 64.44198, 64.42379, 
    64.40524, 64.38634, 64.3671, 64.3475, 64.32755, 64.30725, 64.2866, 
    64.2656, 64.24426, 64.22257, 64.20055, 64.17817, 64.15545, 64.13239, 
    64.10898, 64.08524, 64.06115, 64.03673, 64.01197, 63.98687, 63.96144, 
    63.93568, 63.90958, 63.88315, 63.85638, 63.82929, 63.80187, 63.77412, 
    63.74604, 63.71763, 63.6889, 63.65985, 63.63047, 63.60077, 63.57076, 
    63.54042, 63.50976, 63.47879, 63.44749, 63.41589, 63.38397, 63.35174, 
    63.31919, 63.28634, 63.25317, 63.2197, 63.18592, 63.15184, 63.11745, 
    63.08276, 63.04776, 63.01247, 62.97688, 62.94098, 62.90479, 62.86831, 
    62.83152, 62.79445, 62.75708, 62.71942, 62.68147, 62.64323, 62.60471, 
    62.5659, 62.5268, 62.48742, 62.44776, 62.40782, 62.3676, 62.32709, 
    62.28631, 62.24525, 62.20393, 62.16232, 62.12045, 62.0783, 62.03588, 
    61.99319, 61.95024, 61.90702, 61.86353, 61.81978, 61.77577, 61.7315, 
    61.68697, 61.64218, 61.59713, 61.55183, 61.50627, 61.46046, 61.41439, 
    61.36808, 61.32151, 61.2747, 61.22763, 61.18033, 61.13278, 61.08498, 
    61.03695, 60.98867, 60.94015, 60.89139, 60.8424, 60.79316, 60.7437, 
    60.694, 60.64407, 60.59391, 60.54351, 60.49289, 60.44204, 60.39097, 
    60.33967, 60.28815, 60.2364, 60.18443, 60.13224, 60.07984, 60.02721, 
    59.97437, 59.92131,
  54.29055, 54.35913, 54.42759, 54.49593, 54.56414, 54.63222, 54.70018, 
    54.76801, 54.8357, 54.90328, 54.97072, 55.03803, 55.10521, 55.17225, 
    55.23917, 55.30595, 55.37259, 55.43909, 55.50547, 55.5717, 55.63779, 
    55.70375, 55.76957, 55.83524, 55.90077, 55.96616, 56.03141, 56.09651, 
    56.16146, 56.22627, 56.29093, 56.35545, 56.41981, 56.48403, 56.54809, 
    56.612, 56.67576, 56.73937, 56.80282, 56.86611, 56.92925, 56.99223, 
    57.05506, 57.11772, 57.18022, 57.24257, 57.30474, 57.36676, 57.42861, 
    57.4903, 57.55182, 57.61317, 57.67436, 57.73537, 57.79622, 57.8569, 
    57.9174, 57.97773, 58.03788, 58.09786, 58.15766, 58.21729, 58.27673, 
    58.336, 58.39508, 58.45399, 58.51271, 58.57125, 58.6296, 58.68777, 
    58.74574, 58.80354, 58.86114, 58.91855, 58.97577, 59.03279, 59.08963, 
    59.14627, 59.20271, 59.25896, 59.315, 59.37085, 59.4265, 59.48195, 
    59.53719, 59.59223, 59.64706, 59.70169, 59.75611, 59.81032, 59.86432, 
    59.91811, 59.97169, 60.02505, 60.07821, 60.13114, 60.18386, 60.23636, 
    60.28864, 60.3407, 60.39254, 60.44416, 60.49555, 60.54671, 60.59766, 
    60.64837, 60.69885, 60.7491, 60.79913, 60.84891, 60.89847, 60.94779, 
    60.99687, 61.04572, 61.09432, 61.14269, 61.19081, 61.2387, 61.28634, 
    61.33373, 61.38088, 61.42778, 61.47443, 61.52083, 61.56698, 61.61288, 
    61.65852, 61.7039, 61.74903, 61.79391, 61.83852, 61.88288, 61.92697, 
    61.9708, 62.01436, 62.05766, 62.1007, 62.14346, 62.18596, 62.22818, 
    62.27014, 62.31182, 62.35323, 62.39436, 62.43521, 62.47578, 62.51608, 
    62.5561, 62.59583, 62.63528, 62.67445, 62.71333, 62.75193, 62.79023, 
    62.82825, 62.86597, 62.90341, 62.94055, 62.9774, 63.01395, 63.05021, 
    63.08616, 63.12182, 63.15717, 63.19223, 63.22698, 63.26143, 63.29557, 
    63.32941, 63.36293, 63.39615, 63.42906, 63.46166, 63.49395, 63.52592, 
    63.55758, 63.58891, 63.61994, 63.65064, 63.68103, 63.71109, 63.74084, 
    63.77026, 63.79936, 63.82813, 63.85658, 63.88469, 63.91248, 63.93995, 
    63.96708, 63.99388, 64.02034, 64.04648, 64.07227, 64.09774, 64.12286, 
    64.14765, 64.1721, 64.19621, 64.21999, 64.24342, 64.2665, 64.28925, 
    64.31165, 64.33369, 64.35541, 64.37676, 64.39777, 64.41844, 64.43875, 
    64.45872, 64.47833, 64.49759, 64.51649, 64.53505, 64.55325, 64.57109, 
    64.58858, 64.60571, 64.62248, 64.63889, 64.65495, 64.67065, 64.68598, 
    64.70095, 64.71556, 64.72981, 64.7437, 64.75723, 64.77038, 64.78317, 
    64.7956, 64.80766, 64.81936, 64.83069, 64.84165, 64.85225, 64.86247, 
    64.87233, 64.88181, 64.89093, 64.89968, 64.90806, 64.91606, 64.9237, 
    64.93096, 64.93785, 64.94437, 64.95052, 64.95629, 64.96169, 64.96671, 
    64.97137, 64.97565, 64.97955, 64.98308, 64.98624, 64.98902, 64.99142, 
    64.99346, 64.99512, 64.9964, 64.99731, 64.99784, 64.998, 64.99778, 
    64.99719, 64.99622, 64.99488, 64.99316, 64.99107, 64.9886, 64.98576, 
    64.98254, 64.97896, 64.97499, 64.97066, 64.96594, 64.96086, 64.9554, 
    64.94957, 64.94336, 64.93678, 64.92983, 64.92252, 64.91482, 64.90675, 
    64.89832, 64.88952, 64.88034, 64.8708, 64.86088, 64.85059, 64.83994, 
    64.82893, 64.81754, 64.80579, 64.79366, 64.78117, 64.76833, 64.7551, 
    64.74152, 64.72758, 64.71328, 64.69861, 64.68358, 64.66818, 64.65244, 
    64.63632, 64.61985, 64.60302, 64.58583, 64.56829, 64.55039, 64.53214, 
    64.51353, 64.49457, 64.47525, 64.45558, 64.43556, 64.41519, 64.39448, 
    64.37341, 64.35199, 64.33023, 64.30812, 64.28567, 64.26287, 64.23973, 
    64.21625, 64.19242, 64.16826, 64.14375, 64.11891, 64.09373, 64.06821, 
    64.04237, 64.01618, 63.98966, 63.96281, 63.93562, 63.90811, 63.88027, 
    63.8521, 63.8236, 63.79478, 63.76563, 63.73616, 63.70636, 63.67624, 
    63.64581, 63.61505, 63.58398, 63.55259, 63.52088, 63.48886, 63.45652, 
    63.42388, 63.39092, 63.35765, 63.32407, 63.29019, 63.256, 63.2215, 
    63.1867, 63.1516, 63.1162, 63.08049, 63.04449, 63.00819, 62.97159, 
    62.9347, 62.89751, 62.86003, 62.82225, 62.78419, 62.74584, 62.7072, 
    62.66827, 62.62906, 62.58957, 62.54979, 62.50973, 62.46939, 62.42876, 
    62.38787, 62.34669, 62.30524, 62.26352, 62.22152, 62.17925, 62.13671, 
    62.09391, 62.05083, 62.00749, 61.96388, 61.92001, 61.87588, 61.83148, 
    61.78683, 61.74191, 61.69674, 61.65131, 61.60563, 61.5597, 61.51351, 
    61.46707, 61.42038, 61.37344, 61.32625, 61.27882, 61.23114, 61.18322, 
    61.13506, 61.08665, 61.03801, 60.98912, 60.94, 60.89064, 60.84105, 
    60.79123, 60.74117, 60.69088, 60.64036, 60.58961, 60.53864, 60.48743, 
    60.43601, 60.38436, 60.33248, 60.28039, 60.22807, 60.17554, 60.12278, 
    60.06981, 60.01663,
  54.37465, 54.44334, 54.51191, 54.58035, 54.64867, 54.71686, 54.78493, 
    54.85287, 54.92068, 54.98836, 55.05591, 55.12333, 55.19062, 55.25778, 
    55.3248, 55.39169, 55.45845, 55.52507, 55.59155, 55.6579, 55.72411, 
    55.79017, 55.8561, 55.92189, 55.98754, 56.05304, 56.1184, 56.18362, 
    56.24869, 56.31361, 56.37839, 56.44302, 56.5075, 56.57184, 56.63602, 
    56.70005, 56.76392, 56.82765, 56.89122, 56.95463, 57.01789, 57.08099, 
    57.14394, 57.20672, 57.26934, 57.3318, 57.3941, 57.45624, 57.51822, 
    57.58002, 57.64167, 57.70314, 57.76445, 57.82558, 57.88655, 57.94735, 
    58.00798, 58.06843, 58.1287, 58.18881, 58.24873, 58.30848, 58.36805, 
    58.42744, 58.48666, 58.54568, 58.60453, 58.66319, 58.72167, 58.77996, 
    58.83807, 58.89598, 58.95371, 59.01125, 59.0686, 59.12575, 59.18271, 
    59.23948, 59.29605, 59.35242, 59.40859, 59.46457, 59.52034, 59.57592, 
    59.63129, 59.68645, 59.74141, 59.79617, 59.85072, 59.90506, 59.95918, 
    60.0131, 60.06681, 60.1203, 60.17358, 60.22665, 60.27949, 60.33212, 
    60.38453, 60.43672, 60.48868, 60.54043, 60.59195, 60.64324, 60.69431, 
    60.74515, 60.79576, 60.84614, 60.89629, 60.94621, 60.99589, 61.04533, 
    61.09454, 61.14352, 61.19225, 61.24075, 61.289, 61.33701, 61.38477, 
    61.43229, 61.47956, 61.52659, 61.57336, 61.61989, 61.66616, 61.71219, 
    61.75795, 61.80347, 61.84872, 61.89372, 61.93846, 61.98293, 62.02715, 
    62.0711, 62.11479, 62.15821, 62.20137, 62.24425, 62.28687, 62.32922, 
    62.37129, 62.41309, 62.45462, 62.49587, 62.53684, 62.57754, 62.61795, 
    62.65809, 62.69794, 62.73751, 62.77679, 62.81579, 62.8545, 62.89292, 
    62.93105, 62.96889, 63.00644, 63.04369, 63.08065, 63.11731, 63.15368, 
    63.18975, 63.22551, 63.26098, 63.29614, 63.33101, 63.36556, 63.39981, 
    63.43375, 63.46738, 63.50071, 63.53372, 63.56643, 63.59881, 63.63089, 
    63.66264, 63.69408, 63.72521, 63.75602, 63.7865, 63.81666, 63.8465, 
    63.87602, 63.90521, 63.93408, 63.96262, 63.99083, 64.01871, 64.04626, 
    64.07349, 64.10037, 64.12693, 64.15315, 64.17904, 64.20458, 64.2298, 
    64.25467, 64.27921, 64.3034, 64.32725, 64.35075, 64.37392, 64.39674, 
    64.41922, 64.44135, 64.46313, 64.48456, 64.50565, 64.52638, 64.54677, 
    64.5668, 64.58648, 64.6058, 64.62478, 64.64339, 64.66166, 64.67957, 
    64.69711, 64.7143, 64.73113, 64.7476, 64.76372, 64.77946, 64.79485, 
    64.80988, 64.82455, 64.83884, 64.85278, 64.86636, 64.87956, 64.8924, 
    64.90487, 64.91698, 64.92872, 64.94009, 64.95109, 64.96172, 64.97198, 
    64.98187, 64.99139, 65.00054, 65.00932, 65.01773, 65.02576, 65.03342, 
    65.04072, 65.04763, 65.05418, 65.06034, 65.06614, 65.07156, 65.0766, 
    65.08127, 65.08556, 65.08949, 65.09303, 65.09619, 65.09898, 65.1014, 
    65.10344, 65.10511, 65.10639, 65.10731, 65.10784, 65.108, 65.10778, 
    65.10719, 65.10622, 65.10487, 65.10314, 65.10104, 65.09857, 65.09572, 
    65.09249, 65.08889, 65.08491, 65.08056, 65.07583, 65.07072, 65.06525, 
    65.05939, 65.05316, 65.04656, 65.03959, 65.03224, 65.02452, 65.01643, 
    65.00796, 64.99912, 64.98991, 64.98033, 64.97038, 64.96006, 64.94937, 
    64.93832, 64.92689, 64.91508, 64.90292, 64.8904, 64.87749, 64.86423, 
    64.8506, 64.83661, 64.82225, 64.80753, 64.79245, 64.777, 64.76119, 
    64.74503, 64.72849, 64.71161, 64.69436, 64.67676, 64.65879, 64.64047, 
    64.6218, 64.60278, 64.58339, 64.56365, 64.54356, 64.52312, 64.50233, 
    64.48119, 64.45971, 64.43787, 64.41569, 64.39316, 64.37028, 64.34706, 
    64.32349, 64.29959, 64.27534, 64.25076, 64.22583, 64.20057, 64.17496, 
    64.14902, 64.12275, 64.09615, 64.06921, 64.04193, 64.01433, 63.98639, 
    63.95813, 63.92953, 63.90062, 63.87137, 63.8418, 63.81191, 63.7817, 
    63.75116, 63.72031, 63.68913, 63.65764, 63.62584, 63.59371, 63.56127, 
    63.52852, 63.49546, 63.46209, 63.4284, 63.39441, 63.36012, 63.32551, 
    63.2906, 63.25539, 63.21988, 63.18406, 63.14795, 63.11153, 63.07483, 
    63.03782, 63.00052, 62.96292, 62.92504, 62.88686, 62.84839, 62.80964, 
    62.7706, 62.73127, 62.69165, 62.65176, 62.61158, 62.57112, 62.53038, 
    62.48936, 62.44807, 62.4065, 62.36465, 62.32254, 62.28015, 62.23749, 
    62.19456, 62.15136, 62.10789, 62.06417, 62.02017, 61.97591, 61.9314, 
    61.88662, 61.84158, 61.79628, 61.75073, 61.70493, 61.65886, 61.61255, 
    61.56598, 61.51917, 61.4721, 61.42479, 61.37723, 61.32943, 61.28138, 
    61.23309, 61.18456, 61.13578, 61.08678, 61.03753, 60.98804, 60.93832, 
    60.88837, 60.83818, 60.78777, 60.73712, 60.68624, 60.63514, 60.58381, 
    60.53226, 60.48048, 60.42847, 60.37625, 60.32381, 60.27114, 60.21827, 
    60.16517, 60.11185,
  54.45863, 54.52743, 54.59611, 54.66466, 54.73308, 54.80138, 54.86956, 
    54.93761, 55.00553, 55.07332, 55.14098, 55.20851, 55.27591, 55.34318, 
    55.41032, 55.47732, 55.54419, 55.61092, 55.67751, 55.74397, 55.8103, 
    55.87648, 55.94252, 56.00842, 56.07418, 56.1398, 56.20528, 56.27061, 
    56.3358, 56.40084, 56.46574, 56.53048, 56.59508, 56.65953, 56.72383, 
    56.78798, 56.85197, 56.91582, 56.9795, 57.04304, 57.10641, 57.16964, 
    57.2327, 57.2956, 57.35835, 57.42093, 57.48335, 57.54561, 57.6077, 
    57.66964, 57.7314, 57.793, 57.85443, 57.91569, 57.97678, 58.0377, 
    58.09845, 58.15902, 58.21943, 58.27965, 58.3397, 58.39957, 58.45927, 
    58.51879, 58.57812, 58.63728, 58.69625, 58.75504, 58.81364, 58.87206, 
    58.93029, 58.98833, 59.04619, 59.10385, 59.16132, 59.21861, 59.27569, 
    59.33258, 59.38928, 59.44578, 59.50208, 59.55819, 59.61409, 59.66979, 
    59.72528, 59.78058, 59.83567, 59.89055, 59.94523, 59.99969, 60.05396, 
    60.108, 60.16183, 60.21546, 60.26886, 60.32206, 60.37503, 60.42779, 
    60.48032, 60.53264, 60.58474, 60.63661, 60.68826, 60.73968, 60.79087, 
    60.84184, 60.89258, 60.94309, 60.99337, 61.04341, 61.09322, 61.1428, 
    61.19213, 61.24124, 61.2901, 61.33872, 61.3871, 61.43523, 61.48313, 
    61.53077, 61.57817, 61.62532, 61.67223, 61.71888, 61.76528, 61.81143, 
    61.85732, 61.90296, 61.94834, 61.99346, 62.03832, 62.08292, 62.12726, 
    62.17134, 62.21515, 62.25869, 62.30197, 62.34498, 62.38772, 62.43019, 
    62.47239, 62.51431, 62.55595, 62.59732, 62.63842, 62.67923, 62.71976, 
    62.76002, 62.79999, 62.83967, 62.87907, 62.91819, 62.95701, 62.99555, 
    63.0338, 63.07175, 63.10941, 63.14678, 63.18385, 63.22063, 63.25711, 
    63.29329, 63.32917, 63.36474, 63.40001, 63.43498, 63.46965, 63.50401, 
    63.53806, 63.5718, 63.60522, 63.63834, 63.67115, 63.70364, 63.73582, 
    63.76768, 63.79922, 63.83044, 63.86135, 63.89193, 63.9222, 63.95213, 
    63.98175, 64.01104, 64.04, 64.06863, 64.09694, 64.12491, 64.15256, 
    64.17987, 64.20685, 64.23349, 64.2598, 64.28577, 64.31141, 64.33671, 
    64.36166, 64.38628, 64.41055, 64.43449, 64.45808, 64.48132, 64.50422, 
    64.52677, 64.54897, 64.57083, 64.59234, 64.6135, 64.63431, 64.65476, 
    64.67487, 64.69461, 64.714, 64.73305, 64.75173, 64.77006, 64.78802, 
    64.80563, 64.82288, 64.83978, 64.85631, 64.87247, 64.88828, 64.90372, 
    64.91881, 64.93353, 64.94788, 64.96186, 64.97548, 64.98873, 65.00162, 
    65.01414, 65.02628, 65.03806, 65.04948, 65.06052, 65.07119, 65.08149, 
    65.09142, 65.10097, 65.11015, 65.11897, 65.1274, 65.13547, 65.14316, 
    65.15047, 65.15741, 65.16398, 65.17017, 65.17598, 65.18142, 65.18649, 
    65.19117, 65.19548, 65.19942, 65.20297, 65.20615, 65.20895, 65.21138, 
    65.21342, 65.2151, 65.21638, 65.2173, 65.21784, 65.218, 65.21778, 
    65.21719, 65.21621, 65.21486, 65.21313, 65.21102, 65.20853, 65.20567, 
    65.20244, 65.19882, 65.19482, 65.19045, 65.18571, 65.18059, 65.17509, 
    65.16921, 65.16296, 65.15634, 65.14934, 65.14196, 65.13422, 65.12609, 
    65.11759, 65.10873, 65.09948, 65.08987, 65.07988, 65.06953, 65.05879, 
    65.0477, 65.03622, 65.02439, 65.01218, 64.9996, 64.98666, 64.97335, 
    64.95967, 64.94563, 64.93122, 64.91644, 64.90131, 64.8858, 64.86994, 
    64.85371, 64.83713, 64.82018, 64.80287, 64.78521, 64.76718, 64.74879, 
    64.73006, 64.71096, 64.69151, 64.67171, 64.65155, 64.63104, 64.61018, 
    64.58897, 64.5674, 64.54549, 64.52322, 64.50062, 64.47767, 64.45437, 
    64.43073, 64.40674, 64.38241, 64.35773, 64.33273, 64.30737, 64.28168, 
    64.25566, 64.2293, 64.2026, 64.17557, 64.14821, 64.12051, 64.09248, 
    64.06413, 64.03544, 64.00642, 63.97709, 63.94742, 63.91743, 63.88712, 
    63.85648, 63.82553, 63.79425, 63.76266, 63.73075, 63.69852, 63.66598, 
    63.63313, 63.59996, 63.56648, 63.53269, 63.49859, 63.46418, 63.42947, 
    63.39445, 63.35913, 63.32351, 63.28758, 63.25136, 63.21483, 63.17801, 
    63.14089, 63.10348, 63.06577, 63.02777, 62.98948, 62.95089, 62.91202, 
    62.87286, 62.83342, 62.79368, 62.75367, 62.71337, 62.67279, 62.63194, 
    62.5908, 62.54939, 62.50769, 62.46573, 62.42349, 62.38098, 62.3382, 
    62.29514, 62.25182, 62.20824, 62.16438, 62.12027, 62.07588, 62.03124, 
    61.98634, 61.94117, 61.89576, 61.85007, 61.80414, 61.75796, 61.71152, 
    61.66483, 61.61788, 61.57069, 61.52325, 61.47557, 61.42764, 61.37946, 
    61.33104, 61.28238, 61.23349, 61.18435, 61.13497, 61.08536, 61.03551, 
    60.98543, 60.93512, 60.88457, 60.8338, 60.78279, 60.73156, 60.6801, 
    60.62842, 60.57651, 60.52438, 60.47203, 60.41946, 60.36666, 60.31366, 
    60.26043, 60.20699,
  54.54249, 54.6114, 54.68018, 54.74884, 54.81738, 54.88578, 54.95407, 
    55.02222, 55.09026, 55.15815, 55.22593, 55.29357, 55.36108, 55.42846, 
    55.49571, 55.56282, 55.6298, 55.69665, 55.76336, 55.82993, 55.89637, 
    55.96266, 56.02882, 56.09484, 56.16071, 56.22645, 56.29204, 56.35749, 
    56.42279, 56.48795, 56.55296, 56.61782, 56.68254, 56.74711, 56.81153, 
    56.87579, 56.93991, 57.00387, 57.06768, 57.13133, 57.19482, 57.25817, 
    57.32135, 57.38437, 57.44724, 57.50994, 57.57249, 57.63486, 57.69708, 
    57.75914, 57.82102, 57.88274, 57.94429, 58.00568, 58.06689, 58.12794, 
    58.18881, 58.24951, 58.31004, 58.37038, 58.43056, 58.49056, 58.55038, 
    58.61002, 58.66948, 58.72876, 58.78786, 58.84677, 58.9055, 58.96405, 
    59.0224, 59.08057, 59.13856, 59.19635, 59.25395, 59.31136, 59.36857, 
    59.42559, 59.48241, 59.53904, 59.59547, 59.6517, 59.70773, 59.76356, 
    59.81919, 59.87461, 59.92983, 59.98484, 60.03965, 60.09424, 60.14863, 
    60.2028, 60.25677, 60.31052, 60.36406, 60.41737, 60.47048, 60.52337, 
    60.57603, 60.62848, 60.6807, 60.7327, 60.78448, 60.83603, 60.88736, 
    60.93845, 60.98932, 61.03996, 61.09036, 61.14054, 61.19048, 61.24018, 
    61.28965, 61.33887, 61.38786, 61.43661, 61.48512, 61.53338, 61.5814, 
    61.62918, 61.6767, 61.72398, 61.77101, 61.81779, 61.86432, 61.91059, 
    61.95661, 62.00237, 62.04788, 62.09313, 62.13811, 62.18284, 62.2273, 
    62.2715, 62.31544, 62.35911, 62.40251, 62.44564, 62.4885, 62.53109, 
    62.57341, 62.61546, 62.65722, 62.69872, 62.73993, 62.78086, 62.82152, 
    62.86189, 62.90198, 62.94178, 62.9813, 63.02053, 63.05947, 63.09813, 
    63.13649, 63.17456, 63.21234, 63.24982, 63.28701, 63.3239, 63.36049, 
    63.39678, 63.43277, 63.46846, 63.50384, 63.53892, 63.57369, 63.60816, 
    63.64231, 63.67616, 63.7097, 63.74292, 63.77583, 63.80843, 63.84071, 
    63.87267, 63.90432, 63.93565, 63.96665, 63.99733, 64.02769, 64.05773, 
    64.08744, 64.11683, 64.14588, 64.17461, 64.20301, 64.23108, 64.25882, 
    64.28622, 64.31329, 64.34003, 64.36642, 64.39249, 64.41821, 64.44359, 
    64.46863, 64.49333, 64.51768, 64.5417, 64.56538, 64.5887, 64.61168, 
    64.63431, 64.65659, 64.67852, 64.7001, 64.72134, 64.74222, 64.76274, 
    64.78291, 64.80273, 64.8222, 64.8413, 64.86005, 64.87844, 64.89648, 
    64.91415, 64.93146, 64.94841, 64.965, 64.98122, 64.99709, 65.01259, 
    65.02772, 65.04249, 65.05689, 65.07093, 65.08459, 65.0979, 65.11083, 
    65.12339, 65.13559, 65.14741, 65.15886, 65.16994, 65.18065, 65.19099, 
    65.20095, 65.21054, 65.21976, 65.2286, 65.23707, 65.24516, 65.25288, 
    65.26022, 65.26719, 65.27378, 65.27999, 65.28583, 65.29129, 65.29637, 
    65.30107, 65.3054, 65.30935, 65.31292, 65.31611, 65.31892, 65.32136, 
    65.32341, 65.32509, 65.32639, 65.3273, 65.32784, 65.328, 65.32778, 
    65.32718, 65.3262, 65.32484, 65.32311, 65.32099, 65.3185, 65.31563, 
    65.31238, 65.30875, 65.30474, 65.30035, 65.29559, 65.29045, 65.28493, 
    65.27904, 65.27276, 65.26611, 65.25909, 65.25169, 65.2439, 65.23576, 
    65.22723, 65.21832, 65.20905, 65.1994, 65.18938, 65.17898, 65.16821, 
    65.15707, 65.14556, 65.13368, 65.12143, 65.10881, 65.09582, 65.08246, 
    65.06873, 65.05464, 65.04018, 65.02535, 65.01016, 64.99461, 64.97868, 
    64.96239, 64.94576, 64.92874, 64.91138, 64.89365, 64.87556, 64.85711, 
    64.8383, 64.81914, 64.79962, 64.77975, 64.75952, 64.73894, 64.718, 
    64.69672, 64.67507, 64.65308, 64.63075, 64.60806, 64.58503, 64.56165, 
    64.53793, 64.51385, 64.48945, 64.46469, 64.4396, 64.41416, 64.38838, 
    64.36227, 64.33582, 64.30903, 64.28191, 64.25446, 64.22666, 64.19854, 
    64.17009, 64.14131, 64.1122, 64.08276, 64.053, 64.02291, 63.9925, 
    63.96177, 63.93071, 63.89933, 63.86764, 63.83562, 63.8033, 63.77065, 
    63.73769, 63.70441, 63.67083, 63.63693, 63.60273, 63.56821, 63.53339, 
    63.49826, 63.46283, 63.4271, 63.39106, 63.35472, 63.31808, 63.28115, 
    63.24391, 63.20638, 63.16856, 63.13044, 63.09203, 63.05334, 63.01435, 
    62.97507, 62.9355, 62.89566, 62.85552, 62.81511, 62.77441, 62.73343, 
    62.69217, 62.65063, 62.60883, 62.56674, 62.52438, 62.48174, 62.43884, 
    62.39566, 62.35222, 62.30851, 62.26453, 62.22029, 62.17578, 62.13102, 
    62.08599, 62.0407, 61.99515, 61.94935, 61.90329, 61.85698, 61.81041, 
    61.76359, 61.71652, 61.6692, 61.62164, 61.57382, 61.52576, 61.47746, 
    61.42892, 61.38013, 61.3311, 61.28184, 61.23233, 61.18259, 61.13261, 
    61.08241, 61.03196, 60.98129, 60.93039, 60.87925, 60.82789, 60.7763, 
    60.72449, 60.67245, 60.6202, 60.56771, 60.51501, 60.46209, 60.40895, 
    60.3556, 60.30203,
  54.62622, 54.69524, 54.76413, 54.8329, 54.90154, 54.97006, 55.03845, 
    55.10672, 55.17486, 55.24287, 55.31075, 55.37851, 55.44613, 55.51362, 
    55.58098, 55.6482, 55.7153, 55.78226, 55.84908, 55.91576, 55.98231, 
    56.04873, 56.115, 56.18113, 56.24712, 56.31297, 56.37868, 56.44424, 
    56.50966, 56.57494, 56.64006, 56.70505, 56.76988, 56.83457, 56.8991, 
    56.96349, 57.02772, 57.0918, 57.15573, 57.2195, 57.28312, 57.34658, 
    57.40988, 57.47303, 57.53601, 57.59884, 57.6615, 57.72401, 57.78635, 
    57.84852, 57.91053, 57.97237, 58.03405, 58.09556, 58.15689, 58.21806, 
    58.27906, 58.33988, 58.40053, 58.46101, 58.52131, 58.58143, 58.64138, 
    58.70115, 58.76073, 58.82014, 58.87936, 58.9384, 58.99726, 59.05593, 
    59.11441, 59.17271, 59.23082, 59.28874, 59.34647, 59.404, 59.46135, 
    59.51849, 59.57545, 59.6322, 59.68876, 59.74512, 59.80128, 59.85724, 
    59.91299, 59.96854, 60.02389, 60.07903, 60.13396, 60.18869, 60.24321, 
    60.29751, 60.3516, 60.40549, 60.45915, 60.5126, 60.56583, 60.61885, 
    60.67165, 60.72422, 60.77658, 60.8287, 60.88061, 60.93229, 60.98375, 
    61.03497, 61.08597, 61.13674, 61.18727, 61.23758, 61.28764, 61.33747, 
    61.38707, 61.43643, 61.48555, 61.53442, 61.58306, 61.63145, 61.6796, 
    61.7275, 61.77516, 61.82257, 61.86972, 61.91663, 61.96328, 62.00968, 
    62.05583, 62.10172, 62.14735, 62.19272, 62.23783, 62.28269, 62.32728, 
    62.3716, 62.41566, 62.45946, 62.50298, 62.54624, 62.58922, 62.63194, 
    62.67438, 62.71655, 62.75843, 62.80005, 62.84138, 62.88244, 62.92321, 
    62.9637, 63.00391, 63.04383, 63.08347, 63.12282, 63.16188, 63.20065, 
    63.23913, 63.27732, 63.31521, 63.35281, 63.39011, 63.42711, 63.46382, 
    63.50022, 63.53632, 63.57212, 63.60762, 63.64281, 63.67769, 63.71227, 
    63.74653, 63.78049, 63.81413, 63.84746, 63.88048, 63.91318, 63.94556, 
    63.97763, 64.00938, 64.04081, 64.07191, 64.1027, 64.13316, 64.16329, 
    64.1931, 64.22259, 64.25174, 64.28056, 64.30906, 64.33722, 64.36505, 
    64.39255, 64.41971, 64.44653, 64.47301, 64.49917, 64.52498, 64.55045, 
    64.57558, 64.60036, 64.6248, 64.6489, 64.67265, 64.69605, 64.71911, 
    64.74182, 64.76418, 64.78619, 64.80785, 64.82915, 64.85011, 64.8707, 
    64.89095, 64.91084, 64.93037, 64.94954, 64.96835, 64.98682, 65.00491, 
    65.02264, 65.04002, 65.05703, 65.07368, 65.08997, 65.10588, 65.12144, 
    65.13663, 65.15145, 65.1659, 65.17999, 65.19371, 65.20705, 65.22003, 
    65.23264, 65.24488, 65.25674, 65.26824, 65.27937, 65.29011, 65.30048, 
    65.31049, 65.32011, 65.32936, 65.33823, 65.34673, 65.35486, 65.3626, 
    65.36997, 65.37697, 65.38358, 65.38982, 65.39568, 65.40115, 65.40625, 
    65.41097, 65.41531, 65.41928, 65.42286, 65.42606, 65.42889, 65.43133, 
    65.4334, 65.43507, 65.43638, 65.4373, 65.43784, 65.438, 65.43777, 
    65.43718, 65.4362, 65.43484, 65.43309, 65.43097, 65.42847, 65.42558, 
    65.42232, 65.41868, 65.41466, 65.41026, 65.40547, 65.40031, 65.39478, 
    65.38885, 65.38256, 65.37589, 65.36884, 65.3614, 65.3536, 65.34541, 
    65.33686, 65.32792, 65.31861, 65.30893, 65.29887, 65.28844, 65.27763, 
    65.26645, 65.2549, 65.24297, 65.23067, 65.21801, 65.20497, 65.19156, 
    65.17779, 65.16364, 65.14912, 65.13425, 65.119, 65.10339, 65.08741, 
    65.07107, 65.05436, 65.03729, 65.01986, 65.00207, 64.98392, 64.9654, 
    64.94653, 64.9273, 64.90771, 64.88777, 64.86747, 64.84682, 64.82581, 
    64.80444, 64.78273, 64.76067, 64.73825, 64.71548, 64.69238, 64.66891, 
    64.64511, 64.62096, 64.59646, 64.57162, 64.54644, 64.52092, 64.49506, 
    64.46885, 64.44231, 64.41544, 64.38822, 64.36067, 64.33279, 64.30457, 
    64.27602, 64.24715, 64.21794, 64.18841, 64.15855, 64.12836, 64.09785, 
    64.06702, 64.03586, 64.00438, 63.97258, 63.94046, 63.90803, 63.87527, 
    63.84221, 63.80883, 63.77514, 63.74113, 63.70682, 63.67219, 63.63726, 
    63.60202, 63.56648, 63.53063, 63.49448, 63.45803, 63.42128, 63.38423, 
    63.34688, 63.30924, 63.2713, 63.23307, 63.19454, 63.15572, 63.11662, 
    63.07722, 63.03754, 62.99757, 62.95732, 62.91678, 62.87596, 62.83486, 
    62.79348, 62.75183, 62.70989, 62.66768, 62.6252, 62.58244, 62.53941, 
    62.49611, 62.45255, 62.40871, 62.36461, 62.32024, 62.27561, 62.23072, 
    62.18556, 62.14015, 62.09447, 62.04855, 62.00236, 61.95592, 61.90923, 
    61.86228, 61.81508, 61.76764, 61.71994, 61.672, 61.62381, 61.57538, 
    61.52671, 61.47779, 61.42864, 61.37924, 61.32961, 61.27974, 61.22963, 
    61.17929, 61.12872, 61.07792, 61.02689, 60.97562, 60.92413, 60.87242, 
    60.82048, 60.76831, 60.71592, 60.66331, 60.61048, 60.55743, 60.50416, 
    60.45068, 60.39698,
  54.70984, 54.77895, 54.84795, 54.91683, 54.98558, 55.05421, 55.12271, 
    55.19109, 55.25934, 55.32746, 55.39545, 55.46332, 55.53105, 55.59865, 
    55.66613, 55.73346, 55.80067, 55.86774, 55.93468, 56.00148, 56.06814, 
    56.13467, 56.20105, 56.2673, 56.33341, 56.39937, 56.46519, 56.53088, 
    56.59641, 56.6618, 56.72705, 56.79215, 56.8571, 56.92191, 56.98656, 
    57.05106, 57.11542, 57.17962, 57.24366, 57.30756, 57.3713, 57.43488, 
    57.4983, 57.56157, 57.62468, 57.68762, 57.75041, 57.81303, 57.8755, 
    57.93779, 57.99992, 58.06189, 58.12369, 58.18532, 58.24678, 58.30807, 
    58.3692, 58.43015, 58.49092, 58.55152, 58.61195, 58.6722, 58.73227, 
    58.79216, 58.85188, 58.91141, 58.97076, 59.02993, 59.08891, 59.14771, 
    59.20632, 59.26474, 59.32298, 59.38103, 59.43888, 59.49655, 59.55402, 
    59.61129, 59.66838, 59.72526, 59.78195, 59.83844, 59.89473, 59.95081, 
    60.00669, 60.06238, 60.11786, 60.17313, 60.22819, 60.28304, 60.33769, 
    60.39212, 60.44635, 60.50036, 60.55415, 60.60773, 60.6611, 60.71424, 
    60.76717, 60.81987, 60.87236, 60.92462, 60.97666, 61.02847, 61.08005, 
    61.13141, 61.18254, 61.23343, 61.2841, 61.33453, 61.38473, 61.43469, 
    61.48442, 61.5339, 61.58315, 61.63216, 61.68092, 61.72944, 61.77772, 
    61.82575, 61.87354, 61.92107, 61.96836, 62.01539, 62.06217, 62.1087, 
    62.15497, 62.20099, 62.24675, 62.29225, 62.33749, 62.38247, 62.42718, 
    62.47163, 62.51582, 62.55973, 62.60339, 62.64677, 62.68988, 62.73272, 
    62.77528, 62.81757, 62.85958, 62.90132, 62.94277, 62.98395, 63.02485, 
    63.06546, 63.10579, 63.14583, 63.18559, 63.22506, 63.26423, 63.30312, 
    63.34172, 63.38002, 63.41803, 63.45575, 63.49316, 63.53028, 63.5671, 
    63.60361, 63.63983, 63.67574, 63.71135, 63.74665, 63.78164, 63.81633, 
    63.8507, 63.88477, 63.91852, 63.95196, 63.98508, 64.01789, 64.05038, 
    64.08255, 64.1144, 64.14594, 64.17714, 64.20802, 64.23859, 64.26882, 
    64.29873, 64.32831, 64.35756, 64.38648, 64.41507, 64.44333, 64.47125, 
    64.49884, 64.52609, 64.55301, 64.57959, 64.60583, 64.63172, 64.65728, 
    64.6825, 64.70736, 64.73189, 64.75607, 64.7799, 64.80339, 64.82653, 
    64.84931, 64.87175, 64.89384, 64.91557, 64.93695, 64.95798, 64.97865, 
    64.99897, 65.01893, 65.03853, 65.05777, 65.07665, 65.09517, 65.11333, 
    65.13113, 65.14857, 65.16564, 65.18235, 65.19869, 65.21467, 65.23028, 
    65.24552, 65.2604, 65.2749, 65.28904, 65.30281, 65.31621, 65.32923, 
    65.34189, 65.35417, 65.36608, 65.37762, 65.38878, 65.39957, 65.40997, 
    65.42001, 65.42967, 65.43896, 65.44787, 65.4564, 65.46455, 65.47233, 
    65.47972, 65.48674, 65.49338, 65.49963, 65.50552, 65.51102, 65.51614, 
    65.52087, 65.52523, 65.52921, 65.53281, 65.53602, 65.53886, 65.54131, 
    65.54337, 65.54507, 65.54637, 65.54729, 65.54784, 65.548, 65.54778, 
    65.54717, 65.54619, 65.54482, 65.54308, 65.54094, 65.53843, 65.53554, 
    65.53226, 65.5286, 65.52457, 65.52015, 65.51535, 65.51017, 65.50461, 
    65.49867, 65.49236, 65.48566, 65.47858, 65.47112, 65.46329, 65.45507, 
    65.44648, 65.43752, 65.42817, 65.41845, 65.40836, 65.39788, 65.38704, 
    65.37582, 65.36422, 65.35225, 65.33991, 65.32719, 65.31411, 65.30066, 
    65.28683, 65.27264, 65.25807, 65.24313, 65.22784, 65.21217, 65.19613, 
    65.17973, 65.16296, 65.14584, 65.12834, 65.11048, 65.09226, 65.07368, 
    65.05475, 65.03545, 65.01579, 64.99578, 64.9754, 64.95468, 64.93359, 
    64.91216, 64.89037, 64.86823, 64.84573, 64.82289, 64.7997, 64.77615, 
    64.75227, 64.72803, 64.70345, 64.67853, 64.65326, 64.62765, 64.6017, 
    64.57541, 64.54877, 64.5218, 64.4945, 64.46686, 64.43888, 64.41058, 
    64.38193, 64.35296, 64.32365, 64.29402, 64.26406, 64.23377, 64.20316, 
    64.17223, 64.14097, 64.10938, 64.07748, 64.04526, 64.01272, 63.97986, 
    63.94669, 63.9132, 63.8794, 63.84529, 63.81086, 63.77613, 63.74109, 
    63.70574, 63.67008, 63.63412, 63.59786, 63.56129, 63.52443, 63.48726, 
    63.4498, 63.41204, 63.37399, 63.33563, 63.29699, 63.25806, 63.21883, 
    63.17932, 63.13951, 63.09943, 63.05905, 63.01839, 62.97746, 62.93623, 
    62.89473, 62.85295, 62.8109, 62.76856, 62.72596, 62.68307, 62.63992, 
    62.5965, 62.55281, 62.50885, 62.46462, 62.42012, 62.37537, 62.33035, 
    62.28507, 62.23953, 62.19373, 62.14767, 62.10136, 62.05479, 62.00797, 
    61.96089, 61.91357, 61.86599, 61.81817, 61.7701, 61.72178, 61.67323, 
    61.62442, 61.57537, 61.52609, 61.47657, 61.4268, 61.3768, 61.32657, 
    61.2761, 61.2254, 61.17447, 61.1233, 61.07191, 61.02029, 60.96844, 
    60.91637, 60.86407, 60.81155, 60.75881, 60.70585, 60.65267, 60.59927, 
    60.54566, 60.49183,
  54.79332, 54.86255, 54.93165, 55.00064, 55.0695, 55.13823, 55.20684, 
    55.27533, 55.34369, 55.41192, 55.48003, 55.548, 55.61585, 55.68356, 
    55.75115, 55.8186, 55.88592, 55.9531, 56.02015, 56.08707, 56.15384, 
    56.22048, 56.28698, 56.35335, 56.41957, 56.48565, 56.55159, 56.61739, 
    56.68304, 56.74855, 56.81392, 56.87914, 56.94421, 57.00912, 57.0739, 
    57.13852, 57.203, 57.26731, 57.33148, 57.39549, 57.45935, 57.52306, 
    57.5866, 57.64999, 57.71322, 57.77629, 57.8392, 57.90194, 57.96453, 
    58.02695, 58.0892, 58.15129, 58.21322, 58.27497, 58.33656, 58.39798, 
    58.45922, 58.5203, 58.5812, 58.64192, 58.70248, 58.76285, 58.82305, 
    58.88307, 58.94291, 59.00257, 59.06205, 59.12134, 59.18045, 59.23938, 
    59.29812, 59.35667, 59.41504, 59.47321, 59.53119, 59.58899, 59.64659, 
    59.70399, 59.7612, 59.81821, 59.87503, 59.93165, 59.98807, 60.04428, 
    60.1003, 60.15611, 60.21172, 60.26712, 60.32231, 60.3773, 60.43208, 
    60.48664, 60.54099, 60.59513, 60.64906, 60.70277, 60.75627, 60.80954, 
    60.8626, 60.91544, 60.96805, 61.02044, 61.07261, 61.12455, 61.17627, 
    61.22775, 61.27901, 61.33004, 61.38084, 61.4314, 61.48173, 61.53182, 
    61.58167, 61.63129, 61.68067, 61.7298, 61.7787, 61.82735, 61.87576, 
    61.92392, 61.97183, 62.0195, 62.06691, 62.11407, 62.16098, 62.20764, 
    62.25404, 62.30019, 62.34607, 62.3917, 62.43707, 62.48217, 62.52701, 
    62.57159, 62.6159, 62.65995, 62.70372, 62.74723, 62.79046, 62.83342, 
    62.87611, 62.91853, 62.96066, 63.00252, 63.0441, 63.0854, 63.12642, 
    63.16715, 63.2076, 63.24776, 63.28764, 63.32723, 63.36653, 63.40554, 
    63.44425, 63.48267, 63.5208, 63.55863, 63.59616, 63.6334, 63.67033, 
    63.70696, 63.74329, 63.77931, 63.81503, 63.85044, 63.88555, 63.92035, 
    63.95483, 63.98901, 64.02287, 64.05641, 64.08965, 64.12256, 64.15515, 
    64.18743, 64.21938, 64.25101, 64.28233, 64.31332, 64.34398, 64.37431, 
    64.40433, 64.43401, 64.46336, 64.49237, 64.52106, 64.54941, 64.57742, 
    64.60511, 64.63245, 64.65946, 64.68613, 64.71246, 64.73844, 64.76408, 
    64.78939, 64.81435, 64.83895, 64.86322, 64.88714, 64.91071, 64.93392, 
    64.95679, 64.97931, 65.00147, 65.02328, 65.04474, 65.06583, 65.08658, 
    65.10697, 65.127, 65.14667, 65.16598, 65.18493, 65.20351, 65.22174, 
    65.2396, 65.2571, 65.27424, 65.29101, 65.30741, 65.32344, 65.33911, 
    65.35441, 65.36934, 65.3839, 65.39809, 65.4119, 65.42535, 65.43842, 
    65.45113, 65.46346, 65.4754, 65.48698, 65.49818, 65.50902, 65.51946, 
    65.52954, 65.53924, 65.54855, 65.5575, 65.56606, 65.57424, 65.58205, 
    65.58947, 65.59651, 65.60317, 65.60946, 65.61536, 65.62088, 65.62601, 
    65.63078, 65.63515, 65.63914, 65.64275, 65.64597, 65.64882, 65.65128, 
    65.65336, 65.65505, 65.65636, 65.6573, 65.65784, 65.658, 65.65778, 
    65.65717, 65.65618, 65.65481, 65.65305, 65.65092, 65.64839, 65.64549, 
    65.6422, 65.63853, 65.63448, 65.63004, 65.62523, 65.62003, 65.61445, 
    65.60849, 65.60214, 65.59542, 65.58832, 65.58083, 65.57297, 65.56473, 
    65.55611, 65.5471, 65.53773, 65.52797, 65.51784, 65.50732, 65.49644, 
    65.48518, 65.47354, 65.46152, 65.44914, 65.43639, 65.42325, 65.40974, 
    65.39587, 65.38162, 65.367, 65.35201, 65.33665, 65.32093, 65.30484, 
    65.28838, 65.27155, 65.25436, 65.2368, 65.21888, 65.2006, 65.18195, 
    65.16295, 65.14358, 65.12386, 65.10377, 65.08332, 65.06252, 65.04137, 
    65.01985, 64.99799, 64.97577, 64.95319, 64.93027, 64.907, 64.88338, 
    64.85941, 64.83508, 64.81042, 64.78541, 64.76006, 64.73435, 64.70831, 
    64.68193, 64.65521, 64.62815, 64.60075, 64.57301, 64.54494, 64.51654, 
    64.4878, 64.45873, 64.42933, 64.3996, 64.36954, 64.33915, 64.30844, 
    64.2774, 64.24603, 64.21435, 64.18234, 64.15002, 64.11737, 64.0844, 
    64.05112, 64.01753, 63.98362, 63.9494, 63.91486, 63.88002, 63.84486, 
    63.8094, 63.77364, 63.73756, 63.70119, 63.66451, 63.62753, 63.59024, 
    63.55267, 63.51479, 63.47662, 63.43815, 63.39939, 63.36033, 63.32099, 
    63.28135, 63.24143, 63.20122, 63.16073, 63.11995, 63.07889, 63.03754, 
    62.99592, 62.95402, 62.91183, 62.86938, 62.82665, 62.78364, 62.74036, 
    62.69682, 62.653, 62.60891, 62.56456, 62.51994, 62.47506, 62.42991, 
    62.3845, 62.33883, 62.2929, 62.24672, 62.20028, 62.15358, 62.10663, 
    62.05943, 62.01197, 61.96427, 61.91632, 61.86812, 61.81967, 61.77098, 
    61.72205, 61.67287, 61.62346, 61.5738, 61.52391, 61.47378, 61.42342, 
    61.37281, 61.32198, 61.27092, 61.21962, 61.1681, 61.11635, 61.06437, 
    61.01217, 60.95974, 60.90709, 60.85422, 60.80113, 60.74782, 60.69429, 
    60.64054, 60.58659,
  54.87667, 54.94601, 55.01522, 55.08432, 55.15329, 55.22213, 55.29085, 
    55.35945, 55.42792, 55.49626, 55.56448, 55.63256, 55.70052, 55.76835, 
    55.83604, 55.90361, 55.97104, 56.03834, 56.1055, 56.17253, 56.23942, 
    56.30618, 56.3728, 56.43927, 56.50561, 56.57181, 56.63787, 56.70378, 
    56.76955, 56.83518, 56.90066, 56.966, 57.03119, 57.09623, 57.16112, 
    57.22586, 57.29045, 57.35489, 57.41918, 57.48331, 57.54729, 57.61111, 
    57.67478, 57.73829, 57.80164, 57.86483, 57.92787, 57.99074, 58.05344, 
    58.11599, 58.17837, 58.24058, 58.30263, 58.36451, 58.42622, 58.48776, 
    58.54913, 58.61033, 58.67136, 58.73221, 58.79289, 58.85339, 58.91372, 
    58.97386, 59.03383, 59.09362, 59.15322, 59.21264, 59.27188, 59.33094, 
    59.3898, 59.44849, 59.50698, 59.56528, 59.6234, 59.68132, 59.73905, 
    59.79659, 59.85392, 59.91107, 59.96801, 60.02476, 60.08131, 60.13766, 
    60.1938, 60.24974, 60.30548, 60.36101, 60.41634, 60.47145, 60.52636, 
    60.58106, 60.63554, 60.68982, 60.74387, 60.79771, 60.85134, 60.90475, 
    60.95794, 61.0109, 61.06365, 61.11617, 61.16847, 61.22054, 61.27239, 
    61.32401, 61.3754, 61.42656, 61.47749, 61.52818, 61.57864, 61.62886, 
    61.67885, 61.7286, 61.7781, 61.82737, 61.8764, 61.92518, 61.97371, 
    62.022, 62.07005, 62.11784, 62.16539, 62.21268, 62.25972, 62.3065, 
    62.35303, 62.39931, 62.44532, 62.49108, 62.53657, 62.58181, 62.62677, 
    62.67148, 62.71592, 62.76009, 62.80399, 62.84762, 62.89098, 62.93407, 
    62.97688, 63.01942, 63.06168, 63.10366, 63.14537, 63.18679, 63.22793, 
    63.26878, 63.30936, 63.34964, 63.38964, 63.42935, 63.46877, 63.50789, 
    63.54673, 63.58527, 63.62351, 63.66146, 63.69911, 63.73646, 63.77351, 
    63.81025, 63.8467, 63.88284, 63.91867, 63.95419, 63.98941, 64.02431, 
    64.05891, 64.0932, 64.12717, 64.16082, 64.19416, 64.22718, 64.25989, 
    64.29227, 64.32433, 64.35606, 64.38748, 64.41857, 64.44933, 64.47977, 
    64.50988, 64.53966, 64.56911, 64.59822, 64.62701, 64.65546, 64.68357, 
    64.71134, 64.73878, 64.76588, 64.79264, 64.81906, 64.84514, 64.87086, 
    64.89626, 64.9213, 64.946, 64.97034, 64.99435, 65.018, 65.0413, 65.06425, 
    65.08684, 65.10909, 65.13097, 65.1525, 65.17368, 65.1945, 65.21496, 
    65.23505, 65.2548, 65.27418, 65.29319, 65.31185, 65.33014, 65.34807, 
    65.36563, 65.38282, 65.39965, 65.41611, 65.43221, 65.44793, 65.46329, 
    65.47827, 65.49288, 65.50713, 65.521, 65.53449, 65.54761, 65.56036, 
    65.57273, 65.58472, 65.59635, 65.60759, 65.61846, 65.62895, 65.63906, 
    65.6488, 65.65815, 65.66712, 65.67571, 65.68393, 65.69176, 65.69921, 
    65.70628, 65.71297, 65.71928, 65.7252, 65.73074, 65.73589, 65.74067, 
    65.74506, 65.74907, 65.75269, 65.75593, 65.75878, 65.76125, 65.76334, 
    65.76505, 65.76636, 65.76729, 65.76784, 65.768, 65.76778, 65.76717, 
    65.76617, 65.7648, 65.76304, 65.76089, 65.75836, 65.75544, 65.75214, 
    65.74846, 65.74439, 65.73994, 65.73511, 65.72989, 65.72429, 65.7183, 
    65.71194, 65.70518, 65.69806, 65.69054, 65.68266, 65.67438, 65.66573, 
    65.65669, 65.64728, 65.63749, 65.62731, 65.61677, 65.60584, 65.59454, 
    65.58286, 65.5708, 65.55836, 65.54556, 65.53238, 65.51882, 65.5049, 
    65.4906, 65.47592, 65.46088, 65.44547, 65.42969, 65.41354, 65.39702, 
    65.38013, 65.36288, 65.34525, 65.32727, 65.30892, 65.29021, 65.27113, 
    65.25169, 65.2319, 65.21174, 65.19122, 65.17035, 65.14912, 65.12753, 
    65.10559, 65.08329, 65.06064, 65.03764, 65.01427, 64.99057, 64.96651, 
    64.94212, 64.91736, 64.89227, 64.86682, 64.84103, 64.8149, 64.78843, 
    64.76162, 64.73447, 64.70697, 64.67915, 64.65098, 64.62247, 64.59364, 
    64.56448, 64.53497, 64.50514, 64.47498, 64.44449, 64.41367, 64.38254, 
    64.35107, 64.31927, 64.28716, 64.25473, 64.22198, 64.18891, 64.15552, 
    64.12182, 64.0878, 64.05346, 64.01881, 63.98386, 63.9486, 63.91302, 
    63.87714, 63.84095, 63.80446, 63.76767, 63.73057, 63.69317, 63.65548, 
    63.61748, 63.57919, 63.5406, 63.50172, 63.46255, 63.42308, 63.38333, 
    63.34329, 63.30296, 63.26234, 63.22144, 63.18026, 63.13879, 63.09704, 
    63.05502, 63.01271, 62.97013, 62.92727, 62.88414, 62.84074, 62.79706, 
    62.75312, 62.7089, 62.66442, 62.61968, 62.57467, 62.52939, 62.48386, 
    62.43806, 62.392, 62.34569, 62.29912, 62.25229, 62.20522, 62.15788, 
    62.1103, 62.06247, 62.01438, 61.96605, 61.91748, 61.86866, 61.8196, 
    61.77029, 61.72074, 61.67096, 61.62093, 61.57067, 61.52018, 61.46944, 
    61.41848, 61.36729, 61.31586, 61.26421, 61.21232, 61.16021, 61.10788, 
    61.05532, 61.00254, 60.94954, 60.89631, 60.84287, 60.78921, 60.73534, 
    60.68124,
  54.9599, 55.02935, 55.09867, 55.16787, 55.23695, 55.3059, 55.37473, 
    55.44344, 55.51202, 55.58047, 55.6488, 55.717, 55.78507, 55.85301, 
    55.92082, 55.98849, 56.05604, 56.12345, 56.19073, 56.25787, 56.32488, 
    56.39175, 56.45848, 56.52507, 56.59153, 56.65784, 56.72402, 56.79005, 
    56.85593, 56.92168, 56.98728, 57.05273, 57.11804, 57.1832, 57.24821, 
    57.31308, 57.37778, 57.44234, 57.50676, 57.57101, 57.63511, 57.69905, 
    57.76284, 57.82648, 57.88995, 57.95326, 58.01642, 58.07941, 58.14224, 
    58.20491, 58.26741, 58.32975, 58.39193, 58.45393, 58.51577, 58.57743, 
    58.63893, 58.70026, 58.76141, 58.82239, 58.88319, 58.94382, 59.00427, 
    59.06454, 59.12464, 59.18456, 59.24429, 59.30384, 59.3632, 59.42239, 
    59.48138, 59.5402, 59.59882, 59.65725, 59.71549, 59.77354, 59.83141, 
    59.88907, 59.94654, 60.00381, 60.06089, 60.11777, 60.17445, 60.23093, 
    60.2872, 60.34327, 60.39914, 60.4548, 60.51026, 60.56551, 60.62055, 
    60.67538, 60.72999, 60.7844, 60.83858, 60.89256, 60.94632, 60.99986, 
    61.05318, 61.10628, 61.15915, 61.21181, 61.26424, 61.31644, 61.36842, 
    61.42017, 61.47169, 61.52299, 61.57404, 61.62487, 61.67546, 61.72581, 
    61.77593, 61.82581, 61.87545, 61.92485, 61.97401, 62.02292, 62.07159, 
    62.12001, 62.16818, 62.21611, 62.26378, 62.3112, 62.35838, 62.40529, 
    62.45195, 62.49835, 62.54449, 62.59038, 62.636, 62.68137, 62.72646, 
    62.77129, 62.81586, 62.86016, 62.90419, 62.94794, 62.99143, 63.03465, 
    63.07758, 63.12025, 63.16263, 63.20474, 63.24657, 63.28811, 63.32938, 
    63.37036, 63.41105, 63.45146, 63.49158, 63.53141, 63.57095, 63.61019, 
    63.64915, 63.68781, 63.72617, 63.76424, 63.802, 63.83947, 63.87663, 
    63.9135, 63.95005, 63.98631, 64.02225, 64.05789, 64.09322, 64.12824, 
    64.16295, 64.19735, 64.23142, 64.26519, 64.29864, 64.33176, 64.36458, 
    64.39706, 64.42923, 64.46107, 64.4926, 64.52379, 64.55466, 64.5852, 
    64.6154, 64.64529, 64.67483, 64.70405, 64.73293, 64.76147, 64.78968, 
    64.81755, 64.84509, 64.87228, 64.89912, 64.92564, 64.95181, 64.97762, 
    65.0031, 65.02823, 65.05302, 65.07745, 65.10153, 65.12527, 65.14865, 
    65.17168, 65.19435, 65.21667, 65.23864, 65.26025, 65.2815, 65.30239, 
    65.32292, 65.34309, 65.36291, 65.38235, 65.40144, 65.42017, 65.43852, 
    65.45651, 65.47414, 65.4914, 65.50829, 65.52481, 65.54096, 65.55675, 
    65.57215, 65.5872, 65.60186, 65.61616, 65.63007, 65.64362, 65.65679, 
    65.66959, 65.682, 65.69405, 65.7057, 65.717, 65.7279, 65.73843, 65.74858, 
    65.75835, 65.76774, 65.77674, 65.78537, 65.79361, 65.80148, 65.80895, 
    65.81605, 65.82276, 65.82909, 65.83504, 65.8406, 65.84578, 65.85057, 
    65.85497, 65.85899, 65.86263, 65.86588, 65.86875, 65.87123, 65.87332, 
    65.87503, 65.87635, 65.87729, 65.87784, 65.878, 65.87778, 65.87717, 
    65.87617, 65.87479, 65.87302, 65.87086, 65.86832, 65.86539, 65.86208, 
    65.85838, 65.8543, 65.84984, 65.84499, 65.83974, 65.83412, 65.82812, 
    65.82172, 65.81495, 65.80779, 65.80025, 65.79234, 65.78403, 65.77534, 
    65.76627, 65.75683, 65.74699, 65.73679, 65.7262, 65.71523, 65.70389, 
    65.69216, 65.68006, 65.66759, 65.65473, 65.6415, 65.6279, 65.61391, 
    65.59956, 65.58484, 65.56974, 65.55428, 65.53843, 65.52222, 65.50564, 
    65.48869, 65.47137, 65.45369, 65.43565, 65.41723, 65.39845, 65.3793, 
    65.35979, 65.33993, 65.3197, 65.29911, 65.27816, 65.25685, 65.23519, 
    65.21317, 65.19079, 65.16806, 65.14497, 65.12154, 65.09775, 65.07361, 
    65.04912, 65.02428, 64.99909, 64.97356, 64.94769, 64.92146, 64.89491, 
    64.868, 64.84075, 64.81316, 64.78524, 64.75698, 64.72838, 64.69945, 
    64.67018, 64.64058, 64.61065, 64.58038, 64.5498, 64.51888, 64.48763, 
    64.45606, 64.42416, 64.39194, 64.35941, 64.32655, 64.29337, 64.25987, 
    64.22606, 64.19193, 64.15749, 64.12273, 64.08765, 64.05228, 64.01659, 
    63.98059, 63.94429, 63.90768, 63.87077, 63.83356, 63.79605, 63.75823, 
    63.72012, 63.68171, 63.64301, 63.604, 63.56471, 63.52513, 63.48525, 
    63.44508, 63.40463, 63.36389, 63.32287, 63.28156, 63.23997, 63.1981, 
    63.15595, 63.11352, 63.07081, 63.02783, 62.98457, 62.94104, 62.89724, 
    62.85317, 62.80883, 62.76422, 62.71935, 62.67421, 62.6288, 62.58314, 
    62.53721, 62.49103, 62.44458, 62.39788, 62.35093, 62.30372, 62.25626, 
    62.20854, 62.16058, 62.11237, 62.06391, 62.0152, 61.96625, 61.91705, 
    61.86762, 61.81794, 61.76802, 61.71786, 61.66747, 61.61684, 61.56598, 
    61.51489, 61.46356, 61.412, 61.36022, 61.3082, 61.25596, 61.2035, 
    61.1508, 61.09789, 61.04476, 60.9914, 60.93783, 60.88404, 60.83003, 
    60.7758,
  55.043, 55.11255, 55.18198, 55.25129, 55.32048, 55.38955, 55.45848, 
    55.5273, 55.59599, 55.66456, 55.733, 55.80131, 55.86949, 55.93754, 
    56.00546, 56.07325, 56.14091, 56.20844, 56.27583, 56.34308, 56.41021, 
    56.47719, 56.54404, 56.61075, 56.67732, 56.74375, 56.81004, 56.87619, 
    56.9422, 57.00806, 57.07378, 57.13935, 57.20478, 57.27005, 57.33519, 
    57.40017, 57.465, 57.52968, 57.59421, 57.65858, 57.72281, 57.78687, 
    57.85078, 57.91454, 57.97813, 58.04157, 58.10485, 58.16797, 58.23092, 
    58.29372, 58.35634, 58.4188, 58.4811, 58.54323, 58.60519, 58.66699, 
    58.72861, 58.79006, 58.85134, 58.91245, 58.97338, 59.03413, 59.09472, 
    59.15511, 59.21534, 59.27538, 59.33524, 59.39492, 59.45442, 59.51373, 
    59.57286, 59.63179, 59.69055, 59.74911, 59.80748, 59.86566, 59.92365, 
    59.98145, 60.03905, 60.09645, 60.15366, 60.21067, 60.26748, 60.32409, 
    60.3805, 60.4367, 60.4927, 60.5485, 60.60408, 60.65946, 60.71463, 
    60.7696, 60.82434, 60.87888, 60.9332, 60.98731, 61.04119, 61.09487, 
    61.14832, 61.20155, 61.25456, 61.30735, 61.35992, 61.41225, 61.46436, 
    61.51625, 61.5679, 61.61932, 61.67051, 61.72147, 61.77219, 61.82268, 
    61.87293, 61.92294, 61.97272, 62.02225, 62.07154, 62.12058, 62.16938, 
    62.21793, 62.26624, 62.31429, 62.3621, 62.40965, 62.45695, 62.504, 
    62.55079, 62.59732, 62.64359, 62.68961, 62.73536, 62.78085, 62.82608, 
    62.87104, 62.91573, 62.96016, 63.00431, 63.0482, 63.09181, 63.13515, 
    63.17822, 63.22101, 63.26352, 63.30575, 63.34771, 63.38937, 63.43076, 
    63.47187, 63.51268, 63.55321, 63.59346, 63.63341, 63.67307, 63.71244, 
    63.75151, 63.79029, 63.82877, 63.86695, 63.90484, 63.94242, 63.97971, 
    64.01669, 64.05336, 64.08973, 64.12579, 64.16154, 64.19699, 64.23212, 
    64.26694, 64.30145, 64.33564, 64.36951, 64.40307, 64.43631, 64.46923, 
    64.50182, 64.5341, 64.56605, 64.59767, 64.62897, 64.65994, 64.69058, 
    64.72089, 64.75087, 64.78052, 64.80983, 64.83881, 64.86745, 64.89576, 
    64.92373, 64.95135, 64.97864, 65.00558, 65.03219, 65.05844, 65.08435, 
    65.10992, 65.13514, 65.16, 65.18452, 65.20869, 65.23251, 65.25598, 
    65.27909, 65.30184, 65.32424, 65.34629, 65.36797, 65.38931, 65.41027, 
    65.43088, 65.45112, 65.471, 65.49052, 65.50968, 65.52847, 65.54689, 
    65.56495, 65.58264, 65.59996, 65.61691, 65.63349, 65.6497, 65.66554, 
    65.68102, 65.69611, 65.71083, 65.72517, 65.73914, 65.75274, 65.76596, 
    65.7788, 65.79127, 65.80335, 65.81506, 65.82639, 65.83733, 65.8479, 
    65.85809, 65.8679, 65.87732, 65.88636, 65.89502, 65.9033, 65.91119, 
    65.91869, 65.92582, 65.93256, 65.9389, 65.94488, 65.95045, 65.95565, 
    65.96046, 65.96489, 65.96893, 65.97257, 65.97584, 65.97871, 65.9812, 
    65.98331, 65.98502, 65.98634, 65.98728, 65.98784, 65.988, 65.98778, 
    65.98716, 65.98616, 65.98477, 65.983, 65.98083, 65.97829, 65.97535, 
    65.97202, 65.96832, 65.96421, 65.95973, 65.95486, 65.9496, 65.94395, 
    65.93793, 65.93151, 65.92471, 65.91753, 65.90997, 65.90201, 65.89368, 
    65.88496, 65.87585, 65.86637, 65.85651, 65.84626, 65.83563, 65.82462, 
    65.81323, 65.80147, 65.78932, 65.77679, 65.76389, 65.75062, 65.73696, 
    65.72293, 65.70853, 65.69375, 65.67859, 65.66306, 65.64716, 65.6309, 
    65.61426, 65.59724, 65.57986, 65.56212, 65.54401, 65.52552, 65.50668, 
    65.48746, 65.46788, 65.44794, 65.42764, 65.40697, 65.38595, 65.36457, 
    65.34283, 65.32072, 65.29827, 65.27546, 65.25229, 65.22877, 65.2049, 
    65.18067, 65.1561, 65.13117, 65.1059, 65.08028, 65.05431, 65.028, 
    65.00134, 64.97434, 64.94701, 64.91933, 64.8913, 64.86295, 64.83425, 
    64.80522, 64.77585, 64.74615, 64.71612, 64.68575, 64.65506, 64.62404, 
    64.59269, 64.56101, 64.52901, 64.49669, 64.46404, 64.43108, 64.39778, 
    64.36417, 64.33025, 64.29601, 64.26146, 64.22659, 64.19141, 64.15591, 
    64.12011, 64.084, 64.04758, 64.01086, 63.97383, 63.9365, 63.89887, 
    63.86094, 63.8227, 63.78418, 63.74535, 63.70623, 63.66681, 63.62711, 
    63.58711, 63.54682, 63.50624, 63.46538, 63.42424, 63.3828, 63.34109, 
    63.29909, 63.25681, 63.21426, 63.17142, 63.12831, 63.08493, 63.04128, 
    62.99735, 62.95315, 62.90868, 62.86394, 62.81894, 62.77367, 62.72814, 
    62.68235, 62.63629, 62.58998, 62.5434, 62.49657, 62.44949, 62.40215, 
    62.35455, 62.30671, 62.25861, 62.21027, 62.16167, 62.11284, 62.06376, 
    62.01443, 61.96486, 61.91505, 61.865, 61.81471, 61.76419, 61.71343, 
    61.66243, 61.61121, 61.55975, 61.50806, 61.45613, 61.40399, 61.35162, 
    61.29902, 61.24619, 61.19315, 61.13988, 61.08639, 61.03269, 60.97876, 
    60.92462, 60.87027,
  55.12597, 55.19563, 55.26517, 55.33459, 55.40388, 55.47306, 55.54211, 
    55.61103, 55.67984, 55.74851, 55.81706, 55.88549, 55.95378, 56.02194, 
    56.08998, 56.15788, 56.22565, 56.29329, 56.3608, 56.42817, 56.49541, 
    56.56251, 56.62947, 56.6963, 56.76299, 56.82953, 56.89594, 56.96221, 
    57.02833, 57.09431, 57.16015, 57.22584, 57.29139, 57.35678, 57.42204, 
    57.48714, 57.55209, 57.61689, 57.68154, 57.74604, 57.81038, 57.87457, 
    57.93861, 58.00248, 58.0662, 58.12976, 58.19316, 58.2564, 58.31948, 
    58.3824, 58.44515, 58.50774, 58.57016, 58.63242, 58.69451, 58.75642, 
    58.81818, 58.87975, 58.94116, 59.00239, 59.06345, 59.12433, 59.18504, 
    59.24557, 59.30592, 59.36609, 59.42608, 59.48589, 59.54552, 59.60496, 
    59.66421, 59.72328, 59.78217, 59.84086, 59.89936, 59.95767, 60.01579, 
    60.07372, 60.13145, 60.18899, 60.24633, 60.30347, 60.36041, 60.41715, 
    60.47369, 60.53003, 60.58615, 60.64208, 60.6978, 60.75331, 60.80862, 
    60.86371, 60.91859, 60.97326, 61.02772, 61.08195, 61.13598, 61.18979, 
    61.24337, 61.29673, 61.34988, 61.4028, 61.45549, 61.50797, 61.56021, 
    61.61223, 61.66401, 61.71557, 61.7669, 61.81799, 61.86884, 61.91946, 
    61.96984, 62.01999, 62.06989, 62.11956, 62.16898, 62.21815, 62.26709, 
    62.31577, 62.36421, 62.4124, 62.46033, 62.50801, 62.55545, 62.60262, 
    62.64954, 62.69621, 62.74261, 62.78876, 62.83464, 62.88026, 62.92562, 
    62.97071, 63.01553, 63.06009, 63.10437, 63.14838, 63.19213, 63.23559, 
    63.27879, 63.3217, 63.36434, 63.4067, 63.44878, 63.49057, 63.53209, 
    63.57331, 63.61425, 63.65491, 63.69527, 63.73535, 63.77513, 63.81462, 
    63.85381, 63.89272, 63.93132, 63.96962, 64.00763, 64.04533, 64.08273, 
    64.11983, 64.15662, 64.19311, 64.22928, 64.26515, 64.3007, 64.33595, 
    64.37089, 64.4055, 64.43981, 64.47379, 64.50746, 64.54081, 64.57384, 
    64.60654, 64.63892, 64.67097, 64.70271, 64.73411, 64.76518, 64.79593, 
    64.82635, 64.85642, 64.88618, 64.91559, 64.94466, 64.9734, 65.00181, 
    65.02987, 65.05759, 65.08498, 65.11201, 65.1387, 65.16505, 65.19106, 
    65.21671, 65.24202, 65.26698, 65.29158, 65.31583, 65.33974, 65.36329, 
    65.38648, 65.40932, 65.43179, 65.45392, 65.47569, 65.49709, 65.51813, 
    65.53881, 65.55913, 65.57909, 65.59867, 65.6179, 65.63676, 65.65525, 
    65.67337, 65.69112, 65.70851, 65.72552, 65.74217, 65.75844, 65.77434, 
    65.78986, 65.80502, 65.81979, 65.83419, 65.84821, 65.86185, 65.87512, 
    65.88802, 65.90053, 65.91266, 65.92441, 65.93578, 65.94677, 65.95737, 
    65.9676, 65.97744, 65.9869, 65.99598, 66.00467, 66.01297, 66.0209, 
    66.02843, 66.03558, 66.04234, 66.04872, 66.05471, 66.06032, 66.06553, 
    66.07036, 66.0748, 66.07885, 66.08252, 66.08579, 66.08868, 66.09118, 
    66.09328, 66.09501, 66.09634, 66.09728, 66.09783, 66.098, 66.09777, 
    66.09716, 66.09615, 66.09476, 66.09298, 66.09081, 66.08825, 66.0853, 
    66.08196, 66.07824, 66.07413, 66.06962, 66.06474, 66.05946, 66.05379, 
    66.04774, 66.0413, 66.03448, 66.02726, 66.01967, 66.01169, 66.00332, 
    65.99457, 65.98543, 65.97591, 65.96601, 65.95572, 65.94505, 65.93401, 
    65.92258, 65.91077, 65.89857, 65.886, 65.87305, 65.85973, 65.84602, 
    65.83193, 65.81747, 65.80264, 65.78743, 65.77185, 65.75589, 65.73956, 
    65.72286, 65.70579, 65.68834, 65.67053, 65.65235, 65.6338, 65.61488, 
    65.5956, 65.57595, 65.55594, 65.53556, 65.51482, 65.49373, 65.47227, 
    65.45045, 65.42827, 65.40573, 65.38284, 65.35959, 65.33598, 65.31202, 
    65.28771, 65.26305, 65.23804, 65.21268, 65.18697, 65.16091, 65.13451, 
    65.10776, 65.08067, 65.05323, 65.02545, 64.99734, 64.96888, 64.94009, 
    64.91096, 64.88149, 64.85169, 64.82156, 64.79109, 64.76029, 64.72916, 
    64.69771, 64.66593, 64.63382, 64.60139, 64.56863, 64.53555, 64.50216, 
    64.46844, 64.4344, 64.40005, 64.36538, 64.3304, 64.2951, 64.2595, 
    64.22358, 64.18736, 64.15082, 64.11398, 64.07684, 64.03938, 64.00163, 
    63.96358, 63.92523, 63.88658, 63.84763, 63.80839, 63.76886, 63.72903, 
    63.68891, 63.64849, 63.6078, 63.56681, 63.52554, 63.48398, 63.44214, 
    63.40002, 63.35761, 63.31493, 63.27197, 63.22874, 63.18522, 63.14144, 
    63.09738, 63.05305, 63.00846, 62.96359, 62.91846, 62.87306, 62.8274, 
    62.78148, 62.73529, 62.68884, 62.64214, 62.59518, 62.54796, 62.50049, 
    62.45277, 62.40479, 62.35656, 62.30809, 62.25936, 62.21039, 62.16117, 
    62.11172, 62.06202, 62.01207, 61.96189, 61.91147, 61.86081, 61.80992, 
    61.75879, 61.70743, 61.65584, 61.60402, 61.55196, 61.49968, 61.44717, 
    61.39444, 61.34149, 61.28831, 61.23491, 61.18129, 61.12745, 61.07339, 
    61.01912, 60.96463,
  55.20881, 55.27857, 55.34822, 55.41775, 55.48716, 55.55644, 55.6256, 
    55.69464, 55.76355, 55.83234, 55.901, 55.96954, 56.03794, 56.10622, 
    56.17437, 56.24238, 56.31027, 56.37802, 56.44564, 56.51313, 56.58048, 
    56.6477, 56.71478, 56.78172, 56.84853, 56.91519, 56.98171, 57.0481, 
    57.11434, 57.18044, 57.2464, 57.31221, 57.37787, 57.44339, 57.50876, 
    57.57398, 57.63905, 57.70398, 57.76875, 57.83337, 57.89783, 57.96215, 
    58.0263, 58.0903, 58.15414, 58.21783, 58.28135, 58.34472, 58.40792, 
    58.47096, 58.53384, 58.59655, 58.6591, 58.72149, 58.7837, 58.84575, 
    58.90762, 58.96933, 59.03086, 59.09222, 59.1534, 59.21442, 59.27525, 
    59.33591, 59.39639, 59.45669, 59.51681, 59.57675, 59.6365, 59.69607, 
    59.75546, 59.81466, 59.87367, 59.9325, 59.99113, 60.04957, 60.10782, 
    60.16588, 60.22374, 60.28141, 60.33888, 60.39616, 60.45323, 60.5101, 
    60.56677, 60.62324, 60.67951, 60.73557, 60.79142, 60.84706, 60.9025, 
    60.95773, 61.01274, 61.06754, 61.12213, 61.17651, 61.23066, 61.2846, 
    61.33832, 61.39182, 61.4451, 61.49815, 61.55098, 61.60358, 61.65596, 
    61.70811, 61.76004, 61.81173, 61.86318, 61.91441, 61.9654, 62.01615, 
    62.06667, 62.11694, 62.16698, 62.21678, 62.26633, 62.31564, 62.36471, 
    62.41352, 62.46209, 62.51041, 62.55848, 62.6063, 62.65386, 62.70117, 
    62.74823, 62.79502, 62.84156, 62.88783, 62.93385, 62.9796, 63.02508, 
    63.0703, 63.11525, 63.15994, 63.20435, 63.2485, 63.29237, 63.33596, 
    63.37928, 63.42233, 63.46509, 63.50758, 63.54978, 63.5917, 63.63334, 
    63.67469, 63.71576, 63.75654, 63.79703, 63.83723, 63.87713, 63.91674, 
    63.95606, 63.99508, 64.03381, 64.07224, 64.11036, 64.14818, 64.1857, 
    64.22292, 64.25983, 64.29642, 64.33272, 64.36871, 64.40437, 64.43974, 
    64.47478, 64.50951, 64.54393, 64.57803, 64.61181, 64.64526, 64.6784, 
    64.71121, 64.74371, 64.77586, 64.8077, 64.83921, 64.87039, 64.90124, 
    64.93176, 64.96194, 64.99179, 65.02131, 65.05048, 65.07932, 65.10783, 
    65.13599, 65.1638, 65.19128, 65.21841, 65.2452, 65.27164, 65.29773, 
    65.32348, 65.34888, 65.37392, 65.39861, 65.42295, 65.44694, 65.47057, 
    65.49385, 65.51677, 65.53933, 65.56153, 65.58337, 65.60485, 65.62597, 
    65.64673, 65.66712, 65.68715, 65.70681, 65.7261, 65.74503, 65.76359, 
    65.78178, 65.7996, 65.81705, 65.83413, 65.85083, 65.86716, 65.88312, 
    65.8987, 65.91391, 65.92874, 65.94319, 65.95727, 65.97096, 65.98428, 
    65.99722, 66.00978, 66.02196, 66.03375, 66.04517, 66.05619, 66.06684, 
    66.0771, 66.08698, 66.09648, 66.10559, 66.11431, 66.12265, 66.1306, 
    66.13817, 66.14534, 66.15213, 66.15853, 66.16454, 66.17017, 66.17541, 
    66.18025, 66.18472, 66.18878, 66.19246, 66.19575, 66.19865, 66.20115, 
    66.20327, 66.20499, 66.20634, 66.20728, 66.20783, 66.208, 66.20777, 
    66.20715, 66.20615, 66.20475, 66.20296, 66.20078, 66.19821, 66.19525, 
    66.1919, 66.18816, 66.18404, 66.17951, 66.17461, 66.1693, 66.16362, 
    66.15755, 66.15108, 66.14423, 66.13699, 66.12937, 66.12135, 66.11296, 
    66.10417, 66.095, 66.08545, 66.07551, 66.06519, 66.05447, 66.04338, 
    66.03191, 66.02005, 66.00782, 65.9952, 65.9822, 65.96882, 65.95506, 
    65.94093, 65.92641, 65.91153, 65.89626, 65.88062, 65.8646, 65.84821, 
    65.83145, 65.81432, 65.79681, 65.77893, 65.76068, 65.74207, 65.72308, 
    65.70373, 65.68401, 65.66392, 65.64347, 65.62266, 65.60148, 65.57994, 
    65.55804, 65.53578, 65.51317, 65.49019, 65.46686, 65.44317, 65.41913, 
    65.39473, 65.36998, 65.34488, 65.31943, 65.29362, 65.26748, 65.24098, 
    65.21414, 65.18696, 65.15942, 65.13155, 65.10334, 65.07478, 65.04589, 
    65.01666, 64.98709, 64.95719, 64.92696, 64.89639, 64.86548, 64.83425, 
    64.80269, 64.7708, 64.73859, 64.70605, 64.67318, 64.63999, 64.60648, 
    64.57265, 64.53851, 64.50404, 64.46926, 64.43417, 64.39876, 64.36303, 
    64.327, 64.29066, 64.25401, 64.21705, 64.17979, 64.14222, 64.10435, 
    64.06617, 64.0277, 63.98893, 63.94986, 63.9105, 63.87084, 63.83089, 
    63.79064, 63.75011, 63.70928, 63.66817, 63.62677, 63.58509, 63.54313, 
    63.50087, 63.45834, 63.41553, 63.37245, 63.32909, 63.28545, 63.24153, 
    63.19735, 63.15289, 63.10816, 63.06317, 63.0179, 62.97238, 62.92658, 
    62.88053, 62.83421, 62.78764, 62.7408, 62.69371, 62.64636, 62.59875, 
    62.5509, 62.50279, 62.45443, 62.40582, 62.35696, 62.30786, 62.25851, 
    62.20892, 62.15908, 62.10901, 62.05869, 62.00814, 61.95735, 61.90632, 
    61.85506, 61.80356, 61.75184, 61.69988, 61.64769, 61.59528, 61.54264, 
    61.48977, 61.43668, 61.38337, 61.32984, 61.27608, 61.22211, 61.16792, 
    61.11351, 61.05889,
  55.29151, 55.36139, 55.43114, 55.50078, 55.5703, 55.63969, 55.70897, 
    55.77811, 55.84713, 55.91603, 55.98481, 56.05345, 56.12197, 56.19036, 
    56.25862, 56.32675, 56.39475, 56.46262, 56.53036, 56.59796, 56.66543, 
    56.73276, 56.79995, 56.86701, 56.93393, 57.00072, 57.06736, 57.13386, 
    57.20022, 57.26644, 57.33251, 57.39845, 57.46423, 57.52987, 57.59536, 
    57.6607, 57.72589, 57.79094, 57.85583, 57.92057, 57.98516, 58.04959, 
    58.11388, 58.178, 58.24197, 58.30577, 58.36942, 58.43291, 58.49624, 
    58.55941, 58.62241, 58.68525, 58.74792, 58.81043, 58.87277, 58.93494, 
    58.99695, 59.05878, 59.12044, 59.18193, 59.24324, 59.30438, 59.36535, 
    59.42613, 59.48674, 59.54717, 59.60742, 59.66749, 59.72738, 59.78708, 
    59.84659, 59.90592, 59.96507, 60.02402, 60.08279, 60.14136, 60.19974, 
    60.25793, 60.31593, 60.37373, 60.43133, 60.48874, 60.54594, 60.60295, 
    60.65975, 60.71635, 60.77275, 60.82895, 60.88493, 60.94071, 60.99628, 
    61.05164, 61.10679, 61.16172, 61.21645, 61.27095, 61.32524, 61.37932, 
    61.43317, 61.4868, 61.54022, 61.59341, 61.64637, 61.69911, 61.75162, 
    61.80391, 61.85596, 61.90779, 61.95938, 62.01074, 62.06186, 62.11275, 
    62.1634, 62.21381, 62.26398, 62.31391, 62.3636, 62.41304, 62.46224, 
    62.51119, 62.55989, 62.60835, 62.65655, 62.7045, 62.7522, 62.79964, 
    62.84682, 62.89375, 62.94042, 62.98683, 63.03297, 63.07885, 63.12447, 
    63.16982, 63.2149, 63.25972, 63.30426, 63.34854, 63.39254, 63.43626, 
    63.47971, 63.52288, 63.56578, 63.60839, 63.65072, 63.69277, 63.73453, 
    63.77601, 63.8172, 63.85811, 63.89872, 63.93904, 63.97907, 64.01881, 
    64.05825, 64.0974, 64.13624, 64.17478, 64.21303, 64.25098, 64.28861, 
    64.32594, 64.36298, 64.3997, 64.4361, 64.47221, 64.508, 64.54347, 
    64.57864, 64.61348, 64.64801, 64.68222, 64.71611, 64.74968, 64.78292, 
    64.81585, 64.84844, 64.88071, 64.91266, 64.94427, 64.97556, 65.00652, 
    65.03714, 65.06742, 65.09737, 65.12699, 65.15627, 65.18521, 65.21381, 
    65.24207, 65.26998, 65.29755, 65.32478, 65.35166, 65.3782, 65.40438, 
    65.43021, 65.4557, 65.48083, 65.50562, 65.53004, 65.55412, 65.57784, 
    65.6012, 65.6242, 65.64684, 65.66912, 65.69104, 65.7126, 65.7338, 
    65.75463, 65.77509, 65.7952, 65.81493, 65.8343, 65.85329, 65.87192, 
    65.89017, 65.90807, 65.92558, 65.94272, 65.95948, 65.97588, 65.99189, 
    66.00753, 66.0228, 66.03768, 66.05219, 66.06631, 66.08006, 66.09343, 
    66.10641, 66.11903, 66.13125, 66.14309, 66.15454, 66.16561, 66.1763, 
    66.18661, 66.19652, 66.20605, 66.21519, 66.22395, 66.23232, 66.2403, 
    66.24789, 66.2551, 66.26192, 66.26834, 66.27438, 66.28003, 66.28529, 
    66.29015, 66.29462, 66.29871, 66.3024, 66.3057, 66.30861, 66.31113, 
    66.31326, 66.31499, 66.31633, 66.31728, 66.31783, 66.318, 66.31777, 
    66.31715, 66.31614, 66.31474, 66.31294, 66.31075, 66.30817, 66.30521, 
    66.30184, 66.29809, 66.29394, 66.28941, 66.28448, 66.27916, 66.27345, 
    66.26735, 66.26086, 66.25399, 66.24672, 66.23907, 66.23103, 66.2226, 
    66.21378, 66.20457, 66.19498, 66.185, 66.17464, 66.16389, 66.15276, 
    66.14124, 66.12934, 66.11706, 66.10439, 66.09134, 66.07791, 66.0641, 
    66.04992, 66.03535, 66.02041, 66.00508, 65.98938, 65.9733, 65.95686, 
    65.94003, 65.92283, 65.90526, 65.88731, 65.869, 65.85031, 65.83125, 
    65.81183, 65.79204, 65.77188, 65.75136, 65.73047, 65.70921, 65.6876, 
    65.66562, 65.64328, 65.62058, 65.59753, 65.5741, 65.55033, 65.52621, 
    65.50172, 65.47688, 65.4517, 65.42616, 65.40026, 65.37402, 65.34743, 
    65.3205, 65.29321, 65.26559, 65.23762, 65.2093, 65.18066, 65.15166, 
    65.12233, 65.09266, 65.06265, 65.03232, 65.00164, 64.97063, 64.9393, 
    64.90763, 64.87563, 64.84331, 64.81066, 64.77769, 64.74438, 64.71077, 
    64.67683, 64.64256, 64.60799, 64.57309, 64.53788, 64.50236, 64.46651, 
    64.43037, 64.39391, 64.35714, 64.32006, 64.28268, 64.24499, 64.207, 
    64.16871, 64.13011, 64.09122, 64.05203, 64.01254, 63.97276, 63.93269, 
    63.89231, 63.85166, 63.81071, 63.76947, 63.72795, 63.68613, 63.64404, 
    63.60167, 63.55901, 63.51607, 63.47285, 63.42936, 63.38559, 63.34155, 
    63.29724, 63.25265, 63.20779, 63.16267, 63.11727, 63.07161, 63.02569, 
    62.9795, 62.93306, 62.88634, 62.83938, 62.79215, 62.74467, 62.69693, 
    62.64894, 62.6007, 62.55221, 62.50347, 62.45448, 62.40524, 62.35576, 
    62.30603, 62.25606, 62.20585, 62.1554, 62.10471, 62.05379, 62.00263, 
    61.95123, 61.8996, 61.84774, 61.79565, 61.74333, 61.69078, 61.63801, 
    61.58501, 61.53178, 61.47834, 61.42467, 61.37078, 61.31667, 61.26235, 
    61.20781, 61.15305,
  55.37408, 55.44407, 55.51394, 55.58368, 55.65331, 55.72281, 55.79219, 
    55.86145, 55.93059, 55.9996, 56.06848, 56.13724, 56.20587, 56.27438, 
    56.34275, 56.411, 56.47911, 56.54709, 56.61494, 56.68266, 56.75024, 
    56.81769, 56.885, 56.95218, 57.01921, 57.08612, 57.15288, 57.2195, 
    57.28598, 57.35231, 57.41851, 57.48455, 57.55046, 57.61622, 57.68183, 
    57.7473, 57.81261, 57.87778, 57.94279, 58.00765, 58.07236, 58.13692, 
    58.20132, 58.26557, 58.32966, 58.39359, 58.45737, 58.52098, 58.58443, 
    58.64773, 58.71086, 58.77382, 58.83662, 58.89926, 58.96172, 59.02402, 
    59.08615, 59.14811, 59.2099, 59.27152, 59.33296, 59.39423, 59.45533, 
    59.51624, 59.57698, 59.63754, 59.69792, 59.75811, 59.81813, 59.87796, 
    59.93761, 59.99707, 60.05635, 60.11543, 60.17433, 60.23304, 60.29155, 
    60.34987, 60.408, 60.46593, 60.52367, 60.58121, 60.63855, 60.69569, 
    60.75262, 60.80936, 60.86589, 60.92222, 60.97834, 61.03425, 61.08995, 
    61.14545, 61.20073, 61.2558, 61.31066, 61.3653, 61.41973, 61.47393, 
    61.52792, 61.58169, 61.63524, 61.68856, 61.74166, 61.79454, 61.84718, 
    61.8996, 61.95179, 62.00375, 62.05548, 62.10697, 62.15823, 62.20926, 
    62.26004, 62.31059, 62.36089, 62.41096, 62.46078, 62.51036, 62.55969, 
    62.60878, 62.65761, 62.7062, 62.75454, 62.80262, 62.85045, 62.89803, 
    62.94534, 62.9924, 63.0392, 63.08574, 63.13202, 63.17804, 63.22378, 
    63.26926, 63.31448, 63.35942, 63.4041, 63.44851, 63.49263, 63.53649, 
    63.58007, 63.62337, 63.66639, 63.70913, 63.75159, 63.79377, 63.83566, 
    63.87727, 63.91858, 63.95961, 64.00035, 64.0408, 64.08096, 64.12081, 
    64.16038, 64.19965, 64.23861, 64.27728, 64.31565, 64.35371, 64.39147, 
    64.42892, 64.46607, 64.50291, 64.53944, 64.57566, 64.61156, 64.64716, 
    64.68243, 64.71739, 64.75204, 64.78636, 64.82037, 64.85404, 64.88741, 
    64.92043, 64.95314, 64.98553, 65.01758, 65.0493, 65.08069, 65.11175, 
    65.14248, 65.17287, 65.20292, 65.23264, 65.26202, 65.29106, 65.31976, 
    65.34811, 65.37613, 65.40379, 65.43112, 65.45809, 65.48473, 65.511, 
    65.53693, 65.56251, 65.58773, 65.6126, 65.63712, 65.66127, 65.68507, 
    65.70852, 65.73161, 65.75433, 65.77669, 65.79869, 65.82033, 65.84161, 
    65.86251, 65.88305, 65.90323, 65.92303, 65.94247, 65.96154, 65.98023, 
    65.99856, 66.01651, 66.03409, 66.05129, 66.06812, 66.08457, 66.10065, 
    66.11635, 66.13167, 66.14661, 66.16117, 66.17535, 66.18916, 66.20258, 
    66.21561, 66.22826, 66.24053, 66.25242, 66.26392, 66.27503, 66.28576, 
    66.2961, 66.30605, 66.31562, 66.3248, 66.3336, 66.342, 66.35001, 
    66.35763, 66.36486, 66.3717, 66.37815, 66.38421, 66.38988, 66.39516, 
    66.40004, 66.40453, 66.40863, 66.41234, 66.41565, 66.41857, 66.4211, 
    66.42323, 66.42497, 66.42632, 66.42728, 66.42783, 66.428, 66.42777, 
    66.42715, 66.42613, 66.42472, 66.42292, 66.42072, 66.41814, 66.41515, 
    66.41178, 66.40801, 66.40385, 66.39929, 66.39435, 66.38901, 66.38328, 
    66.37716, 66.37064, 66.36374, 66.35645, 66.34876, 66.34069, 66.33223, 
    66.32337, 66.31413, 66.3045, 66.29449, 66.28409, 66.2733, 66.26212, 
    66.25056, 66.23862, 66.22629, 66.21357, 66.20048, 66.187, 66.17313, 
    66.1589, 66.14427, 66.12927, 66.11389, 66.09814, 66.082, 66.06548, 
    66.0486, 66.03133, 66.01369, 65.99568, 65.9773, 65.95855, 65.93942, 
    65.91992, 65.90006, 65.87983, 65.85923, 65.83826, 65.81693, 65.79523, 
    65.77318, 65.75076, 65.72797, 65.70483, 65.68134, 65.65748, 65.63326, 
    65.60869, 65.58376, 65.55849, 65.53285, 65.50687, 65.48054, 65.45385, 
    65.42682, 65.39944, 65.37172, 65.34365, 65.31524, 65.28649, 65.25739, 
    65.22796, 65.19819, 65.16808, 65.13764, 65.10686, 65.07574, 65.0443, 
    65.01253, 64.98042, 64.94799, 64.91523, 64.88215, 64.84874, 64.815, 
    64.78095, 64.74657, 64.71188, 64.67687, 64.64155, 64.6059, 64.56995, 
    64.53368, 64.49711, 64.46022, 64.42302, 64.38552, 64.34771, 64.3096, 
    64.27119, 64.23247, 64.19345, 64.15414, 64.11452, 64.07462, 64.03442, 
    63.99393, 63.95314, 63.91207, 63.8707, 63.82905, 63.78711, 63.74489, 
    63.70239, 63.6596, 63.61654, 63.57319, 63.52957, 63.48567, 63.4415, 
    63.39705, 63.35233, 63.30735, 63.26209, 63.21656, 63.17077, 63.12472, 
    63.0784, 63.03182, 62.98497, 62.93787, 62.89051, 62.8429, 62.79503, 
    62.74691, 62.69853, 62.64991, 62.60103, 62.5519, 62.50253, 62.45292, 
    62.40306, 62.35295, 62.30261, 62.25202, 62.2012, 62.15014, 62.09884, 
    62.04731, 61.99555, 61.94355, 61.89133, 61.83887, 61.78619, 61.73328, 
    61.68014, 61.62678, 61.5732, 61.5194, 61.46537, 61.41113, 61.35667, 
    61.302, 61.24711,
  55.45652, 55.52662, 55.59659, 55.66645, 55.73618, 55.8058, 55.87529, 
    55.94466, 56.0139, 56.08303, 56.15202, 56.22089, 56.28964, 56.35826, 
    56.42674, 56.4951, 56.56333, 56.63143, 56.69939, 56.76723, 56.83493, 
    56.90249, 56.96992, 57.03721, 57.10437, 57.17138, 57.23826, 57.305, 
    57.3716, 57.43805, 57.50437, 57.57054, 57.63656, 57.70244, 57.76817, 
    57.83376, 57.8992, 57.96449, 58.02962, 58.09461, 58.15944, 58.22412, 
    58.28865, 58.35302, 58.41723, 58.48129, 58.54519, 58.60893, 58.67251, 
    58.73592, 58.79918, 58.86227, 58.9252, 58.98796, 59.05056, 59.11298, 
    59.17524, 59.23733, 59.29924, 59.36099, 59.42256, 59.48396, 59.54518, 
    59.60623, 59.6671, 59.72779, 59.7883, 59.84863, 59.90877, 59.96873, 
    60.02851, 60.0881, 60.14751, 60.20673, 60.26576, 60.3246, 60.38325, 
    60.4417, 60.49996, 60.55803, 60.6159, 60.67357, 60.73104, 60.78831, 
    60.84539, 60.90226, 60.95892, 61.01538, 61.07164, 61.12769, 61.18353, 
    61.23915, 61.29457, 61.34978, 61.40477, 61.45955, 61.51411, 61.56845, 
    61.62257, 61.67648, 61.73016, 61.78362, 61.83686, 61.88987, 61.94265, 
    61.9952, 62.04753, 62.09962, 62.15149, 62.20312, 62.25451, 62.30567, 
    62.35659, 62.40727, 62.45771, 62.50792, 62.55787, 62.60759, 62.65705, 
    62.70627, 62.75525, 62.80397, 62.85244, 62.90065, 62.94862, 62.99633, 
    63.04378, 63.09097, 63.13791, 63.18458, 63.23099, 63.27714, 63.32302, 
    63.36863, 63.41398, 63.45906, 63.50386, 63.5484, 63.59266, 63.63664, 
    63.68035, 63.72378, 63.76693, 63.80981, 63.85239, 63.8947, 63.93672, 
    63.97845, 64.0199, 64.06105, 64.10192, 64.14249, 64.18277, 64.22276, 
    64.26244, 64.30183, 64.34093, 64.37972, 64.41821, 64.45639, 64.49428, 
    64.53185, 64.56911, 64.60608, 64.64272, 64.67906, 64.71508, 64.75079, 
    64.78619, 64.82126, 64.85602, 64.89046, 64.92458, 64.95837, 64.99184, 
    65.02498, 65.0578, 65.09029, 65.12245, 65.15428, 65.18578, 65.21695, 
    65.24778, 65.27827, 65.30843, 65.33826, 65.36774, 65.39687, 65.42567, 
    65.45413, 65.48225, 65.51001, 65.53743, 65.5645, 65.59122, 65.61759, 
    65.64362, 65.66928, 65.6946, 65.71956, 65.74416, 65.7684, 65.79229, 
    65.81582, 65.83899, 65.86179, 65.88424, 65.90632, 65.92804, 65.94939, 
    65.97038, 65.99099, 66.01124, 66.03112, 66.05063, 66.06977, 66.08853, 
    66.10693, 66.12495, 66.14259, 66.15986, 66.17675, 66.19327, 66.2094, 
    66.22516, 66.24054, 66.25554, 66.27015, 66.28439, 66.29824, 66.31171, 
    66.32479, 66.33749, 66.34981, 66.36174, 66.37328, 66.38445, 66.39521, 
    66.40559, 66.41559, 66.42519, 66.4344, 66.44323, 66.45166, 66.4597, 
    66.46735, 66.47462, 66.48148, 66.48796, 66.49404, 66.49973, 66.50503, 
    66.50993, 66.51444, 66.51855, 66.52228, 66.5256, 66.52853, 66.53107, 
    66.53322, 66.53497, 66.53632, 66.53727, 66.53783, 66.538, 66.53777, 
    66.53715, 66.53613, 66.53471, 66.53291, 66.5307, 66.5281, 66.5251, 
    66.52171, 66.51793, 66.51376, 66.50919, 66.50422, 66.49886, 66.4931, 
    66.48696, 66.48042, 66.4735, 66.46617, 66.45846, 66.45036, 66.44186, 
    66.43297, 66.4237, 66.41403, 66.40398, 66.39353, 66.38271, 66.37148, 
    66.35988, 66.34789, 66.33551, 66.32275, 66.3096, 66.29607, 66.28216, 
    66.26787, 66.25319, 66.23813, 66.22269, 66.20687, 66.19067, 66.1741, 
    66.15715, 66.13982, 66.12212, 66.10404, 66.08559, 66.06676, 66.04757, 
    66.028, 66.00806, 65.98775, 65.96708, 65.94604, 65.92463, 65.90285, 
    65.88071, 65.85822, 65.83535, 65.81213, 65.78854, 65.7646, 65.74029, 
    65.71563, 65.69061, 65.66525, 65.63952, 65.61345, 65.58702, 65.56024, 
    65.53311, 65.50564, 65.47782, 65.44965, 65.42114, 65.39229, 65.3631, 
    65.33356, 65.30369, 65.27348, 65.24293, 65.21204, 65.18082, 65.14927, 
    65.11739, 65.08517, 65.05263, 65.01976, 64.98656, 64.95304, 64.9192, 
    64.88503, 64.85054, 64.81573, 64.78061, 64.74516, 64.7094, 64.67333, 
    64.63695, 64.60025, 64.56324, 64.52592, 64.4883, 64.45037, 64.41214, 
    64.3736, 64.33476, 64.29562, 64.25619, 64.21645, 64.17642, 64.13609, 
    64.09547, 64.05457, 64.01336, 63.97187, 63.93009, 63.88803, 63.84568, 
    63.80304, 63.76013, 63.71693, 63.67346, 63.6297, 63.58567, 63.54137, 
    63.49679, 63.45194, 63.40683, 63.36143, 63.31578, 63.26986, 63.22367, 
    63.17721, 63.1305, 63.08352, 63.03629, 62.9888, 62.94105, 62.89304, 
    62.84478, 62.79628, 62.74751, 62.6985, 62.64924, 62.59974, 62.54998, 
    62.49999, 62.44975, 62.39927, 62.34855, 62.29759, 62.2464, 62.19497, 
    62.1433, 62.0914, 62.03927, 61.9869, 61.93431, 61.8815, 61.82845, 
    61.77518, 61.72168, 61.66796, 61.61403, 61.55987, 61.50549, 61.4509, 
    61.39609, 61.34106,
  55.53883, 55.60903, 55.67912, 55.74908, 55.81892, 55.88865, 55.95825, 
    56.02773, 56.09709, 56.16632, 56.23543, 56.30442, 56.37328, 56.44201, 
    56.5106, 56.57908, 56.64742, 56.71563, 56.78371, 56.85166, 56.91948, 
    56.98716, 57.0547, 57.12211, 57.18939, 57.25652, 57.32352, 57.39038, 
    57.45709, 57.52367, 57.5901, 57.65639, 57.72253, 57.78854, 57.85439, 
    57.9201, 57.98566, 58.05106, 58.11633, 58.18143, 58.24639, 58.3112, 
    58.37584, 58.44034, 58.50468, 58.56886, 58.63288, 58.69675, 58.76045, 
    58.824, 58.88738, 58.9506, 59.01365, 59.07654, 59.13926, 59.20182, 
    59.2642, 59.32642, 59.38847, 59.45034, 59.51204, 59.57357, 59.63492, 
    59.6961, 59.7571, 59.81792, 59.87856, 59.93901, 59.99929, 60.05939, 
    60.1193, 60.17902, 60.23856, 60.29791, 60.35707, 60.41605, 60.47483, 
    60.53342, 60.59181, 60.65001, 60.70801, 60.76582, 60.82343, 60.88083, 
    60.93804, 60.99504, 61.05185, 61.10844, 61.16483, 61.22102, 61.27699, 
    61.33275, 61.38831, 61.44365, 61.49878, 61.55369, 61.60838, 61.66286, 
    61.71712, 61.77116, 61.82498, 61.87858, 61.93195, 61.9851, 62.03801, 
    62.09071, 62.14317, 62.1954, 62.2474, 62.29916, 62.3507, 62.40199, 
    62.45304, 62.50386, 62.55444, 62.60478, 62.65487, 62.70472, 62.75432, 
    62.80368, 62.85279, 62.90165, 62.95025, 62.9986, 63.0467, 63.09454, 
    63.14213, 63.18946, 63.23653, 63.28333, 63.32988, 63.37616, 63.42217, 
    63.46792, 63.5134, 63.55861, 63.60355, 63.64822, 63.69261, 63.73672, 
    63.78056, 63.82413, 63.86741, 63.91041, 63.95313, 63.99556, 64.03771, 
    64.07957, 64.12115, 64.16243, 64.20342, 64.24412, 64.28453, 64.32464, 
    64.36445, 64.40397, 64.44318, 64.4821, 64.52071, 64.55902, 64.59702, 
    64.63472, 64.6721, 64.70918, 64.74596, 64.78241, 64.81855, 64.85438, 
    64.88988, 64.92508, 64.95995, 64.99451, 65.02874, 65.06264, 65.09623, 
    65.12949, 65.16241, 65.19501, 65.22729, 65.25922, 65.29083, 65.32211, 
    65.35304, 65.38364, 65.41391, 65.44383, 65.47342, 65.50266, 65.53156, 
    65.56011, 65.58833, 65.61619, 65.64371, 65.67088, 65.69769, 65.72416, 
    65.75027, 65.77603, 65.80144, 65.82648, 65.85117, 65.87551, 65.89948, 
    65.9231, 65.94635, 65.96925, 65.99177, 66.01393, 66.03573, 66.05716, 
    66.07822, 66.09892, 66.11924, 66.13919, 66.15878, 66.17798, 66.19682, 
    66.21528, 66.23337, 66.25108, 66.26841, 66.28536, 66.30194, 66.31814, 
    66.33395, 66.3494, 66.36445, 66.37912, 66.39341, 66.40732, 66.42084, 
    66.43398, 66.44672, 66.45908, 66.47106, 66.48265, 66.49385, 66.50466, 
    66.51508, 66.52511, 66.53475, 66.544, 66.55286, 66.56133, 66.5694, 
    66.57708, 66.58437, 66.59126, 66.59776, 66.60387, 66.60958, 66.6149, 
    66.61982, 66.62435, 66.62848, 66.63222, 66.63556, 66.6385, 66.64104, 
    66.6432, 66.64495, 66.64631, 66.64727, 66.64783, 66.64799, 66.64777, 
    66.64714, 66.64612, 66.6447, 66.64288, 66.64067, 66.63806, 66.63506, 
    66.63165, 66.62785, 66.62366, 66.61907, 66.61408, 66.6087, 66.60293, 
    66.59676, 66.5902, 66.58324, 66.57589, 66.56815, 66.56001, 66.55148, 
    66.54256, 66.53325, 66.52355, 66.51346, 66.50298, 66.4921, 66.48084, 
    66.46919, 66.45715, 66.44473, 66.43192, 66.41872, 66.40514, 66.39117, 
    66.37682, 66.36209, 66.34698, 66.33148, 66.31561, 66.29935, 66.28271, 
    66.26569, 66.2483, 66.23053, 66.21239, 66.19386, 66.17496, 66.1557, 
    66.13606, 66.11605, 66.09566, 66.07491, 66.05379, 66.0323, 66.01045, 
    65.98823, 65.96564, 65.9427, 65.91939, 65.89571, 65.87169, 65.8473, 
    65.82255, 65.79744, 65.77198, 65.74616, 65.71999, 65.69347, 65.6666, 
    65.63937, 65.61181, 65.58389, 65.55562, 65.52701, 65.49805, 65.46876, 
    65.43913, 65.40914, 65.37882, 65.34817, 65.31718, 65.28585, 65.2542, 
    65.2222, 65.18988, 65.15723, 65.12424, 65.09093, 65.0573, 65.02335, 
    64.98906, 64.95446, 64.91953, 64.88429, 64.84873, 64.81285, 64.77666, 
    64.74016, 64.70334, 64.66621, 64.62878, 64.59103, 64.55298, 64.51463, 
    64.47596, 64.437, 64.39774, 64.35818, 64.31831, 64.27815, 64.2377, 
    64.19695, 64.15591, 64.11459, 64.07297, 64.03106, 63.98887, 63.94639, 
    63.90363, 63.86058, 63.81725, 63.77365, 63.72976, 63.6856, 63.64117, 
    63.59646, 63.55148, 63.50623, 63.4607, 63.41491, 63.36885, 63.32253, 
    63.27595, 63.2291, 63.18199, 63.13462, 63.08699, 63.03911, 62.99097, 
    62.94258, 62.89393, 62.84504, 62.79589, 62.74649, 62.69685, 62.64697, 
    62.59683, 62.54646, 62.49584, 62.44498, 62.39389, 62.34256, 62.29099, 
    62.23919, 62.18715, 62.13488, 62.08239, 62.02966, 61.9767, 61.92352, 
    61.87011, 61.81648, 61.76263, 61.70856, 61.65426, 61.59975, 61.54502, 
    61.49007, 61.43491,
  55.621, 55.69131, 55.7615, 55.83158, 55.90153, 55.97137, 56.04108, 
    56.11067, 56.18014, 56.24949, 56.31871, 56.3878, 56.45678, 56.52562, 
    56.59433, 56.66292, 56.73138, 56.79971, 56.8679, 56.93597, 57.00389, 
    57.07169, 57.13936, 57.20688, 57.27428, 57.34153, 57.40864, 57.47562, 
    57.54245, 57.60915, 57.6757, 57.74211, 57.80838, 57.8745, 57.94048, 
    58.0063, 58.07198, 58.13752, 58.2029, 58.26813, 58.33321, 58.39814, 
    58.46291, 58.52753, 58.592, 58.6563, 58.72045, 58.78444, 58.84827, 
    58.91195, 58.97545, 59.0388, 59.10198, 59.165, 59.22784, 59.29053, 
    59.35304, 59.41539, 59.47757, 59.53957, 59.6014, 59.66306, 59.72454, 
    59.78585, 59.84697, 59.90792, 59.9687, 60.02929, 60.0897, 60.14993, 
    60.20997, 60.26982, 60.3295, 60.38898, 60.44828, 60.50738, 60.5663, 
    60.62502, 60.68354, 60.74188, 60.80001, 60.85796, 60.9157, 60.97324, 
    61.03058, 61.08772, 61.14466, 61.20139, 61.25792, 61.31424, 61.37035, 
    61.42625, 61.48193, 61.53741, 61.59268, 61.64772, 61.70256, 61.75718, 
    61.81157, 61.86575, 61.9197, 61.97343, 62.02694, 62.08023, 62.13328, 
    62.18611, 62.23871, 62.29108, 62.34321, 62.39511, 62.44678, 62.49821, 
    62.54941, 62.60036, 62.65108, 62.70155, 62.75178, 62.80177, 62.85151, 
    62.901, 62.95024, 62.99923, 63.04798, 63.09647, 63.1447, 63.19268, 
    63.2404, 63.28786, 63.33507, 63.38201, 63.42869, 63.4751, 63.52125, 
    63.56713, 63.61275, 63.65809, 63.70316, 63.74796, 63.79248, 63.83673, 
    63.8807, 63.9244, 63.96781, 64.01094, 64.05379, 64.09635, 64.13863, 
    64.18063, 64.22233, 64.26374, 64.30486, 64.34569, 64.38622, 64.42646, 
    64.4664, 64.50603, 64.54538, 64.58442, 64.62315, 64.66158, 64.69971, 
    64.73753, 64.77504, 64.81224, 64.84913, 64.8857, 64.92197, 64.95791, 
    64.99354, 65.02885, 65.06384, 65.0985, 65.13285, 65.16688, 65.20057, 
    65.23394, 65.26698, 65.2997, 65.33208, 65.36413, 65.39584, 65.42722, 
    65.45827, 65.48898, 65.51935, 65.54938, 65.57906, 65.60841, 65.63741, 
    65.66607, 65.69437, 65.72234, 65.74995, 65.77722, 65.80413, 65.83069, 
    65.8569, 65.88275, 65.90825, 65.93339, 65.95817, 65.98259, 66.00665, 
    66.03036, 66.0537, 66.07667, 66.09928, 66.12152, 66.1434, 66.16491, 
    66.18605, 66.20682, 66.22722, 66.24725, 66.2669, 66.28618, 66.30509, 
    66.32362, 66.34177, 66.35955, 66.37695, 66.39397, 66.41061, 66.42686, 
    66.44275, 66.45824, 66.47335, 66.48808, 66.50243, 66.51638, 66.52995, 
    66.54314, 66.55594, 66.56835, 66.58038, 66.592, 66.60325, 66.6141, 
    66.62457, 66.63464, 66.64431, 66.65359, 66.66249, 66.67099, 66.67909, 
    66.68681, 66.69412, 66.70104, 66.70757, 66.7137, 66.71944, 66.72477, 
    66.72971, 66.73426, 66.7384, 66.74216, 66.74551, 66.74846, 66.75101, 
    66.75317, 66.75494, 66.7563, 66.75726, 66.75783, 66.758, 66.75777, 
    66.75714, 66.75611, 66.75468, 66.75286, 66.75064, 66.74802, 66.745, 
    66.74158, 66.73778, 66.73357, 66.72896, 66.72395, 66.71855, 66.71275, 
    66.70657, 66.69997, 66.69299, 66.68561, 66.67784, 66.66967, 66.66111, 
    66.65215, 66.64281, 66.63306, 66.62293, 66.61241, 66.60149, 66.59019, 
    66.5785, 66.56641, 66.55394, 66.54108, 66.52783, 66.5142, 66.50018, 
    66.48578, 66.47099, 66.45582, 66.44026, 66.42432, 66.408, 66.3913, 
    66.37422, 66.35677, 66.33893, 66.32071, 66.30212, 66.28316, 66.26382, 
    66.2441, 66.22401, 66.20356, 66.18273, 66.16153, 66.13996, 66.11803, 
    66.09573, 66.07306, 66.05003, 66.02663, 66.00288, 65.97875, 65.95428, 
    65.92944, 65.90424, 65.87868, 65.85278, 65.82652, 65.7999, 65.77293, 
    65.74561, 65.71794, 65.68992, 65.66155, 65.63284, 65.60379, 65.57439, 
    65.54465, 65.51456, 65.48414, 65.45338, 65.42228, 65.39085, 65.35908, 
    65.32697, 65.29454, 65.26178, 65.22868, 65.19526, 65.16151, 65.12744, 
    65.09304, 65.05833, 65.02328, 64.98792, 64.95225, 64.91625, 64.87994, 
    64.84332, 64.80637, 64.76913, 64.73157, 64.6937, 64.65553, 64.61705, 
    64.57826, 64.53918, 64.49979, 64.4601, 64.42011, 64.37983, 64.33925, 
    64.29837, 64.25721, 64.21575, 64.174, 64.13197, 64.08964, 64.04703, 
    64.00414, 63.96096, 63.9175, 63.87377, 63.82975, 63.78546, 63.74089, 
    63.69605, 63.65094, 63.60555, 63.55989, 63.51397, 63.46778, 63.42132, 
    63.3746, 63.32762, 63.28037, 63.23287, 63.18511, 63.13709, 63.08881, 
    63.04028, 62.9915, 62.94247, 62.89318, 62.84365, 62.79388, 62.74385, 
    62.69358, 62.64307, 62.59232, 62.54133, 62.4901, 62.43863, 62.38692, 
    62.33498, 62.28281, 62.2304, 62.17777, 62.1249, 62.07181, 62.01849, 
    61.96495, 61.91118, 61.85719, 61.80298, 61.74855, 61.6939, 61.63903, 
    61.58395, 61.52865,
  55.70303, 55.77345, 55.84375, 55.91394, 55.984, 56.05395, 56.12377, 
    56.19347, 56.26305, 56.33251, 56.40185, 56.47105, 56.54014, 56.6091, 
    56.67793, 56.74663, 56.8152, 56.88364, 56.95195, 57.02013, 57.08818, 
    57.1561, 57.22388, 57.29152, 57.35903, 57.4264, 57.49363, 57.56073, 
    57.62769, 57.6945, 57.76117, 57.8277, 57.89409, 57.96033, 58.02643, 
    58.09238, 58.15818, 58.22384, 58.28934, 58.3547, 58.4199, 58.48495, 
    58.54985, 58.6146, 58.67918, 58.74362, 58.80789, 58.87201, 58.93597, 
    58.99976, 59.0634, 59.12687, 59.19018, 59.25333, 59.3163, 59.37912, 
    59.44176, 59.50423, 59.56654, 59.62867, 59.69064, 59.75242, 59.81403, 
    59.87547, 59.93673, 59.99781, 60.05872, 60.11944, 60.17999, 60.24034, 
    60.30052, 60.36051, 60.42031, 60.47993, 60.53936, 60.5986, 60.65765, 
    60.7165, 60.77517, 60.83363, 60.89191, 60.94998, 61.00786, 61.06554, 
    61.12301, 61.18029, 61.23736, 61.29423, 61.35089, 61.40734, 61.46359, 
    61.51963, 61.57545, 61.63107, 61.68647, 61.74166, 61.79663, 61.85138, 
    61.90591, 61.96023, 62.01432, 62.06819, 62.12183, 62.17525, 62.22845, 
    62.28141, 62.33415, 62.38666, 62.43893, 62.49097, 62.54278, 62.59435, 
    62.64568, 62.69677, 62.74762, 62.79823, 62.8486, 62.89872, 62.9486, 
    62.99823, 63.04761, 63.09674, 63.14561, 63.19424, 63.24261, 63.29073, 
    63.33858, 63.38618, 63.43352, 63.4806, 63.52741, 63.57396, 63.62025, 
    63.66626, 63.71201, 63.75749, 63.80269, 63.84763, 63.89228, 63.93666, 
    63.98077, 64.0246, 64.06814, 64.1114, 64.15438, 64.19707, 64.23949, 
    64.28161, 64.32344, 64.36498, 64.40623, 64.44719, 64.48785, 64.52821, 
    64.56828, 64.60805, 64.64751, 64.68668, 64.72554, 64.76409, 64.80235, 
    64.84029, 64.87792, 64.91524, 64.95225, 64.98895, 65.02533, 65.06139, 
    65.09714, 65.13257, 65.16767, 65.20246, 65.23692, 65.27106, 65.30487, 
    65.33836, 65.37151, 65.40434, 65.43682, 65.46899, 65.50081, 65.5323, 
    65.56345, 65.59427, 65.62474, 65.65488, 65.68467, 65.71412, 65.74323, 
    65.77198, 65.80039, 65.82845, 65.85617, 65.88353, 65.91054, 65.93719, 
    65.9635, 65.98945, 66.01504, 66.04027, 66.06514, 66.08965, 66.1138, 
    66.13759, 66.16101, 66.18407, 66.20676, 66.22909, 66.25105, 66.27264, 
    66.29385, 66.3147, 66.33518, 66.35529, 66.37502, 66.39436, 66.41335, 
    66.43195, 66.45016, 66.46801, 66.48547, 66.50256, 66.51926, 66.53558, 
    66.55152, 66.56708, 66.58224, 66.59703, 66.61143, 66.62544, 66.63907, 
    66.65231, 66.66515, 66.67761, 66.68968, 66.70135, 66.71265, 66.72354, 
    66.73404, 66.74415, 66.75387, 66.76318, 66.77212, 66.78065, 66.78878, 
    66.79652, 66.80387, 66.81082, 66.81737, 66.82352, 66.82928, 66.83464, 
    66.8396, 66.84416, 66.84833, 66.85209, 66.85546, 66.85842, 66.86099, 
    66.86316, 66.86493, 66.86629, 66.86726, 66.86783, 66.868, 66.86777, 
    66.86713, 66.8661, 66.86467, 66.86284, 66.86061, 66.85798, 66.85495, 
    66.85152, 66.84769, 66.84347, 66.83884, 66.83382, 66.8284, 66.82258, 
    66.81636, 66.80975, 66.80273, 66.79533, 66.78752, 66.77932, 66.77073, 
    66.76174, 66.75236, 66.74258, 66.73241, 66.72184, 66.71088, 66.69954, 
    66.6878, 66.67567, 66.66315, 66.65024, 66.63694, 66.62325, 66.60918, 
    66.59472, 66.57987, 66.56464, 66.54903, 66.53303, 66.51665, 66.49989, 
    66.48274, 66.46522, 66.44731, 66.42902, 66.41037, 66.39133, 66.37192, 
    66.35213, 66.33196, 66.31143, 66.29053, 66.26925, 66.2476, 66.22559, 
    66.2032, 66.18045, 66.15733, 66.13385, 66.11001, 66.0858, 66.06123, 
    66.0363, 66.01101, 65.98537, 65.95937, 65.93301, 65.9063, 65.87923, 
    65.85181, 65.82404, 65.79592, 65.76746, 65.73864, 65.70948, 65.67998, 
    65.65013, 65.61994, 65.58942, 65.55855, 65.52734, 65.4958, 65.46392, 
    65.43171, 65.39916, 65.36629, 65.33308, 65.29955, 65.26568, 65.23149, 
    65.19698, 65.16214, 65.12698, 65.09151, 65.05571, 65.01959, 64.98316, 
    64.94642, 64.90936, 64.87199, 64.8343, 64.79632, 64.75802, 64.71941, 
    64.6805, 64.64129, 64.60178, 64.56196, 64.52185, 64.48144, 64.44073, 
    64.39973, 64.35843, 64.31684, 64.27496, 64.2328, 64.19035, 64.14761, 
    64.10458, 64.06127, 64.01768, 63.97381, 63.92966, 63.88524, 63.84054, 
    63.79556, 63.75031, 63.70479, 63.659, 63.61294, 63.56662, 63.52003, 
    63.47317, 63.42605, 63.37867, 63.33103, 63.28313, 63.23498, 63.18657, 
    63.1379, 63.08898, 63.03981, 62.99039, 62.94072, 62.89081, 62.84065, 
    62.79024, 62.73959, 62.68871, 62.63757, 62.5862, 62.5346, 62.48275, 
    62.43068, 62.37837, 62.32582, 62.27305, 62.22005, 62.16682, 62.11337, 
    62.05968, 62.00578, 61.95165, 61.8973, 61.84273, 61.78794, 61.73294, 
    61.67772, 61.62229,
  55.78492, 55.85545, 55.92587, 55.99616, 56.06633, 56.13639, 56.20633, 
    56.27614, 56.34583, 56.4154, 56.48485, 56.55417, 56.62337, 56.69244, 
    56.76138, 56.8302, 56.89889, 56.96745, 57.03587, 57.10417, 57.17233, 
    57.24036, 57.30826, 57.37602, 57.44365, 57.51114, 57.57849, 57.64571, 
    57.71278, 57.77972, 57.84651, 57.91316, 57.97967, 58.04603, 58.11225, 
    58.17833, 58.24425, 58.31003, 58.37566, 58.44114, 58.50646, 58.57164, 
    58.63666, 58.70153, 58.76625, 58.8308, 58.89521, 58.95945, 59.02353, 
    59.08746, 59.15122, 59.21482, 59.27826, 59.34153, 59.40464, 59.46758, 
    59.53035, 59.59296, 59.65539, 59.71766, 59.77975, 59.84166, 59.90341, 
    59.96498, 60.02637, 60.08758, 60.14862, 60.20947, 60.27015, 60.33064, 
    60.39095, 60.45107, 60.51101, 60.57076, 60.63033, 60.6897, 60.74888, 
    60.80787, 60.86667, 60.92527, 60.98368, 61.04189, 61.0999, 61.15772, 
    61.21533, 61.27274, 61.32995, 61.38696, 61.44375, 61.50035, 61.55673, 
    61.6129, 61.66887, 61.72462, 61.78016, 61.83548, 61.89059, 61.94548, 
    62.00015, 62.0546, 62.10883, 62.16284, 62.21663, 62.27018, 62.32352, 
    62.37662, 62.42949, 62.48214, 62.53455, 62.58673, 62.63867, 62.69038, 
    62.74185, 62.79308, 62.84407, 62.89482, 62.94532, 62.99558, 63.0456, 
    63.09536, 63.14488, 63.19415, 63.24316, 63.29193, 63.34044, 63.38869, 
    63.43668, 63.48442, 63.53189, 63.57911, 63.62606, 63.67274, 63.71916, 
    63.76531, 63.8112, 63.85681, 63.90215, 63.94722, 63.99201, 64.03652, 
    64.08076, 64.12472, 64.1684, 64.21179, 64.25491, 64.29773, 64.34027, 
    64.38252, 64.42448, 64.46616, 64.50754, 64.54862, 64.58941, 64.62991, 
    64.6701, 64.70999, 64.74959, 64.78888, 64.82787, 64.86655, 64.90492, 
    64.94299, 64.98074, 65.01819, 65.05532, 65.09213, 65.12864, 65.16483, 
    65.20069, 65.23624, 65.27146, 65.30637, 65.34094, 65.3752, 65.40912, 
    65.44272, 65.47599, 65.50893, 65.54153, 65.5738, 65.60574, 65.63734, 
    65.6686, 65.69952, 65.7301, 65.76035, 65.79025, 65.81979, 65.84901, 
    65.87786, 65.90638, 65.93454, 65.96235, 65.98981, 66.01692, 66.04367, 
    66.07007, 66.09612, 66.1218, 66.14712, 66.17208, 66.19669, 66.22092, 
    66.2448, 66.26831, 66.29145, 66.31423, 66.33664, 66.35868, 66.38035, 
    66.40165, 66.42257, 66.44312, 66.4633, 66.48311, 66.50253, 66.52158, 
    66.54025, 66.55855, 66.57646, 66.59399, 66.61114, 66.62791, 66.64429, 
    66.66029, 66.6759, 66.69113, 66.70597, 66.72043, 66.7345, 66.74817, 
    66.76146, 66.77436, 66.78687, 66.79898, 66.8107, 66.82204, 66.83297, 
    66.84351, 66.85366, 66.86342, 66.87277, 66.88174, 66.8903, 66.89847, 
    66.90624, 66.91362, 66.92059, 66.92717, 66.93335, 66.93913, 66.94451, 
    66.94949, 66.95407, 66.95825, 66.96203, 66.96541, 66.96838, 66.97096, 
    66.97314, 66.97491, 66.97629, 66.97726, 66.97783, 66.978, 66.97777, 
    66.97713, 66.9761, 66.97466, 66.97282, 66.97058, 66.96794, 66.9649, 
    66.96146, 66.95762, 66.95337, 66.94873, 66.94369, 66.93824, 66.9324, 
    66.92616, 66.91952, 66.91248, 66.90504, 66.89721, 66.88898, 66.88035, 
    66.87132, 66.8619, 66.85208, 66.84187, 66.83127, 66.82027, 66.80888, 
    66.79709, 66.78491, 66.77235, 66.75938, 66.74603, 66.73229, 66.71817, 
    66.70365, 66.68875, 66.67346, 66.65778, 66.64172, 66.62528, 66.60845, 
    66.59124, 66.57365, 66.55568, 66.53732, 66.51859, 66.49949, 66.48, 
    66.46014, 66.4399, 66.41929, 66.3983, 66.37695, 66.35522, 66.33311, 
    66.31065, 66.28781, 66.26461, 66.24104, 66.21711, 66.19282, 66.16816, 
    66.14314, 66.11775, 66.09202, 66.06592, 66.03947, 66.01266, 65.9855, 
    65.95798, 65.93011, 65.90189, 65.87332, 65.84441, 65.81515, 65.78554, 
    65.75558, 65.72529, 65.69466, 65.66367, 65.63236, 65.60071, 65.56872, 
    65.53639, 65.50374, 65.47075, 65.43742, 65.40378, 65.3698, 65.33549, 
    65.30087, 65.26591, 65.23064, 65.19504, 65.15912, 65.12289, 65.08633, 
    65.04946, 65.01228, 64.97479, 64.93698, 64.89887, 64.86044, 64.82172, 
    64.78268, 64.74334, 64.7037, 64.66376, 64.62352, 64.58298, 64.54214, 
    64.50101, 64.45959, 64.41787, 64.37586, 64.33356, 64.29098, 64.2481, 
    64.20495, 64.16151, 64.11778, 64.07378, 64.0295, 63.98494, 63.94011, 
    63.895, 63.84961, 63.80396, 63.75803, 63.71184, 63.66537, 63.61865, 
    63.57166, 63.5244, 63.47689, 63.42911, 63.38107, 63.33278, 63.28423, 
    63.23543, 63.18637, 63.13707, 63.08751, 63.0377, 62.98765, 62.93735, 
    62.88681, 62.83602, 62.78499, 62.73372, 62.68222, 62.63047, 62.57849, 
    62.52628, 62.47383, 62.42115, 62.36824, 62.31509, 62.26173, 62.20813, 
    62.15431, 62.10027, 62.04601, 61.99152, 61.93681, 61.88189, 61.82674, 
    61.77139, 61.71581,
  55.86668, 55.93732, 56.00784, 56.07824, 56.14853, 56.21869, 56.28874, 
    56.35867, 56.42847, 56.49815, 56.56771, 56.63715, 56.70646, 56.77564, 
    56.8447, 56.91363, 56.98244, 57.05111, 57.11965, 57.18806, 57.25635, 
    57.32449, 57.39251, 57.46039, 57.52813, 57.59575, 57.66322, 57.73055, 
    57.79774, 57.8648, 57.93171, 57.99849, 58.06511, 58.1316, 58.19794, 
    58.26414, 58.33018, 58.39608, 58.46184, 58.52744, 58.59289, 58.6582, 
    58.72334, 58.78834, 58.85318, 58.91786, 58.98239, 59.04676, 59.11097, 
    59.17502, 59.23891, 59.30264, 59.3662, 59.42961, 59.49284, 59.55591, 
    59.61882, 59.68155, 59.74411, 59.80651, 59.86873, 59.93078, 59.99266, 
    60.05436, 60.11588, 60.17723, 60.2384, 60.29939, 60.36019, 60.42082, 
    60.48126, 60.54152, 60.60159, 60.66147, 60.72117, 60.78068, 60.84, 
    60.89912, 60.95806, 61.0168, 61.07534, 61.13369, 61.19183, 61.24979, 
    61.30753, 61.36508, 61.42243, 61.47957, 61.53651, 61.59324, 61.64976, 
    61.70607, 61.76217, 61.81806, 61.87374, 61.9292, 61.98444, 62.03947, 
    62.09428, 62.14887, 62.20324, 62.25739, 62.31131, 62.36501, 62.41848, 
    62.47172, 62.52473, 62.57752, 62.63007, 62.68239, 62.73447, 62.78632, 
    62.83792, 62.88929, 62.94042, 62.99131, 63.04195, 63.09235, 63.14251, 
    63.19241, 63.24207, 63.29147, 63.34063, 63.38953, 63.43817, 63.48656, 
    63.53469, 63.58257, 63.63018, 63.67753, 63.72462, 63.77144, 63.818, 
    63.86428, 63.9103, 63.95605, 64.00153, 64.04673, 64.09165, 64.13631, 
    64.18068, 64.22477, 64.26858, 64.31211, 64.35535, 64.39831, 64.44099, 
    64.48337, 64.52546, 64.56726, 64.60877, 64.64999, 64.69091, 64.73153, 
    64.77185, 64.81187, 64.85159, 64.89101, 64.93013, 64.96893, 65.00743, 
    65.04562, 65.0835, 65.12107, 65.15833, 65.19527, 65.2319, 65.2682, 
    65.30418, 65.33985, 65.3752, 65.41022, 65.44492, 65.47929, 65.51333, 
    65.54704, 65.58042, 65.61347, 65.64619, 65.67857, 65.71062, 65.74233, 
    65.7737, 65.80473, 65.83543, 65.86578, 65.89577, 65.92544, 65.95475, 
    65.98371, 66.01233, 66.04059, 66.0685, 66.09606, 66.12327, 66.15012, 
    66.17661, 66.20275, 66.22852, 66.25394, 66.279, 66.30369, 66.32802, 
    66.35198, 66.37558, 66.39881, 66.42167, 66.44417, 66.46629, 66.48804, 
    66.50941, 66.53042, 66.55105, 66.5713, 66.59119, 66.61069, 66.62981, 
    66.64855, 66.66691, 66.68489, 66.70249, 66.7197, 66.73653, 66.75298, 
    66.76904, 66.78472, 66.8, 66.8149, 66.82941, 66.84354, 66.85727, 
    66.87061, 66.88355, 66.89611, 66.90827, 66.92004, 66.93142, 66.9424, 
    66.95298, 66.96317, 66.97296, 66.98236, 66.99136, 66.99995, 67.00816, 
    67.01596, 67.02336, 67.03036, 67.03697, 67.04317, 67.04897, 67.05437, 
    67.05938, 67.06397, 67.06817, 67.07197, 67.07536, 67.07835, 67.08093, 
    67.08312, 67.0849, 67.08628, 67.08726, 67.08783, 67.088, 67.08777, 
    67.08713, 67.08609, 67.08465, 67.0828, 67.08055, 67.0779, 67.07484, 
    67.0714, 67.06754, 67.06327, 67.05861, 67.05355, 67.04808, 67.04222, 
    67.03595, 67.02928, 67.02222, 67.01475, 67.00689, 66.99862, 66.98996, 
    66.9809, 66.97144, 66.96159, 66.95133, 66.94069, 66.92964, 66.91821, 
    66.90638, 66.89415, 66.88153, 66.86852, 66.85513, 66.84133, 66.82715, 
    66.81258, 66.79762, 66.78226, 66.76653, 66.7504, 66.7339, 66.71701, 
    66.69973, 66.68208, 66.66403, 66.64561, 66.62681, 66.60763, 66.58807, 
    66.56813, 66.54781, 66.52712, 66.50606, 66.48462, 66.46281, 66.44063, 
    66.41808, 66.39516, 66.37187, 66.34821, 66.3242, 66.2998, 66.27505, 
    66.24995, 66.22447, 66.19864, 66.17245, 66.1459, 66.11899, 66.09173, 
    66.06411, 66.03614, 66.00782, 65.97916, 65.95013, 65.92077, 65.89105, 
    65.86099, 65.8306, 65.79985, 65.76876, 65.73734, 65.70557, 65.67348, 
    65.64104, 65.60827, 65.57516, 65.54173, 65.50797, 65.47387, 65.43945, 
    65.4047, 65.36963, 65.33423, 65.29852, 65.26247, 65.22612, 65.18945, 
    65.15246, 65.11515, 65.07754, 65.0396, 65.00137, 64.96281, 64.92396, 
    64.8848, 64.84534, 64.80556, 64.7655, 64.72512, 64.68446, 64.64349, 
    64.60223, 64.56067, 64.51882, 64.47668, 64.43425, 64.39153, 64.34853, 
    64.30524, 64.26167, 64.21781, 64.17368, 64.12926, 64.08456, 64.0396, 
    63.99435, 63.94883, 63.90304, 63.85698, 63.81065, 63.76405, 63.71719, 
    63.67006, 63.62267, 63.57501, 63.5271, 63.47892, 63.4305, 63.38181, 
    63.33287, 63.28367, 63.23423, 63.18453, 63.13459, 63.0844, 63.03396, 
    62.98328, 62.93235, 62.88118, 62.82978, 62.77813, 62.72625, 62.67413, 
    62.62177, 62.56919, 62.51637, 62.46331, 62.41004, 62.35653, 62.3028, 
    62.24884, 62.19466, 62.14025, 62.08563, 62.03078, 61.97572, 61.92044, 
    61.86494, 61.80923,
  55.9483, 56.01904, 56.08967, 56.16019, 56.23058, 56.30086, 56.37102, 
    56.44106, 56.51097, 56.58077, 56.65044, 56.71999, 56.78941, 56.85871, 
    56.92788, 56.99693, 57.06585, 57.13464, 57.2033, 57.27182, 57.34022, 
    57.40849, 57.47662, 57.54462, 57.61248, 57.68021, 57.7478, 57.81525, 
    57.88257, 57.94975, 58.01678, 58.08367, 58.15042, 58.21703, 58.2835, 
    58.34981, 58.41599, 58.48201, 58.54789, 58.61361, 58.67919, 58.74461, 
    58.80989, 58.87501, 58.93998, 59.00478, 59.06944, 59.13394, 59.19828, 
    59.26245, 59.32647, 59.39033, 59.45403, 59.51756, 59.58092, 59.64412, 
    59.70715, 59.77002, 59.83271, 59.89524, 59.95759, 60.01977, 60.08178, 
    60.14361, 60.20527, 60.26675, 60.32805, 60.38917, 60.45011, 60.51087, 
    60.57145, 60.63184, 60.69204, 60.75206, 60.8119, 60.87154, 60.93099, 
    60.99026, 61.04932, 61.1082, 61.16688, 61.22536, 61.28365, 61.34174, 
    61.39962, 61.45731, 61.51479, 61.57207, 61.62915, 61.68601, 61.74267, 
    61.79912, 61.85536, 61.91139, 61.96721, 62.0228, 62.07819, 62.13336, 
    62.18831, 62.24304, 62.29755, 62.35183, 62.40589, 62.45973, 62.51334, 
    62.56672, 62.61988, 62.6728, 62.72549, 62.77795, 62.83017, 62.88215, 
    62.9339, 62.98541, 63.03668, 63.0877, 63.13849, 63.18903, 63.23932, 
    63.28936, 63.33916, 63.3887, 63.438, 63.48703, 63.53582, 63.58435, 
    63.63262, 63.68063, 63.72838, 63.77587, 63.82309, 63.87005, 63.91674, 
    63.96317, 64.00932, 64.05521, 64.10082, 64.14616, 64.19122, 64.23601, 
    64.28052, 64.32474, 64.36868, 64.41235, 64.45573, 64.49882, 64.54163, 
    64.58414, 64.62637, 64.6683, 64.70995, 64.75129, 64.79234, 64.83309, 
    64.87354, 64.9137, 64.95354, 64.99309, 65.03233, 65.07127, 65.10989, 
    65.14821, 65.18621, 65.22391, 65.26128, 65.29835, 65.33509, 65.37152, 
    65.40763, 65.44341, 65.47888, 65.51402, 65.54884, 65.58332, 65.61749, 
    65.65131, 65.68481, 65.71798, 65.75081, 65.7833, 65.81547, 65.84728, 
    65.87877, 65.90991, 65.9407, 65.97116, 66.00127, 66.03104, 66.06046, 
    66.08952, 66.11824, 66.14661, 66.17462, 66.20228, 66.22958, 66.25653, 
    66.28313, 66.30936, 66.33523, 66.36074, 66.38589, 66.41067, 66.43509, 
    66.45914, 66.48283, 66.50614, 66.52909, 66.55167, 66.57388, 66.59571, 
    66.61716, 66.63825, 66.65896, 66.67929, 66.69924, 66.71882, 66.73801, 
    66.75683, 66.77526, 66.79331, 66.81097, 66.82826, 66.84515, 66.86166, 
    66.87779, 66.89352, 66.90887, 66.92383, 66.93839, 66.95257, 66.96635, 
    66.97974, 66.99274, 67.00535, 67.01756, 67.02937, 67.04079, 67.05182, 
    67.06245, 67.07268, 67.0825, 67.09193, 67.10097, 67.1096, 67.11784, 
    67.12567, 67.1331, 67.14014, 67.14677, 67.15299, 67.15882, 67.16424, 
    67.16926, 67.17388, 67.17809, 67.1819, 67.18531, 67.18831, 67.19091, 
    67.1931, 67.19489, 67.19627, 67.19725, 67.19783, 67.198, 67.19776, 
    67.19713, 67.19608, 67.19463, 67.19278, 67.19052, 67.18786, 67.1848, 
    67.18133, 67.17745, 67.17317, 67.1685, 67.16341, 67.15792, 67.15204, 
    67.14574, 67.13905, 67.13196, 67.12446, 67.11656, 67.10827, 67.09957, 
    67.09047, 67.08098, 67.07108, 67.06079, 67.0501, 67.03902, 67.02753, 
    67.01566, 67.00338, 66.99072, 66.97765, 66.9642, 66.95036, 66.93612, 
    66.92149, 66.90647, 66.89106, 66.87527, 66.85908, 66.84251, 66.82555, 
    66.80821, 66.79048, 66.77237, 66.75388, 66.735, 66.71575, 66.69611, 
    66.6761, 66.65571, 66.63494, 66.6138, 66.59228, 66.57039, 66.54813, 
    66.52549, 66.50248, 66.4791, 66.45536, 66.43125, 66.40678, 66.38194, 
    66.35673, 66.33116, 66.30523, 66.27895, 66.2523, 66.22529, 66.19793, 
    66.17021, 66.14214, 66.11372, 66.08495, 66.05582, 66.02635, 65.99654, 
    65.96637, 65.93586, 65.90501, 65.87381, 65.84228, 65.8104, 65.77818, 
    65.74564, 65.71275, 65.67953, 65.64598, 65.6121, 65.57789, 65.54335, 
    65.50848, 65.47329, 65.43777, 65.40194, 65.36578, 65.3293, 65.2925, 
    65.25539, 65.21796, 65.18022, 65.14217, 65.1038, 65.06512, 65.02615, 
    64.98685, 64.94726, 64.90736, 64.86716, 64.82666, 64.78587, 64.74477, 
    64.70338, 64.66169, 64.61971, 64.57744, 64.53487, 64.49202, 64.44888, 
    64.40546, 64.36176, 64.31776, 64.27349, 64.22894, 64.18411, 64.13901, 
    64.09363, 64.04797, 64.00204, 63.95584, 63.90938, 63.86264, 63.81564, 
    63.76838, 63.72084, 63.67305, 63.625, 63.57669, 63.52812, 63.47929, 
    63.43021, 63.38088, 63.3313, 63.28146, 63.23138, 63.18105, 63.13047, 
    63.07965, 63.02858, 62.97728, 62.92573, 62.87395, 62.82192, 62.76966, 
    62.71717, 62.66444, 62.61148, 62.55829, 62.50488, 62.45123, 62.39736, 
    62.34326, 62.28894, 62.23439, 62.17963, 62.12465, 62.06944, 62.01402, 
    61.95839, 61.90254,
  56.02977, 56.10062, 56.17137, 56.24199, 56.3125, 56.38288, 56.45316, 
    56.5233, 56.59333, 56.66324, 56.73302, 56.80269, 56.87223, 56.94164, 
    57.01093, 57.08009, 57.14912, 57.21803, 57.2868, 57.35545, 57.42396, 
    57.49234, 57.5606, 57.62871, 57.69669, 57.76454, 57.83225, 57.89983, 
    57.96726, 58.03456, 58.10171, 58.16873, 58.2356, 58.30233, 58.36892, 
    58.43536, 58.50165, 58.5678, 58.6338, 58.69965, 58.76535, 58.8309, 
    58.8963, 58.96155, 59.02664, 59.09158, 59.15636, 59.22098, 59.28545, 
    59.34976, 59.4139, 59.47789, 59.54171, 59.60537, 59.66887, 59.7322, 
    59.79536, 59.85836, 59.92118, 59.98384, 60.04633, 60.10863, 60.17078, 
    60.23274, 60.29453, 60.35614, 60.41758, 60.47883, 60.53991, 60.6008, 
    60.66151, 60.72204, 60.78238, 60.84253, 60.9025, 60.96228, 61.02187, 
    61.08127, 61.14047, 61.19949, 61.2583, 61.31693, 61.37535, 61.43357, 
    61.4916, 61.54942, 61.60704, 61.66446, 61.72167, 61.77868, 61.83547, 
    61.89206, 61.94844, 62.00461, 62.06056, 62.1163, 62.17183, 62.22713, 
    62.28222, 62.33709, 62.39174, 62.44617, 62.50037, 62.55434, 62.6081, 
    62.66162, 62.71491, 62.76797, 62.8208, 62.8734, 62.92577, 62.97789, 
    63.02978, 63.08143, 63.13284, 63.18401, 63.23493, 63.28561, 63.33604, 
    63.38622, 63.43616, 63.48584, 63.53527, 63.58445, 63.63338, 63.68204, 
    63.73045, 63.7786, 63.82649, 63.87412, 63.92148, 63.96858, 64.01541, 
    64.06197, 64.10827, 64.15429, 64.20004, 64.24551, 64.29071, 64.33563, 
    64.38027, 64.42464, 64.46872, 64.51251, 64.55603, 64.59926, 64.6422, 
    64.68484, 64.7272, 64.76927, 64.81104, 64.85252, 64.8937, 64.93459, 
    64.97517, 65.01545, 65.05543, 65.0951, 65.13447, 65.17353, 65.21229, 
    65.25072, 65.28886, 65.32668, 65.36418, 65.40137, 65.43824, 65.47479, 
    65.51102, 65.54693, 65.58251, 65.61777, 65.65271, 65.68732, 65.72159, 
    65.75554, 65.78915, 65.82243, 65.85538, 65.88799, 65.92027, 65.95219, 
    65.98379, 66.01505, 66.04595, 66.07652, 66.10674, 66.1366, 66.16613, 
    66.1953, 66.22412, 66.25259, 66.28071, 66.30846, 66.33587, 66.36292, 
    66.38961, 66.41593, 66.4419, 66.46751, 66.49274, 66.51762, 66.54214, 
    66.56628, 66.59005, 66.61346, 66.63649, 66.65915, 66.68144, 66.70335, 
    66.7249, 66.74606, 66.76685, 66.78726, 66.80729, 66.82694, 66.84621, 
    66.8651, 66.8836, 66.90172, 66.91945, 66.9368, 66.95377, 66.97034, 
    66.98653, 67.00232, 67.01772, 67.03274, 67.04736, 67.0616, 67.07543, 
    67.08888, 67.10193, 67.11459, 67.12685, 67.1387, 67.15017, 67.16124, 
    67.17191, 67.18217, 67.19205, 67.20152, 67.21059, 67.21925, 67.22752, 
    67.23538, 67.24284, 67.2499, 67.25656, 67.26281, 67.26866, 67.27411, 
    67.27914, 67.28378, 67.28801, 67.29184, 67.29526, 67.29827, 67.30088, 
    67.30308, 67.30488, 67.30627, 67.30725, 67.30783, 67.308, 67.30776, 
    67.30712, 67.30608, 67.30462, 67.30276, 67.30049, 67.29782, 67.29474, 
    67.29126, 67.28737, 67.28307, 67.27837, 67.27327, 67.26776, 67.26185, 
    67.25553, 67.24882, 67.24169, 67.23416, 67.22623, 67.2179, 67.20918, 
    67.20004, 67.19051, 67.18057, 67.17024, 67.15952, 67.14838, 67.13686, 
    67.12493, 67.11261, 67.09989, 67.08678, 67.07327, 67.05937, 67.04508, 
    67.0304, 67.01531, 66.99985, 66.98399, 66.96774, 66.9511, 66.93408, 
    66.91667, 66.89888, 66.8807, 66.86213, 66.84319, 66.82385, 66.80415, 
    66.78406, 66.76359, 66.74274, 66.72151, 66.69991, 66.67794, 66.65559, 
    66.63287, 66.60978, 66.58631, 66.56248, 66.53828, 66.51371, 66.48878, 
    66.46348, 66.43782, 66.4118, 66.38541, 66.35867, 66.33156, 66.3041, 
    66.27628, 66.24811, 66.21959, 66.19071, 66.16148, 66.1319, 66.10197, 
    66.0717, 66.04108, 66.01012, 65.97881, 65.94717, 65.91518, 65.88286, 
    65.85019, 65.81719, 65.78386, 65.75019, 65.71619, 65.68186, 65.6472, 
    65.61222, 65.5769, 65.54127, 65.50531, 65.46903, 65.43243, 65.39551, 
    65.35827, 65.32072, 65.28284, 65.24467, 65.20618, 65.16737, 65.12827, 
    65.08884, 65.04913, 65.00909, 64.96877, 64.92814, 64.88721, 64.84598, 
    64.80445, 64.76263, 64.72052, 64.67812, 64.63542, 64.59244, 64.54916, 
    64.50561, 64.46176, 64.41764, 64.37323, 64.32854, 64.28358, 64.23833, 
    64.19282, 64.14703, 64.10096, 64.05463, 64.00802, 63.96115, 63.91401, 
    63.8666, 63.81894, 63.771, 63.72281, 63.67436, 63.62566, 63.57669, 
    63.52747, 63.478, 63.42828, 63.3783, 63.32808, 63.27761, 63.22689, 
    63.17593, 63.12472, 63.07328, 63.02159, 62.96966, 62.9175, 62.8651, 
    62.81247, 62.7596, 62.7065, 62.65317, 62.59961, 62.54582, 62.49181, 
    62.43757, 62.38311, 62.32843, 62.27353, 62.2184, 62.16306, 62.1075, 
    62.05173, 61.99574,
  56.1111, 56.18207, 56.25292, 56.32365, 56.39427, 56.46477, 56.53515, 
    56.60541, 56.67555, 56.74557, 56.81547, 56.88525, 56.9549, 57.02443, 
    57.09383, 57.16311, 57.23225, 57.30127, 57.37017, 57.43893, 57.50756, 
    57.57606, 57.64443, 57.71267, 57.78077, 57.84873, 57.91656, 57.98426, 
    58.05181, 58.11923, 58.1865, 58.25364, 58.32064, 58.38749, 58.4542, 
    58.52076, 58.58718, 58.65345, 58.71958, 58.78555, 58.85138, 58.91706, 
    58.98258, 59.04795, 59.11317, 59.17824, 59.24314, 59.3079, 59.37249, 
    59.43693, 59.5012, 59.56532, 59.62927, 59.69306, 59.75668, 59.82014, 
    59.88344, 59.94656, 60.00952, 60.07231, 60.13493, 60.19737, 60.25965, 
    60.32174, 60.38367, 60.44541, 60.50698, 60.56837, 60.62958, 60.69061, 
    60.75145, 60.81211, 60.87259, 60.93288, 60.99298, 61.0529, 61.11263, 
    61.17216, 61.2315, 61.29065, 61.34961, 61.40836, 61.46693, 61.52529, 
    61.58345, 61.64141, 61.69917, 61.75673, 61.81408, 61.87122, 61.92816, 
    61.98489, 62.04141, 62.09772, 62.15381, 62.20969, 62.26535, 62.3208, 
    62.37603, 62.43104, 62.48583, 62.54039, 62.59474, 62.64886, 62.70275, 
    62.75641, 62.80984, 62.86305, 62.91602, 62.96876, 63.02126, 63.07353, 
    63.12556, 63.17735, 63.2289, 63.2802, 63.33127, 63.38209, 63.43266, 
    63.48299, 63.53306, 63.58289, 63.63246, 63.68178, 63.73084, 63.77965, 
    63.8282, 63.87649, 63.92452, 63.97228, 64.01978, 64.06702, 64.11399, 
    64.16069, 64.20712, 64.25329, 64.29917, 64.34478, 64.39012, 64.43518, 
    64.47996, 64.52446, 64.56867, 64.61261, 64.65626, 64.69962, 64.74269, 
    64.78548, 64.82796, 64.87016, 64.91207, 64.95368, 64.995, 65.03601, 
    65.07672, 65.11713, 65.15724, 65.19705, 65.23655, 65.27573, 65.31462, 
    65.35319, 65.39145, 65.42939, 65.46702, 65.50433, 65.54133, 65.578, 
    65.61436, 65.65038, 65.6861, 65.72147, 65.75653, 65.79125, 65.82565, 
    65.85972, 65.89345, 65.92684, 65.95991, 65.99263, 66.02502, 66.05707, 
    66.08877, 66.12013, 66.15115, 66.18182, 66.21215, 66.24213, 66.27176, 
    66.30104, 66.32996, 66.35854, 66.38676, 66.41462, 66.44212, 66.46927, 
    66.49606, 66.52248, 66.54855, 66.57425, 66.59958, 66.62455, 66.64915, 
    66.67339, 66.69725, 66.72074, 66.74387, 66.76661, 66.78899, 66.81099, 
    66.83261, 66.85385, 66.87472, 66.89521, 66.91531, 66.93504, 66.95438, 
    66.97334, 66.99192, 67.01011, 67.02791, 67.04533, 67.06236, 67.07899, 
    67.09525, 67.1111, 67.12657, 67.14165, 67.15633, 67.17062, 67.18451, 
    67.19801, 67.21111, 67.22381, 67.23611, 67.24802, 67.25954, 67.27065, 
    67.28136, 67.29167, 67.30157, 67.31109, 67.32019, 67.3289, 67.3372, 
    67.34509, 67.35258, 67.35967, 67.36636, 67.37263, 67.3785, 67.38397, 
    67.38903, 67.39368, 67.39793, 67.40177, 67.4052, 67.40823, 67.41085, 
    67.41306, 67.41486, 67.41626, 67.41724, 67.41782, 67.418, 67.41776, 
    67.41712, 67.41607, 67.4146, 67.41273, 67.41046, 67.40778, 67.40469, 
    67.40119, 67.39729, 67.39297, 67.38826, 67.38313, 67.3776, 67.37167, 
    67.36533, 67.35857, 67.35143, 67.34386, 67.33591, 67.32755, 67.31878, 
    67.30961, 67.30004, 67.29006, 67.27969, 67.26891, 67.25774, 67.24617, 
    67.2342, 67.22182, 67.20906, 67.19589, 67.18233, 67.16838, 67.15403, 
    67.13929, 67.12415, 67.10862, 67.0927, 67.07639, 67.05968, 67.0426, 
    67.02512, 67.00726, 66.98901, 66.97037, 66.95135, 66.93195, 66.91216, 
    66.89199, 66.87144, 66.85052, 66.82922, 66.80753, 66.78547, 66.76304, 
    66.74023, 66.71705, 66.6935, 66.66958, 66.64529, 66.62063, 66.5956, 
    66.57021, 66.54445, 66.51833, 66.49184, 66.465, 66.4378, 66.41024, 
    66.38232, 66.35404, 66.32542, 66.29643, 66.2671, 66.23741, 66.20738, 
    66.17699, 66.14627, 66.1152, 66.08378, 66.05202, 66.01992, 65.98748, 
    65.9547, 65.92159, 65.88813, 65.85435, 65.82023, 65.78578, 65.75101, 
    65.7159, 65.68047, 65.64471, 65.60863, 65.57222, 65.5355, 65.49845, 
    65.46109, 65.42341, 65.38541, 65.34711, 65.30849, 65.26956, 65.23032, 
    65.19077, 65.15092, 65.11076, 65.0703, 65.02954, 64.98848, 64.94712, 
    64.90546, 64.86351, 64.82127, 64.77872, 64.73589, 64.69278, 64.64937, 
    64.60567, 64.5617, 64.51743, 64.47289, 64.42807, 64.38297, 64.33759, 
    64.29193, 64.246, 64.1998, 64.15333, 64.10658, 64.05957, 64.01229, 
    63.96474, 63.91694, 63.86887, 63.82054, 63.77195, 63.7231, 63.674, 
    63.62463, 63.57502, 63.52516, 63.47504, 63.42468, 63.37407, 63.32321, 
    63.27211, 63.22076, 63.16917, 63.11734, 63.06528, 63.01297, 62.96043, 
    62.90766, 62.85465, 62.80141, 62.74794, 62.69424, 62.64031, 62.58616, 
    62.53178, 62.47718, 62.42235, 62.36731, 62.31205, 62.25656, 62.20086, 
    62.14495, 62.08882,
  56.19229, 56.26337, 56.33433, 56.40517, 56.4759, 56.54651, 56.617, 
    56.68738, 56.75763, 56.82776, 56.89777, 56.96766, 57.03743, 57.10707, 
    57.17659, 57.24598, 57.31524, 57.38438, 57.45339, 57.52227, 57.59102, 
    57.65964, 57.72813, 57.79648, 57.8647, 57.93279, 58.00074, 58.06855, 
    58.13623, 58.20376, 58.27116, 58.33842, 58.40554, 58.47251, 58.53934, 
    58.60603, 58.67257, 58.73897, 58.80522, 58.87132, 58.93727, 59.00307, 
    59.06873, 59.13422, 59.19957, 59.26476, 59.3298, 59.39468, 59.4594, 
    59.52396, 59.58837, 59.65261, 59.71669, 59.78061, 59.84437, 59.90796, 
    59.97139, 60.03465, 60.09773, 60.16065, 60.2234, 60.28598, 60.34838, 
    60.41062, 60.47268, 60.53455, 60.59626, 60.65778, 60.71912, 60.78028, 
    60.84127, 60.90207, 60.96268, 61.02311, 61.08334, 61.1434, 61.20326, 
    61.26293, 61.32241, 61.3817, 61.44079, 61.49969, 61.55838, 61.61689, 
    61.67519, 61.73329, 61.79119, 61.84888, 61.90637, 61.96366, 62.02073, 
    62.0776, 62.13426, 62.19071, 62.24694, 62.30296, 62.35877, 62.41436, 
    62.46973, 62.52488, 62.57981, 62.63451, 62.689, 62.74326, 62.79729, 
    62.8511, 62.90467, 62.95802, 63.01113, 63.06401, 63.11665, 63.16906, 
    63.22123, 63.27317, 63.32486, 63.37631, 63.42751, 63.47847, 63.52919, 
    63.57965, 63.62987, 63.67984, 63.72955, 63.77901, 63.82822, 63.87716, 
    63.92585, 63.97429, 64.02245, 64.07036, 64.118, 64.16537, 64.21249, 
    64.25933, 64.3059, 64.3522, 64.39822, 64.44397, 64.48945, 64.53465, 
    64.57956, 64.6242, 64.66855, 64.71262, 64.7564, 64.7999, 64.84311, 
    64.88603, 64.92866, 64.97099, 65.01303, 65.05477, 65.09622, 65.13737, 
    65.17822, 65.21876, 65.259, 65.29893, 65.33856, 65.37788, 65.41689, 
    65.45559, 65.49397, 65.53204, 65.5698, 65.60724, 65.64436, 65.68116, 
    65.71764, 65.75379, 65.78962, 65.82513, 65.8603, 65.89514, 65.92966, 
    65.96384, 65.9977, 66.03121, 66.06438, 66.09723, 66.12973, 66.16189, 
    66.19371, 66.22518, 66.25632, 66.28709, 66.31754, 66.34762, 66.37736, 
    66.40675, 66.43578, 66.46445, 66.49277, 66.52074, 66.54835, 66.57559, 
    66.60248, 66.62901, 66.65517, 66.68096, 66.70639, 66.73145, 66.75615, 
    66.78047, 66.80443, 66.828, 66.85122, 66.87405, 66.89651, 66.91859, 
    66.9403, 66.96162, 66.98257, 67.00314, 67.02332, 67.04313, 67.06255, 
    67.08157, 67.10023, 67.11848, 67.13636, 67.15384, 67.17094, 67.18764, 
    67.20396, 67.21988, 67.2354, 67.25053, 67.26527, 67.27962, 67.29357, 
    67.30712, 67.32027, 67.33303, 67.34538, 67.35735, 67.3689, 67.38005, 
    67.39081, 67.40116, 67.41111, 67.42065, 67.42979, 67.43854, 67.44687, 
    67.4548, 67.46232, 67.46944, 67.47614, 67.48244, 67.48834, 67.49383, 
    67.49891, 67.50359, 67.50785, 67.5117, 67.51515, 67.51819, 67.52082, 
    67.52304, 67.52485, 67.52625, 67.52724, 67.52782, 67.528, 67.52776, 
    67.52711, 67.52606, 67.52459, 67.52272, 67.52043, 67.51774, 67.51463, 
    67.51112, 67.5072, 67.50288, 67.49814, 67.49299, 67.48743, 67.48148, 
    67.47511, 67.46834, 67.46115, 67.45357, 67.44558, 67.43718, 67.42838, 
    67.41917, 67.40956, 67.39955, 67.38913, 67.37832, 67.3671, 67.35548, 
    67.34346, 67.33104, 67.31822, 67.305, 67.29139, 67.27738, 67.26297, 
    67.24817, 67.23297, 67.21738, 67.2014, 67.18503, 67.16826, 67.1511, 
    67.13356, 67.11562, 67.0973, 67.07859, 67.05949, 67.04002, 67.02016, 
    66.99991, 66.97929, 66.95827, 66.93689, 66.91512, 66.89298, 66.87046, 
    66.84757, 66.8243, 66.80066, 66.77665, 66.75227, 66.72751, 66.70239, 
    66.6769, 66.65105, 66.62483, 66.59825, 66.5713, 66.54401, 66.51634, 
    66.48832, 66.45994, 66.43121, 66.40211, 66.37268, 66.34289, 66.31274, 
    66.28225, 66.25141, 66.22023, 66.1887, 66.15682, 66.12461, 66.09206, 
    66.05916, 66.02593, 65.99236, 65.95846, 65.92422, 65.88966, 65.85476, 
    65.81953, 65.78397, 65.74809, 65.71189, 65.67536, 65.63851, 65.60134, 
    65.56385, 65.52605, 65.48792, 65.44949, 65.41074, 65.37168, 65.33231, 
    65.29263, 65.25266, 65.21236, 65.17178, 65.13088, 65.08968, 65.04819, 
    65.0064, 64.96432, 64.92194, 64.87926, 64.8363, 64.79304, 64.7495, 
    64.70567, 64.66155, 64.61716, 64.57247, 64.52751, 64.48227, 64.43675, 
    64.39096, 64.34489, 64.29855, 64.25194, 64.20506, 64.15791, 64.11048, 
    64.0628, 64.01485, 63.96664, 63.91817, 63.86944, 63.82045, 63.77121, 
    63.7217, 63.67195, 63.62194, 63.57169, 63.52118, 63.47043, 63.41943, 
    63.36818, 63.3167, 63.26497, 63.213, 63.16079, 63.10835, 63.05566, 
    63.00274, 62.9496, 62.89621, 62.8426, 62.78876, 62.73469, 62.6804, 
    62.62588, 62.57113, 62.51617, 62.46098, 62.40558, 62.34996, 62.29412, 
    62.23806, 62.18179,
  56.27334, 56.34452, 56.4156, 56.48655, 56.55739, 56.62811, 56.69872, 
    56.7692, 56.83957, 56.90981, 56.97993, 57.04994, 57.11982, 57.18958, 
    57.25921, 57.32871, 57.39809, 57.46735, 57.53647, 57.60547, 57.67434, 
    57.74307, 57.81168, 57.88015, 57.94849, 58.0167, 58.08477, 58.1527, 
    58.2205, 58.28816, 58.35568, 58.42306, 58.4903, 58.5574, 58.62435, 
    58.69116, 58.75783, 58.82435, 58.89072, 58.95695, 59.02303, 59.08895, 
    59.15473, 59.22036, 59.28583, 59.35115, 59.41631, 59.48132, 59.54617, 
    59.61087, 59.6754, 59.73977, 59.80399, 59.86804, 59.93192, 59.99564, 
    60.0592, 60.12259, 60.18581, 60.24886, 60.31175, 60.37446, 60.437, 
    60.49936, 60.56155, 60.62357, 60.6854, 60.74706, 60.80854, 60.86984, 
    60.93096, 60.99189, 61.05264, 61.1132, 61.17358, 61.23377, 61.29377, 
    61.35358, 61.4132, 61.47262, 61.53185, 61.59089, 61.64972, 61.70836, 
    61.7668, 61.82505, 61.88308, 61.94092, 61.99855, 62.05597, 62.11319, 
    62.1702, 62.227, 62.28359, 62.33996, 62.39613, 62.45207, 62.5078, 
    62.56331, 62.61861, 62.67368, 62.72853, 62.78315, 62.83755, 62.89173, 
    62.94567, 62.99939, 63.05288, 63.10614, 63.15916, 63.21194, 63.2645, 
    63.31681, 63.36889, 63.42072, 63.47231, 63.52365, 63.57476, 63.62561, 
    63.67622, 63.72658, 63.77669, 63.82655, 63.87615, 63.9255, 63.97459, 
    64.02341, 64.07199, 64.1203, 64.16834, 64.21613, 64.26365, 64.3109, 
    64.35788, 64.40459, 64.45103, 64.49719, 64.54308, 64.58869, 64.63403, 
    64.67908, 64.72385, 64.76835, 64.81255, 64.85648, 64.90011, 64.94346, 
    64.98651, 65.02927, 65.07175, 65.11392, 65.1558, 65.19737, 65.23866, 
    65.27963, 65.32031, 65.36069, 65.40075, 65.44051, 65.47996, 65.5191, 
    65.55793, 65.59644, 65.63464, 65.67252, 65.71009, 65.74734, 65.78426, 
    65.82086, 65.85714, 65.8931, 65.92872, 65.96402, 65.99899, 66.03362, 
    66.06792, 66.10189, 66.13553, 66.16882, 66.20177, 66.2344, 66.26667, 
    66.29861, 66.33019, 66.36143, 66.39233, 66.42287, 66.45307, 66.48292, 
    66.51241, 66.54155, 66.57033, 66.59875, 66.62682, 66.65453, 66.68188, 
    66.70887, 66.73549, 66.76175, 66.78764, 66.81316, 66.83833, 66.86311, 
    66.88753, 66.91158, 66.93525, 66.95854, 66.98147, 67.00401, 67.02618, 
    67.04797, 67.06937, 67.09041, 67.11105, 67.13132, 67.15119, 67.17068, 
    67.1898, 67.20851, 67.22684, 67.24479, 67.26234, 67.2795, 67.29627, 
    67.31265, 67.32864, 67.34422, 67.35942, 67.37422, 67.38862, 67.40263, 
    67.41623, 67.42944, 67.44224, 67.45464, 67.46665, 67.47826, 67.48946, 
    67.50025, 67.51064, 67.52064, 67.53022, 67.5394, 67.54817, 67.55653, 
    67.5645, 67.57205, 67.57919, 67.58593, 67.59226, 67.59818, 67.60369, 
    67.6088, 67.61349, 67.61777, 67.62164, 67.6251, 67.62815, 67.63079, 
    67.63302, 67.63484, 67.63625, 67.63724, 67.63783, 67.638, 67.63776, 
    67.63711, 67.63605, 67.63457, 67.6327, 67.6304, 67.62769, 67.62458, 
    67.62106, 67.61712, 67.61277, 67.60802, 67.60284, 67.59727, 67.59129, 
    67.58489, 67.57809, 67.57088, 67.56326, 67.55524, 67.54681, 67.53797, 
    67.52873, 67.51908, 67.50903, 67.49857, 67.48771, 67.47645, 67.46478, 
    67.45271, 67.44024, 67.42738, 67.4141, 67.40044, 67.38637, 67.3719, 
    67.35704, 67.34179, 67.32613, 67.31009, 67.29365, 67.27682, 67.25959, 
    67.24198, 67.22398, 67.20558, 67.1868, 67.16763, 67.14807, 67.12814, 
    67.10781, 67.0871, 67.06602, 67.04455, 67.0227, 67.00047, 66.97787, 
    66.95488, 66.93153, 66.9078, 66.88369, 66.85921, 66.83437, 66.80915, 
    66.78357, 66.75762, 66.7313, 66.70462, 66.67758, 66.65018, 66.62241, 
    66.59428, 66.5658, 66.53696, 66.50777, 66.47822, 66.44832, 66.41807, 
    66.38747, 66.35651, 66.32522, 66.29357, 66.26159, 66.22926, 66.19659, 
    66.16357, 66.13023, 66.09654, 66.06252, 66.02816, 65.99348, 65.95846, 
    65.9231, 65.88743, 65.85143, 65.81509, 65.77844, 65.74146, 65.70417, 
    65.66655, 65.62862, 65.59037, 65.5518, 65.51293, 65.47374, 65.43424, 
    65.39443, 65.35432, 65.3139, 65.27317, 65.23215, 65.19082, 65.14919, 
    65.10727, 65.06505, 65.02253, 64.97972, 64.93662, 64.89323, 64.84955, 
    64.80558, 64.76133, 64.7168, 64.67197, 64.62688, 64.5815, 64.53584, 
    64.48991, 64.4437, 64.39722, 64.35046, 64.30344, 64.25615, 64.20859, 
    64.16077, 64.11267, 64.06432, 64.01571, 63.96684, 63.91771, 63.86832, 
    63.81868, 63.76878, 63.71864, 63.66824, 63.61759, 63.56669, 63.51555, 
    63.46416, 63.41253, 63.36066, 63.30855, 63.2562, 63.20361, 63.15079, 
    63.09773, 63.04443, 62.99091, 62.93716, 62.88317, 62.82896, 62.77452, 
    62.71986, 62.66498, 62.60987, 62.55455, 62.499, 62.44324, 62.38726, 
    62.33106, 62.27465,
  56.35424, 56.42554, 56.49672, 56.56778, 56.63873, 56.70956, 56.78028, 
    56.85088, 56.92136, 56.99171, 57.06195, 57.13207, 57.20206, 57.27193, 
    57.34168, 57.4113, 57.4808, 57.55017, 57.61942, 57.68853, 57.75751, 
    57.82637, 57.89509, 57.96368, 58.03214, 58.10047, 58.16866, 58.23671, 
    58.30463, 58.37241, 58.44005, 58.50756, 58.57492, 58.64214, 58.70922, 
    58.77615, 58.84295, 58.90959, 58.97609, 59.04244, 59.10864, 59.1747, 
    59.2406, 59.30635, 59.37196, 59.4374, 59.50269, 59.56783, 59.63281, 
    59.69763, 59.7623, 59.8268, 59.89114, 59.95532, 60.01934, 60.08319, 
    60.14688, 60.2104, 60.27376, 60.33694, 60.39996, 60.4628, 60.52547, 
    60.58797, 60.6503, 60.71245, 60.77442, 60.83622, 60.89783, 60.95926, 
    61.02052, 61.08159, 61.14248, 61.20317, 61.26369, 61.32402, 61.38415, 
    61.4441, 61.50386, 61.56342, 61.62279, 61.68196, 61.74094, 61.79972, 
    61.8583, 61.91668, 61.97486, 62.03284, 62.09061, 62.14817, 62.20553, 
    62.26268, 62.31962, 62.37635, 62.43287, 62.48917, 62.54526, 62.60113, 
    62.65678, 62.71222, 62.76743, 62.82243, 62.87719, 62.93174, 62.98606, 
    63.04015, 63.09401, 63.14764, 63.20103, 63.2542, 63.30713, 63.35983, 
    63.41228, 63.4645, 63.51648, 63.56821, 63.6197, 63.67094, 63.72195, 
    63.7727, 63.8232, 63.87345, 63.92345, 63.97319, 64.02268, 64.07191, 
    64.12089, 64.1696, 64.21806, 64.26624, 64.31416, 64.36182, 64.40922, 
    64.45634, 64.50319, 64.54977, 64.59607, 64.64211, 64.68786, 64.73333, 
    64.77853, 64.82344, 64.86806, 64.91241, 64.95647, 65.00024, 65.04372, 
    65.08692, 65.12981, 65.17242, 65.21474, 65.25674, 65.29846, 65.33987, 
    65.38099, 65.4218, 65.4623, 65.5025, 65.54239, 65.58197, 65.62125, 
    65.6602, 65.69884, 65.73717, 65.77518, 65.81288, 65.85025, 65.88731, 
    65.92403, 65.96043, 65.99651, 66.03226, 66.06768, 66.10277, 66.13753, 
    66.17195, 66.20604, 66.23979, 66.27321, 66.30628, 66.33901, 66.37141, 
    66.40345, 66.43516, 66.46651, 66.49752, 66.52818, 66.55848, 66.58844, 
    66.61803, 66.64729, 66.67617, 66.7047, 66.73288, 66.76069, 66.78814, 
    66.81522, 66.84195, 66.86831, 66.89429, 66.91991, 66.94517, 66.97005, 
    66.99456, 67.0187, 67.04246, 67.06585, 67.08886, 67.11149, 67.13374, 
    67.15562, 67.17711, 67.19822, 67.21895, 67.23929, 67.25925, 67.27882, 
    67.298, 67.31679, 67.3352, 67.35321, 67.37083, 67.38806, 67.4049, 
    67.42134, 67.43739, 67.45304, 67.46829, 67.48315, 67.49761, 67.51167, 
    67.52533, 67.53859, 67.55145, 67.5639, 67.57595, 67.5876, 67.59885, 
    67.60969, 67.62012, 67.63016, 67.63978, 67.64899, 67.65781, 67.66621, 
    67.67419, 67.68178, 67.68896, 67.69572, 67.70207, 67.70802, 67.71355, 
    67.71867, 67.72339, 67.72768, 67.73158, 67.73505, 67.73811, 67.74076, 
    67.743, 67.74483, 67.74624, 67.74724, 67.74783, 67.748, 67.74776, 
    67.74711, 67.74604, 67.74457, 67.74268, 67.74037, 67.73766, 67.73453, 
    67.73099, 67.72704, 67.72266, 67.71789, 67.71271, 67.70711, 67.7011, 
    67.69468, 67.68785, 67.68061, 67.67296, 67.6649, 67.65644, 67.64757, 
    67.63828, 67.62859, 67.6185, 67.608, 67.5971, 67.58578, 67.57407, 
    67.56196, 67.54944, 67.53651, 67.52319, 67.50947, 67.49535, 67.48083, 
    67.4659, 67.45059, 67.43488, 67.41876, 67.40226, 67.38536, 67.36807, 
    67.35039, 67.33231, 67.31384, 67.29499, 67.27574, 67.25611, 67.23609, 
    67.21569, 67.19491, 67.17374, 67.15218, 67.13025, 67.10793, 67.08524, 
    67.06217, 67.03873, 67.01491, 66.99071, 66.96614, 66.9412, 66.91589, 
    66.89021, 66.86416, 66.83775, 66.81097, 66.78382, 66.75631, 66.72845, 
    66.70022, 66.67162, 66.64268, 66.61338, 66.58372, 66.55371, 66.52335, 
    66.49264, 66.46157, 66.43016, 66.39841, 66.3663, 66.33386, 66.30107, 
    66.26794, 66.23447, 66.20067, 66.16653, 66.13205, 66.09724, 66.0621, 
    66.02663, 65.99083, 65.9547, 65.91824, 65.88146, 65.84436, 65.80694, 
    65.7692, 65.73113, 65.69276, 65.65406, 65.61505, 65.57574, 65.5361, 
    65.49616, 65.45592, 65.41536, 65.3745, 65.33334, 65.29189, 65.25012, 
    65.20806, 65.1657, 65.12305, 65.08011, 65.03687, 64.99334, 64.94952, 
    64.90542, 64.86102, 64.81635, 64.77139, 64.72616, 64.68063, 64.63484, 
    64.58877, 64.54242, 64.4958, 64.4489, 64.40174, 64.3543, 64.3066, 
    64.25864, 64.2104, 64.16191, 64.11316, 64.06414, 64.01487, 63.96534, 
    63.91556, 63.86552, 63.81523, 63.76469, 63.71389, 63.66286, 63.61157, 
    63.56004, 63.50827, 63.45625, 63.404, 63.35151, 63.29877, 63.24581, 
    63.1926, 63.13917, 63.0855, 63.0316, 62.97748, 62.92313, 62.86855, 
    62.81374, 62.75871, 62.70346, 62.64799, 62.59231, 62.5364, 62.48028, 
    62.42394, 62.36739,
  56.435, 56.5064, 56.57769, 56.64886, 56.71993, 56.79087, 56.8617, 56.93241, 
    57.003, 57.07347, 57.14383, 57.21405, 57.28416, 57.35415, 57.42401, 
    57.49375, 57.56336, 57.63285, 57.70221, 57.77144, 57.84055, 57.90952, 
    57.97836, 58.04707, 58.11565, 58.18409, 58.2524, 58.32058, 58.38862, 
    58.45652, 58.52429, 58.59191, 58.6594, 58.72674, 58.79394, 58.861, 
    58.92792, 58.99469, 59.06131, 59.12779, 59.19412, 59.2603, 59.32633, 
    59.39221, 59.45794, 59.52351, 59.58894, 59.6542, 59.71931, 59.78426, 
    59.84906, 59.91369, 59.97816, 60.04248, 60.10662, 60.17061, 60.23443, 
    60.29808, 60.36157, 60.42489, 60.48804, 60.55102, 60.61382, 60.67646, 
    60.73892, 60.8012, 60.86331, 60.92524, 60.98699, 61.04856, 61.10995, 
    61.17116, 61.23218, 61.29302, 61.35367, 61.41413, 61.47441, 61.5345, 
    61.59439, 61.65409, 61.7136, 61.77292, 61.83204, 61.89095, 61.94968, 
    62.0082, 62.06652, 62.12463, 62.18254, 62.24025, 62.29775, 62.35504, 
    62.41212, 62.469, 62.52566, 62.5821, 62.63833, 62.69435, 62.75014, 
    62.80572, 62.86108, 62.91621, 62.97113, 63.02581, 63.08027, 63.13451, 
    63.18851, 63.24229, 63.29583, 63.34914, 63.40221, 63.45505, 63.50765, 
    63.56001, 63.61213, 63.66401, 63.71564, 63.76703, 63.81818, 63.86907, 
    63.91972, 63.97011, 64.02025, 64.07014, 64.11977, 64.16914, 64.21826, 
    64.26712, 64.31571, 64.36404, 64.41212, 64.45992, 64.50745, 64.55471, 
    64.6017, 64.64842, 64.69487, 64.74104, 64.78693, 64.83255, 64.87788, 
    64.92294, 64.9677, 65.01219, 65.05639, 65.1003, 65.14392, 65.18725, 
    65.23029, 65.27303, 65.31548, 65.35762, 65.39948, 65.44102, 65.48227, 
    65.52322, 65.56385, 65.60419, 65.64421, 65.68392, 65.72333, 65.76241, 
    65.80119, 65.83965, 65.87778, 65.91561, 65.95311, 65.99029, 66.02715, 
    66.06367, 66.09988, 66.13575, 66.1713, 66.2065, 66.24139, 66.27593, 
    66.31014, 66.34401, 66.37755, 66.41074, 66.44359, 66.4761, 66.50826, 
    66.54008, 66.57155, 66.60267, 66.63344, 66.66386, 66.69392, 66.72363, 
    66.75298, 66.78197, 66.81062, 66.83889, 66.86681, 66.89436, 66.92155, 
    66.94837, 66.97483, 67.00092, 67.02664, 67.05199, 67.07697, 67.10157, 
    67.12579, 67.14965, 67.17313, 67.19623, 67.21895, 67.24129, 67.26324, 
    67.28482, 67.30602, 67.32682, 67.34724, 67.36728, 67.38692, 67.40618, 
    67.42505, 67.44353, 67.46161, 67.4793, 67.4966, 67.5135, 67.53001, 
    67.54613, 67.56184, 67.57716, 67.59207, 67.60659, 67.6207, 67.63442, 
    67.64774, 67.66064, 67.67315, 67.68525, 67.69695, 67.70824, 67.71912, 
    67.7296, 67.73967, 67.74934, 67.75859, 67.76743, 67.77587, 67.7839, 
    67.79151, 67.79871, 67.8055, 67.81188, 67.81786, 67.82341, 67.82855, 
    67.83328, 67.8376, 67.84151, 67.84499, 67.84807, 67.85073, 67.85298, 
    67.85481, 67.85623, 67.85723, 67.85783, 67.858, 67.85776, 67.8571, 
    67.85603, 67.85455, 67.85265, 67.85034, 67.84761, 67.84447, 67.84091, 
    67.83694, 67.83257, 67.82777, 67.82256, 67.81694, 67.81091, 67.80446, 
    67.7976, 67.79033, 67.78265, 67.77456, 67.76606, 67.75715, 67.74783, 
    67.73811, 67.72797, 67.71743, 67.70648, 67.69512, 67.68336, 67.6712, 
    67.65863, 67.64565, 67.63228, 67.6185, 67.60432, 67.58974, 67.57476, 
    67.55938, 67.5436, 67.52743, 67.51086, 67.49389, 67.47653, 67.45878, 
    67.44063, 67.42209, 67.40316, 67.38384, 67.36414, 67.34404, 67.32355, 
    67.30269, 67.28143, 67.2598, 67.23778, 67.21538, 67.1926, 67.16944, 
    67.1459, 67.12199, 67.0977, 67.07304, 67.048, 67.0226, 66.99682, 
    66.97067, 66.94415, 66.91727, 66.89003, 66.86242, 66.83444, 66.80611, 
    66.77741, 66.74836, 66.71896, 66.68919, 66.65907, 66.62859, 66.59777, 
    66.56659, 66.53506, 66.5032, 66.47098, 66.43842, 66.40551, 66.37226, 
    66.33868, 66.30475, 66.27048, 66.23589, 66.20096, 66.1657, 66.1301, 
    66.09417, 66.05791, 66.02133, 65.98443, 65.9472, 65.90965, 65.87177, 
    65.83359, 65.79507, 65.75625, 65.71711, 65.67766, 65.6379, 65.59782, 
    65.55745, 65.51676, 65.47577, 65.43447, 65.39288, 65.35098, 65.30878, 
    65.26629, 65.2235, 65.18041, 65.13704, 65.09337, 65.04942, 65.00517, 
    64.96064, 64.91582, 64.87073, 64.82536, 64.77969, 64.73376, 64.68754, 
    64.64105, 64.59429, 64.54725, 64.49995, 64.45237, 64.40453, 64.35642, 
    64.30804, 64.25941, 64.21051, 64.16135, 64.11194, 64.06226, 64.01234, 
    63.96215, 63.91172, 63.86103, 63.8101, 63.75892, 63.70749, 63.65582, 
    63.6039, 63.55174, 63.49934, 63.4467, 63.39383, 63.34072, 63.28737, 
    63.2338, 63.17999, 63.12594, 63.07167, 63.01718, 62.96246, 62.90751, 
    62.85234, 62.79694, 62.74133, 62.6855, 62.62945, 62.57319, 62.51671, 
    62.46001,
  56.51561, 56.58712, 56.65852, 56.7298, 56.80098, 56.87203, 56.94297, 
    57.01379, 57.0845, 57.15508, 57.22555, 57.29589, 57.36612, 57.43622, 
    57.5062, 57.57605, 57.64578, 57.71538, 57.78486, 57.85421, 57.92343, 
    57.99252, 58.06148, 58.13031, 58.19901, 58.26758, 58.33601, 58.4043, 
    58.47247, 58.54049, 58.60838, 58.67612, 58.74373, 58.8112, 58.87853, 
    58.94571, 59.01275, 59.07965, 59.1464, 59.213, 59.27946, 59.34576, 
    59.41192, 59.47793, 59.54379, 59.60949, 59.67504, 59.74043, 59.80567, 
    59.87075, 59.93568, 60.00044, 60.06505, 60.12949, 60.19377, 60.25789, 
    60.32184, 60.38563, 60.44925, 60.5127, 60.57598, 60.6391, 60.70204, 
    60.7648, 60.8274, 60.88982, 60.95206, 61.01413, 61.07602, 61.13773, 
    61.19925, 61.2606, 61.32176, 61.38273, 61.44352, 61.50413, 61.56454, 
    61.62477, 61.6848, 61.74464, 61.80429, 61.86375, 61.923, 61.98206, 
    62.04093, 62.09959, 62.15805, 62.2163, 62.27436, 62.33221, 62.38985, 
    62.44728, 62.50451, 62.56152, 62.61833, 62.67492, 62.73129, 62.78745, 
    62.84339, 62.89911, 62.95461, 63.00989, 63.06495, 63.11977, 63.17438, 
    63.22876, 63.28291, 63.33682, 63.39051, 63.44397, 63.49718, 63.55016, 
    63.60291, 63.65541, 63.70768, 63.7597, 63.81148, 63.86301, 63.9143, 
    63.96534, 64.01614, 64.06667, 64.11696, 64.16699, 64.21677, 64.26629, 
    64.31554, 64.36455, 64.41328, 64.46176, 64.50997, 64.55791, 64.60559, 
    64.65299, 64.70013, 64.74699, 64.79358, 64.83989, 64.88593, 64.93169, 
    64.97716, 65.02235, 65.06726, 65.11189, 65.15623, 65.20027, 65.24403, 
    65.28751, 65.33068, 65.37356, 65.41615, 65.45843, 65.50041, 65.5421, 
    65.58348, 65.62457, 65.66534, 65.7058, 65.74596, 65.7858, 65.82534, 
    65.86456, 65.90347, 65.94205, 65.98032, 66.01828, 66.05591, 66.09322, 
    66.1302, 66.16685, 66.20318, 66.23918, 66.27485, 66.31019, 66.34519, 
    66.37986, 66.41419, 66.44818, 66.48183, 66.51514, 66.54812, 66.58074, 
    66.61302, 66.64495, 66.67654, 66.70777, 66.73866, 66.76919, 66.79936, 
    66.82918, 66.85864, 66.88775, 66.91649, 66.94488, 66.97289, 67.00055, 
    67.02784, 67.05477, 67.08132, 67.10751, 67.13333, 67.15878, 67.18385, 
    67.20855, 67.23287, 67.25681, 67.28038, 67.30357, 67.32638, 67.34881, 
    67.37085, 67.39251, 67.41379, 67.43468, 67.45518, 67.47529, 67.49502, 
    67.51435, 67.53329, 67.55184, 67.57, 67.58776, 67.60513, 67.6221, 
    67.63868, 67.65485, 67.67063, 67.686, 67.70098, 67.71556, 67.72974, 
    67.74351, 67.75687, 67.76983, 67.78239, 67.79454, 67.80628, 67.81762, 
    67.82855, 67.83907, 67.84918, 67.85889, 67.86818, 67.87706, 67.88553, 
    67.89359, 67.90123, 67.90847, 67.91529, 67.92169, 67.92769, 67.93327, 
    67.93843, 67.94318, 67.94752, 67.95144, 67.95494, 67.95803, 67.9607, 
    67.96296, 67.9648, 67.96622, 67.96723, 67.96783, 67.968, 67.96776, 
    67.9671, 67.96603, 67.96454, 67.96263, 67.9603, 67.95757, 67.95441, 
    67.95084, 67.94686, 67.94246, 67.93764, 67.93241, 67.92677, 67.92071, 
    67.91424, 67.90735, 67.90005, 67.89234, 67.88422, 67.87568, 67.86674, 
    67.85738, 67.84761, 67.83743, 67.82685, 67.81586, 67.80445, 67.79265, 
    67.78043, 67.76781, 67.75478, 67.74136, 67.72752, 67.71328, 67.69864, 
    67.6836, 67.66816, 67.65232, 67.63608, 67.61945, 67.60241, 67.58498, 
    67.56715, 67.54893, 67.53032, 67.51131, 67.49192, 67.47214, 67.45196, 
    67.4314, 67.41045, 67.38911, 67.36739, 67.34528, 67.3228, 67.29993, 
    67.27668, 67.25305, 67.22905, 67.20467, 67.17991, 67.15478, 67.12927, 
    67.10339, 67.07715, 67.05054, 67.02355, 66.9962, 66.96849, 66.94041, 
    66.91197, 66.88316, 66.854, 66.82449, 66.79461, 66.76438, 66.7338, 
    66.70286, 66.67156, 66.63992, 66.60794, 66.57561, 66.54292, 66.5099, 
    66.47653, 66.44283, 66.40878, 66.3744, 66.33968, 66.30462, 66.26923, 
    66.23351, 66.19746, 66.16108, 66.12437, 66.08733, 66.04998, 66.0123, 
    65.9743, 65.93597, 65.89733, 65.85838, 65.81911, 65.77953, 65.73962, 
    65.69942, 65.65891, 65.61809, 65.57696, 65.53553, 65.49379, 65.45176, 
    65.40942, 65.36679, 65.32387, 65.28065, 65.23713, 65.19333, 65.14923, 
    65.10485, 65.06018, 65.01522, 64.96999, 64.92446, 64.87866, 64.83259, 
    64.78623, 64.73959, 64.69269, 64.64552, 64.59807, 64.55035, 64.50236, 
    64.45411, 64.40559, 64.35681, 64.30777, 64.25847, 64.20891, 64.1591, 
    64.10902, 64.05869, 64.00812, 63.95729, 63.90621, 63.85488, 63.80331, 
    63.75149, 63.69943, 63.64713, 63.59458, 63.5418, 63.48878, 63.43552, 
    63.38203, 63.32831, 63.27436, 63.22017, 63.16576, 63.11111, 63.05625, 
    63.00116, 62.94584, 62.89031, 62.83455, 62.77858, 62.72239, 62.66598, 
    62.60936, 62.55252,
  56.59607, 56.66769, 56.7392, 56.8106, 56.88188, 56.95304, 57.0241, 
    57.09503, 57.16585, 57.23655, 57.30713, 57.37759, 57.44793, 57.51814, 
    57.58823, 57.6582, 57.72805, 57.79777, 57.86736, 57.93683, 58.00617, 
    58.07538, 58.14446, 58.21341, 58.28223, 58.35091, 58.41947, 58.48788, 
    58.55617, 58.62431, 58.69232, 58.76019, 58.82793, 58.89552, 58.96297, 
    59.03028, 59.09744, 59.16446, 59.23134, 59.29807, 59.36465, 59.43109, 
    59.49737, 59.56351, 59.62949, 59.69532, 59.761, 59.82653, 59.8919, 
    59.95711, 60.02216, 60.08706, 60.15179, 60.21637, 60.28078, 60.34503, 
    60.40911, 60.47304, 60.53679, 60.60038, 60.6638, 60.72704, 60.79012, 
    60.85302, 60.91575, 60.97831, 61.04069, 61.10289, 61.16491, 61.22676, 
    61.28842, 61.3499, 61.41121, 61.47232, 61.53325, 61.59399, 61.65454, 
    61.71491, 61.77508, 61.83506, 61.89486, 61.95445, 62.01385, 62.07305, 
    62.13205, 62.19086, 62.24946, 62.30786, 62.36605, 62.42405, 62.48183, 
    62.53941, 62.59678, 62.65393, 62.71088, 62.76761, 62.82413, 62.88043, 
    62.93652, 62.99238, 63.04802, 63.10345, 63.15865, 63.21362, 63.26838, 
    63.3229, 63.37719, 63.43125, 63.48508, 63.53868, 63.59205, 63.64518, 
    63.69806, 63.75071, 63.80312, 63.85529, 63.90722, 63.9589, 64.01033, 
    64.06152, 64.11245, 64.16313, 64.21356, 64.26374, 64.31366, 64.36333, 
    64.41273, 64.46188, 64.51076, 64.55938, 64.60773, 64.65582, 64.70364, 
    64.75119, 64.79847, 64.84547, 64.8922, 64.93866, 64.98483, 65.03073, 
    65.07635, 65.12169, 65.16674, 65.2115, 65.25598, 65.30017, 65.34407, 
    65.38768, 65.43099, 65.47401, 65.51673, 65.55916, 65.60128, 65.6431, 
    65.68462, 65.72584, 65.76675, 65.80735, 65.84764, 65.88762, 65.92729, 
    65.96664, 66.00568, 66.0444, 66.0828, 66.12089, 66.15865, 66.19608, 
    66.23319, 66.26997, 66.30643, 66.34256, 66.37835, 66.41382, 66.44894, 
    66.48373, 66.51819, 66.5523, 66.58607, 66.61951, 66.6526, 66.68534, 
    66.71774, 66.74979, 66.78149, 66.81284, 66.84383, 66.87447, 66.90476, 
    66.93469, 66.96426, 66.99348, 67.02233, 67.05082, 67.07895, 67.1067, 
    67.1341, 67.16113, 67.18779, 67.21407, 67.23999, 67.26553, 67.2907, 
    67.3155, 67.33991, 67.36395, 67.38761, 67.41089, 67.43378, 67.4563, 
    67.47843, 67.50018, 67.52154, 67.54251, 67.5631, 67.58328, 67.60309, 
    67.6225, 67.64152, 67.66014, 67.67838, 67.69621, 67.71365, 67.73068, 
    67.74732, 67.76357, 67.77941, 67.79485, 67.80988, 67.82452, 67.83875, 
    67.85258, 67.866, 67.87901, 67.89162, 67.90382, 67.91562, 67.927, 
    67.93797, 67.94854, 67.95869, 67.96844, 67.97776, 67.98668, 67.99519, 
    68.00328, 68.01096, 68.01822, 68.02507, 68.0315, 68.03752, 68.04312, 
    68.04831, 68.05308, 68.05743, 68.06137, 68.06489, 68.06799, 68.07067, 
    68.07294, 68.07478, 68.07622, 68.07722, 68.07782, 68.078, 68.07776, 
    68.0771, 68.07602, 68.07452, 68.07261, 68.07027, 68.06753, 68.06435, 
    68.06078, 68.05677, 68.05235, 68.04752, 68.04227, 68.0366, 68.03051, 
    68.02401, 68.0171, 68.00977, 68.00203, 67.99387, 67.9853, 67.97632, 
    67.96692, 67.95712, 67.94689, 67.93626, 67.92522, 67.91378, 67.90192, 
    67.88966, 67.87698, 67.86391, 67.85042, 67.83652, 67.82224, 67.80753, 
    67.79243, 67.77693, 67.76102, 67.74472, 67.72801, 67.71091, 67.69341, 
    67.67551, 67.65723, 67.63853, 67.61945, 67.59998, 67.58012, 67.55986, 
    67.53922, 67.51819, 67.49677, 67.47496, 67.45277, 67.43019, 67.40723, 
    67.3839, 67.36018, 67.33607, 67.3116, 67.28675, 67.26152, 67.23592, 
    67.20995, 67.18359, 67.15688, 67.12979, 67.10234, 67.07452, 67.04634, 
    67.01779, 66.98888, 66.95961, 66.92999, 66.89999, 66.86965, 66.83895, 
    66.8079, 66.7765, 66.74474, 66.71264, 66.68018, 66.64738, 66.61424, 
    66.58076, 66.54693, 66.51276, 66.47825, 66.44341, 66.40823, 66.37271, 
    66.33687, 66.30069, 66.26418, 66.22734, 66.19019, 66.15269, 66.11488, 
    66.07675, 66.0383, 65.99953, 65.96044, 65.92104, 65.88132, 65.84129, 
    65.80095, 65.7603, 65.71934, 65.67808, 65.63651, 65.59464, 65.55247, 
    65.50999, 65.46722, 65.42416, 65.3808, 65.33714, 65.2932, 65.24896, 
    65.20444, 65.15963, 65.11453, 65.06915, 65.02349, 64.97755, 64.93133, 
    64.88483, 64.83805, 64.79101, 64.74368, 64.69609, 64.64823, 64.6001, 
    64.5517, 64.50304, 64.45412, 64.40493, 64.35548, 64.30579, 64.25582, 
    64.2056, 64.15514, 64.10441, 64.05344, 64.00221, 63.95074, 63.89902, 
    63.84706, 63.79485, 63.7424, 63.68971, 63.63679, 63.58362, 63.53022, 
    63.47659, 63.42272, 63.36862, 63.31429, 63.25973, 63.20494, 63.14993, 
    63.0947, 63.03924, 62.98356, 62.92766, 62.87154, 62.8152, 62.75865, 
    62.70189, 62.64491,
  56.67638, 56.74811, 56.81973, 56.89124, 56.96263, 57.03391, 57.10508, 
    57.17612, 57.24705, 57.31786, 57.38856, 57.45913, 57.52958, 57.59991, 
    57.67012, 57.74021, 57.81017, 57.88001, 57.94972, 58.01931, 58.08876, 
    58.15809, 58.22729, 58.29636, 58.3653, 58.4341, 58.50278, 58.57132, 
    58.63972, 58.70799, 58.77612, 58.84412, 58.91197, 58.97969, 59.04726, 
    59.1147, 59.18199, 59.24913, 59.31614, 59.38299, 59.4497, 59.51627, 
    59.58268, 59.64894, 59.71505, 59.78102, 59.84682, 59.91248, 59.97798, 
    60.04332, 60.10851, 60.17353, 60.2384, 60.3031, 60.36765, 60.43203, 
    60.49625, 60.56031, 60.6242, 60.68792, 60.75146, 60.81485, 60.87806, 
    60.9411, 61.00397, 61.06666, 61.12917, 61.19151, 61.25368, 61.31566, 
    61.37746, 61.43908, 61.50052, 61.56177, 61.62284, 61.68372, 61.74442, 
    61.80492, 61.86524, 61.92536, 61.98529, 62.04502, 62.10456, 62.16391, 
    62.22305, 62.282, 62.34074, 62.39929, 62.45763, 62.51576, 62.57369, 
    62.63141, 62.68892, 62.74622, 62.80331, 62.86019, 62.91685, 62.9733, 
    63.02953, 63.08553, 63.14132, 63.19689, 63.25224, 63.30736, 63.36226, 
    63.41692, 63.47136, 63.52557, 63.57955, 63.63329, 63.6868, 63.74007, 
    63.79311, 63.84591, 63.89846, 63.95078, 64.00285, 64.05467, 64.10625, 
    64.15759, 64.20866, 64.25949, 64.31007, 64.36039, 64.41046, 64.46027, 
    64.50982, 64.55911, 64.60814, 64.6569, 64.7054, 64.75363, 64.8016, 
    64.84929, 64.89671, 64.94386, 64.99074, 65.03734, 65.08366, 65.1297, 
    65.17546, 65.22093, 65.26613, 65.31104, 65.35565, 65.39999, 65.44402, 
    65.48778, 65.53123, 65.57439, 65.61725, 65.65981, 65.70207, 65.74403, 
    65.78569, 65.82704, 65.86809, 65.90883, 65.94926, 65.98937, 66.02917, 
    66.06866, 66.10783, 66.14668, 66.18522, 66.22343, 66.26132, 66.29889, 
    66.33613, 66.37304, 66.40962, 66.44588, 66.4818, 66.51739, 66.55264, 
    66.58755, 66.62213, 66.65637, 66.69027, 66.72382, 66.75703, 66.78989, 
    66.82241, 66.85458, 66.88639, 66.91785, 66.94897, 66.97972, 67.01012, 
    67.04016, 67.06985, 67.09917, 67.12813, 67.15673, 67.18496, 67.21283, 
    67.24033, 67.26746, 67.29422, 67.32061, 67.34663, 67.37227, 67.39753, 
    67.42242, 67.44693, 67.47106, 67.49482, 67.51819, 67.54118, 67.56377, 
    67.58599, 67.60783, 67.62927, 67.65032, 67.67099, 67.69126, 67.71114, 
    67.73064, 67.74973, 67.76842, 67.78673, 67.80463, 67.82214, 67.83926, 
    67.85596, 67.87227, 67.88818, 67.90368, 67.91878, 67.93347, 67.94776, 
    67.96165, 67.97512, 67.98819, 68.00085, 68.0131, 68.02494, 68.03637, 
    68.04739, 68.058, 68.06819, 68.07798, 68.08735, 68.0963, 68.10484, 
    68.11297, 68.12067, 68.12797, 68.13485, 68.1413, 68.14735, 68.15298, 
    68.15819, 68.16297, 68.16734, 68.1713, 68.17483, 68.17795, 68.18064, 
    68.18291, 68.18477, 68.18621, 68.18723, 68.18782, 68.188, 68.18775, 
    68.1871, 68.18601, 68.18451, 68.18259, 68.18024, 68.17748, 68.1743, 
    68.1707, 68.16668, 68.16225, 68.15739, 68.15211, 68.14642, 68.14031, 
    68.13379, 68.12685, 68.11948, 68.11171, 68.10352, 68.09491, 68.08589, 
    68.07645, 68.06661, 68.05635, 68.04568, 68.03459, 68.02309, 68.01119, 
    67.99887, 67.98615, 67.97301, 67.95947, 67.94553, 67.93118, 67.91641, 
    67.90125, 67.88569, 67.86972, 67.85335, 67.83657, 67.8194, 67.80183, 
    67.78386, 67.7655, 67.74673, 67.72758, 67.70802, 67.68808, 67.66775, 
    67.64702, 67.6259, 67.6044, 67.5825, 67.56023, 67.53756, 67.51452, 
    67.49108, 67.46727, 67.44308, 67.41851, 67.39356, 67.36823, 67.34253, 
    67.31646, 67.29001, 67.26319, 67.236, 67.20844, 67.18052, 67.15223, 
    67.12357, 67.09456, 67.06518, 67.03544, 67.00534, 66.97488, 66.94407, 
    66.9129, 66.88138, 66.84951, 66.81728, 66.78471, 66.7518, 66.71854, 
    66.68493, 66.65098, 66.61668, 66.58205, 66.54709, 66.51178, 66.47614, 
    66.44016, 66.40386, 66.36723, 66.33026, 66.29297, 66.25535, 66.21741, 
    66.17915, 66.14056, 66.10165, 66.06243, 66.0229, 65.98305, 65.94288, 
    65.9024, 65.86162, 65.82053, 65.77912, 65.73742, 65.69541, 65.6531, 
    65.61049, 65.56758, 65.52438, 65.48087, 65.43708, 65.39299, 65.34862, 
    65.30395, 65.259, 65.21376, 65.16824, 65.12244, 65.07635, 65.02998, 
    64.98334, 64.93642, 64.88923, 64.84177, 64.79403, 64.74602, 64.69775, 
    64.64921, 64.6004, 64.55133, 64.502, 64.45241, 64.40256, 64.35245, 
    64.30209, 64.25147, 64.2006, 64.14948, 64.09811, 64.04649, 63.99463, 
    63.94252, 63.89017, 63.83757, 63.78474, 63.73166, 63.67835, 63.62481, 
    63.57103, 63.51701, 63.46276, 63.40829, 63.35359, 63.29866, 63.2435, 
    63.18812, 63.13251, 63.07669, 63.02065, 62.96438, 62.9079, 62.8512, 
    62.7943, 62.73717,
  56.75654, 56.82838, 56.90011, 56.97173, 57.04324, 57.11463, 57.1859, 
    57.25706, 57.32811, 57.39903, 57.46984, 57.54052, 57.61109, 57.68154, 
    57.75187, 57.82207, 57.89215, 57.9621, 58.03193, 58.10163, 58.17121, 
    58.24066, 58.30997, 58.37917, 58.44822, 58.51715, 58.58595, 58.65461, 
    58.72313, 58.79152, 58.85978, 58.92789, 58.99588, 59.06371, 59.13141, 
    59.19897, 59.26639, 59.33366, 59.40079, 59.46777, 59.53461, 59.6013, 
    59.66784, 59.73423, 59.80048, 59.86657, 59.9325, 59.99829, 60.06392, 
    60.12939, 60.19471, 60.25986, 60.32486, 60.38971, 60.45438, 60.5189, 
    60.58325, 60.64744, 60.71146, 60.77531, 60.839, 60.90252, 60.96587, 
    61.02904, 61.09204, 61.15487, 61.21753, 61.28, 61.3423, 61.40442, 
    61.46637, 61.52813, 61.5897, 61.65109, 61.7123, 61.77332, 61.83416, 
    61.89481, 61.95526, 62.01552, 62.0756, 62.13547, 62.19516, 62.25464, 
    62.31393, 62.37302, 62.4319, 62.49059, 62.54907, 62.60735, 62.66542, 
    62.72329, 62.78094, 62.83839, 62.89562, 62.95264, 63.00945, 63.06604, 
    63.12241, 63.17857, 63.2345, 63.29022, 63.34571, 63.40098, 63.45602, 
    63.51083, 63.56542, 63.61977, 63.6739, 63.72779, 63.78144, 63.83487, 
    63.88805, 63.94099, 63.99369, 64.04616, 64.09837, 64.15034, 64.20207, 
    64.25355, 64.30477, 64.35575, 64.40647, 64.45695, 64.50716, 64.55711, 
    64.60681, 64.65624, 64.70542, 64.75433, 64.80297, 64.85135, 64.89946, 
    64.9473, 64.99487, 65.04216, 65.08918, 65.13593, 65.18239, 65.22858, 
    65.27448, 65.3201, 65.36543, 65.41048, 65.45525, 65.49972, 65.5439, 
    65.58779, 65.63139, 65.67468, 65.71769, 65.76039, 65.8028, 65.84489, 
    65.88669, 65.92818, 65.96936, 66.01023, 66.0508, 66.09105, 66.13099, 
    66.17061, 66.20992, 66.2489, 66.28757, 66.32591, 66.36394, 66.40163, 
    66.439, 66.47604, 66.51276, 66.54914, 66.58519, 66.6209, 66.65628, 
    66.69132, 66.72603, 66.76038, 66.7944, 66.82808, 66.86141, 66.89439, 
    66.92703, 66.95931, 66.99125, 67.02283, 67.05405, 67.08493, 67.11544, 
    67.1456, 67.17539, 67.20483, 67.23389, 67.2626, 67.29094, 67.31892, 
    67.34652, 67.37376, 67.40062, 67.42711, 67.45322, 67.47897, 67.50433, 
    67.52932, 67.55392, 67.57815, 67.602, 67.62546, 67.64854, 67.67123, 
    67.69353, 67.71545, 67.73698, 67.75812, 67.77887, 67.79922, 67.81918, 
    67.83875, 67.85793, 67.87669, 67.89507, 67.91306, 67.93063, 67.94781, 
    67.96458, 67.98096, 67.99693, 68.0125, 68.02766, 68.04241, 68.05676, 
    68.0707, 68.08424, 68.09736, 68.11007, 68.12237, 68.13426, 68.14574, 
    68.15681, 68.16746, 68.1777, 68.18752, 68.19692, 68.20592, 68.21449, 
    68.22265, 68.23039, 68.23772, 68.24462, 68.25111, 68.25718, 68.26283, 
    68.26806, 68.27287, 68.27726, 68.28123, 68.28477, 68.2879, 68.29061, 
    68.29289, 68.29476, 68.2962, 68.29722, 68.29782, 68.298, 68.29775, 
    68.29709, 68.296, 68.29449, 68.29256, 68.29021, 68.28744, 68.28424, 
    68.28062, 68.27659, 68.27213, 68.26726, 68.26196, 68.25625, 68.25011, 
    68.24356, 68.23659, 68.22919, 68.22139, 68.21317, 68.20452, 68.19547, 
    68.18599, 68.1761, 68.16579, 68.15508, 68.14395, 68.13241, 68.12045, 
    68.10809, 68.09531, 68.08212, 68.06852, 68.05452, 68.04011, 68.02528, 
    68.01006, 67.99443, 67.97839, 67.96196, 67.94512, 67.92788, 67.91023, 
    67.8922, 67.87376, 67.85492, 67.83568, 67.81606, 67.79603, 67.77561, 
    67.7548, 67.7336, 67.71201, 67.69003, 67.66766, 67.64491, 67.62177, 
    67.59825, 67.57434, 67.55006, 67.52539, 67.50034, 67.47492, 67.44912, 
    67.42294, 67.39639, 67.36947, 67.34218, 67.31451, 67.28648, 67.25809, 
    67.22932, 67.2002, 67.1707, 67.14085, 67.11064, 67.08007, 67.04914, 
    67.01786, 66.98622, 66.95423, 66.92189, 66.8892, 66.85616, 66.82278, 
    66.78905, 66.75497, 66.72056, 66.68581, 66.65071, 66.61528, 66.57951, 
    66.54341, 66.50697, 66.47021, 66.43311, 66.39569, 66.35794, 66.31987, 
    66.28147, 66.24276, 66.20372, 66.16436, 66.12469, 66.0847, 66.0444, 
    66.00379, 65.96287, 65.92163, 65.8801, 65.83825, 65.7961, 65.75365, 
    65.71091, 65.66785, 65.62451, 65.58087, 65.53693, 65.49271, 65.44819, 
    65.40337, 65.35828, 65.3129, 65.26723, 65.22128, 65.17506, 65.12855, 
    65.08176, 65.0347, 64.98736, 64.93975, 64.89187, 64.84372, 64.7953, 
    64.74661, 64.69765, 64.64845, 64.59897, 64.54922, 64.49923, 64.44897, 
    64.39847, 64.3477, 64.29669, 64.24542, 64.1939, 64.14214, 64.09013, 
    64.03787, 63.98537, 63.93263, 63.87965, 63.82643, 63.77298, 63.71928, 
    63.66535, 63.61119, 63.5568, 63.50218, 63.44733, 63.39225, 63.33695, 
    63.28142, 63.22567, 63.1697, 63.11351, 63.0571, 63.00048, 62.94364, 
    62.88658, 62.82932,
  56.83655, 56.9085, 56.98034, 57.05207, 57.12369, 57.19519, 57.26658, 
    57.33785, 57.40901, 57.48005, 57.55097, 57.62177, 57.69245, 57.76302, 
    57.83345, 57.90377, 57.97397, 58.04404, 58.11399, 58.18381, 58.25351, 
    58.32307, 58.39251, 58.46182, 58.531, 58.60005, 58.66896, 58.73774, 
    58.80639, 58.87491, 58.94328, 59.01152, 59.07963, 59.14759, 59.21542, 
    59.2831, 59.35064, 59.41804, 59.4853, 59.55241, 59.61937, 59.68619, 
    59.75286, 59.81938, 59.88575, 59.95197, 60.01804, 60.08395, 60.14971, 
    60.21532, 60.28077, 60.34605, 60.41119, 60.47616, 60.54097, 60.60562, 
    60.6701, 60.73443, 60.79858, 60.86258, 60.9264, 60.99005, 61.05354, 
    61.11684, 61.17999, 61.24295, 61.30574, 61.36836, 61.43079, 61.49305, 
    61.55513, 61.61703, 61.67875, 61.74028, 61.80163, 61.86279, 61.92377, 
    61.98455, 62.04515, 62.10556, 62.16577, 62.22579, 62.28561, 62.34524, 
    62.40467, 62.46391, 62.52293, 62.58176, 62.64039, 62.69881, 62.75703, 
    62.81504, 62.87284, 62.93043, 62.98781, 63.04498, 63.10193, 63.15866, 
    63.21519, 63.27149, 63.32757, 63.38343, 63.43907, 63.49448, 63.54967, 
    63.60463, 63.65936, 63.71387, 63.76814, 63.82217, 63.87598, 63.92955, 
    63.98288, 64.03596, 64.08881, 64.14143, 64.19379, 64.24591, 64.29778, 
    64.34941, 64.40078, 64.4519, 64.50278, 64.55339, 64.60375, 64.65385, 
    64.7037, 64.75328, 64.8026, 64.85166, 64.90045, 64.94897, 64.99723, 
    65.04522, 65.09293, 65.14037, 65.18754, 65.23442, 65.28103, 65.32736, 
    65.37341, 65.41917, 65.46465, 65.50985, 65.55476, 65.59937, 65.64369, 
    65.68773, 65.73146, 65.7749, 65.81805, 65.86089, 65.90343, 65.94567, 
    65.98761, 66.02924, 66.07056, 66.11157, 66.15227, 66.19266, 66.23273, 
    66.27249, 66.31194, 66.35105, 66.38985, 66.42834, 66.46649, 66.50432, 
    66.54182, 66.57899, 66.61584, 66.65234, 66.68852, 66.72437, 66.75987, 
    66.79504, 66.82986, 66.86435, 66.89849, 66.93229, 66.96574, 66.99885, 
    67.03161, 67.06401, 67.09606, 67.12776, 67.1591, 67.19009, 67.22072, 
    67.25098, 67.2809, 67.31044, 67.33962, 67.36844, 67.39689, 67.42496, 
    67.45267, 67.48002, 67.50698, 67.53358, 67.55979, 67.58563, 67.6111, 
    67.63618, 67.66089, 67.68521, 67.70914, 67.7327, 67.75587, 67.77866, 
    67.80105, 67.82305, 67.84467, 67.86589, 67.88673, 67.90716, 67.9272, 
    67.94685, 67.9661, 67.98495, 68.0034, 68.02145, 68.0391, 68.05635, 
    68.0732, 68.08964, 68.10567, 68.12131, 68.13653, 68.15134, 68.16575, 
    68.17975, 68.19334, 68.20651, 68.21928, 68.23163, 68.24357, 68.2551, 
    68.26621, 68.27691, 68.28719, 68.29705, 68.3065, 68.31553, 68.32414, 
    68.33234, 68.34011, 68.34747, 68.3544, 68.36092, 68.367, 68.37268, 
    68.37793, 68.38276, 68.38717, 68.39116, 68.39472, 68.39786, 68.40058, 
    68.40287, 68.40475, 68.4062, 68.40722, 68.40782, 68.408, 68.40775, 
    68.40708, 68.40599, 68.40448, 68.40254, 68.40018, 68.39739, 68.39419, 
    68.39056, 68.3865, 68.38203, 68.37713, 68.37181, 68.36607, 68.35991, 
    68.35333, 68.34633, 68.33891, 68.33106, 68.32281, 68.31413, 68.30503, 
    68.29552, 68.28559, 68.27524, 68.26448, 68.2533, 68.24171, 68.22971, 
    68.21729, 68.20446, 68.19122, 68.17756, 68.1635, 68.14902, 68.13415, 
    68.11886, 68.10316, 68.08707, 68.07056, 68.05365, 68.03634, 68.01862, 
    68.00051, 67.98199, 67.96308, 67.94377, 67.92406, 67.90395, 67.88345, 
    67.86256, 67.84128, 67.8196, 67.79753, 67.77508, 67.75224, 67.729, 
    67.70539, 67.68139, 67.65701, 67.63224, 67.60709, 67.58157, 67.55567, 
    67.5294, 67.50274, 67.47572, 67.44832, 67.42055, 67.39241, 67.36391, 
    67.33503, 67.30579, 67.27619, 67.24622, 67.2159, 67.18521, 67.15417, 
    67.12277, 67.09102, 67.05891, 67.02644, 66.99364, 66.96048, 66.92697, 
    66.89312, 66.85892, 66.82438, 66.7895, 66.75428, 66.71872, 66.68282, 
    66.64659, 66.61003, 66.57314, 66.53591, 66.49835, 66.46047, 66.42227, 
    66.38374, 66.34489, 66.30572, 66.26622, 66.22642, 66.18629, 66.14585, 
    66.1051, 66.06404, 66.02267, 65.981, 65.93901, 65.89672, 65.85413, 
    65.81124, 65.76805, 65.72456, 65.68078, 65.6367, 65.59233, 65.54767, 
    65.50272, 65.45748, 65.41196, 65.36614, 65.32005, 65.27368, 65.22703, 
    65.18009, 65.13288, 65.0854, 65.03764, 64.98962, 64.94131, 64.89275, 
    64.84392, 64.79482, 64.74546, 64.69583, 64.64595, 64.5958, 64.5454, 
    64.49474, 64.44383, 64.39267, 64.34126, 64.2896, 64.23768, 64.18552, 
    64.13312, 64.08047, 64.02759, 63.97446, 63.92109, 63.86749, 63.81364, 
    63.75957, 63.70526, 63.65072, 63.59595, 63.54095, 63.48573, 63.43028, 
    63.37461, 63.31871, 63.2626, 63.20626, 63.14971, 63.09293, 63.03595, 
    62.97875, 62.92133,
  56.9164, 56.98847, 57.06042, 57.13226, 57.20399, 57.2756, 57.3471, 
    57.41849, 57.48976, 57.56091, 57.63195, 57.70286, 57.77366, 57.84434, 
    57.91489, 57.98533, 58.05564, 58.12583, 58.1959, 58.26583, 58.33565, 
    58.40533, 58.4749, 58.54432, 58.61362, 58.68279, 58.75183, 58.82073, 
    58.8895, 58.95814, 59.02664, 59.09501, 59.16323, 59.23132, 59.29927, 
    59.36708, 59.43475, 59.50227, 59.56966, 59.63689, 59.70399, 59.77093, 
    59.83773, 59.90438, 59.97088, 60.03723, 60.10343, 60.16947, 60.23536, 
    60.3011, 60.36668, 60.4321, 60.49737, 60.56247, 60.62742, 60.6922, 
    60.75682, 60.82128, 60.88557, 60.9497, 61.01365, 61.07744, 61.14106, 
    61.20451, 61.26779, 61.33089, 61.39382, 61.45657, 61.51915, 61.58155, 
    61.64377, 61.70581, 61.76766, 61.82933, 61.89082, 61.95213, 62.01324, 
    62.07417, 62.13491, 62.19546, 62.25581, 62.31598, 62.37594, 62.43571, 
    62.49529, 62.55466, 62.61384, 62.67281, 62.73159, 62.79015, 62.84851, 
    62.90667, 62.96461, 63.02235, 63.07988, 63.13719, 63.19429, 63.25117, 
    63.30784, 63.36428, 63.42051, 63.47652, 63.53231, 63.58787, 63.6432, 
    63.69831, 63.75319, 63.80784, 63.86226, 63.91645, 63.9704, 64.02412, 
    64.07759, 64.13083, 64.18383, 64.23659, 64.2891, 64.34137, 64.39339, 
    64.44516, 64.49668, 64.54796, 64.59898, 64.64974, 64.70025, 64.7505, 
    64.80049, 64.85022, 64.89969, 64.94889, 64.99783, 65.0465, 65.09491, 
    65.14304, 65.1909, 65.23849, 65.2858, 65.33283, 65.37959, 65.42606, 
    65.47225, 65.51817, 65.56379, 65.60913, 65.65417, 65.69894, 65.74341, 
    65.78758, 65.83146, 65.87505, 65.91833, 65.96131, 66.004, 66.04638, 
    66.08846, 66.13022, 66.17168, 66.21283, 66.25367, 66.2942, 66.33441, 
    66.37431, 66.41388, 66.45314, 66.49207, 66.53069, 66.56898, 66.60694, 
    66.64457, 66.68188, 66.71885, 66.75549, 66.7918, 66.82777, 66.8634, 
    66.8987, 66.93365, 66.96826, 67.00253, 67.03645, 67.07003, 67.10326, 
    67.13613, 67.16866, 67.20083, 67.23264, 67.26411, 67.29521, 67.32595, 
    67.35634, 67.38636, 67.41602, 67.4453, 67.47424, 67.50279, 67.53098, 
    67.5588, 67.58624, 67.61331, 67.64001, 67.66633, 67.69228, 67.71783, 
    67.74302, 67.76782, 67.79224, 67.81628, 67.83992, 67.86318, 67.88605, 
    67.90854, 67.93063, 67.95234, 67.97365, 67.99456, 68.01508, 68.0352, 
    68.05493, 68.07426, 68.09319, 68.11171, 68.12984, 68.14756, 68.16488, 
    68.18179, 68.1983, 68.21441, 68.2301, 68.24538, 68.26026, 68.27473, 
    68.28879, 68.30243, 68.31567, 68.32848, 68.34089, 68.35287, 68.36445, 
    68.37561, 68.38635, 68.39668, 68.40658, 68.41607, 68.42513, 68.43378, 
    68.44201, 68.44982, 68.45721, 68.46417, 68.47071, 68.47683, 68.48253, 
    68.4878, 68.49265, 68.49708, 68.50108, 68.50466, 68.50782, 68.51054, 
    68.51285, 68.51473, 68.51619, 68.51721, 68.51782, 68.518, 68.51775, 
    68.51708, 68.51598, 68.51447, 68.51251, 68.51015, 68.50735, 68.50413, 
    68.50048, 68.49641, 68.49191, 68.487, 68.48166, 68.47589, 68.4697, 
    68.4631, 68.45606, 68.44862, 68.44073, 68.43244, 68.42373, 68.4146, 
    68.40504, 68.39507, 68.38468, 68.37387, 68.36265, 68.35101, 68.33895, 
    68.32648, 68.3136, 68.3003, 68.28659, 68.27247, 68.25794, 68.243, 
    68.22765, 68.21188, 68.19572, 68.17915, 68.16217, 68.14478, 68.127, 
    68.10881, 68.09022, 68.07123, 68.05183, 68.03205, 68.01186, 67.99128, 
    67.9703, 67.94893, 67.92717, 67.90501, 67.88247, 67.85953, 67.8362, 
    67.8125, 67.78841, 67.76392, 67.73906, 67.71382, 67.68819, 67.66219, 
    67.63581, 67.60905, 67.58192, 67.55442, 67.52654, 67.4983, 67.46968, 
    67.4407, 67.41135, 67.38164, 67.35155, 67.32111, 67.29031, 67.25916, 
    67.22764, 67.19576, 67.16354, 67.13096, 67.09802, 67.06474, 67.03111, 
    66.99713, 66.96281, 66.92815, 66.89314, 66.85779, 66.82211, 66.78608, 
    66.74972, 66.71303, 66.676, 66.63864, 66.60095, 66.56294, 66.5246, 
    66.48594, 66.44695, 66.40765, 66.36801, 66.32807, 66.28781, 66.24723, 
    66.20634, 66.16515, 66.12363, 66.08182, 66.0397, 65.99727, 65.95454, 
    65.9115, 65.86817, 65.82454, 65.78061, 65.73639, 65.69188, 65.64707, 
    65.60197, 65.55659, 65.51093, 65.46497, 65.41873, 65.37221, 65.32541, 
    65.27833, 65.23097, 65.18335, 65.13544, 65.08727, 65.03883, 64.99011, 
    64.94113, 64.89188, 64.84237, 64.7926, 64.74257, 64.69228, 64.64172, 
    64.59092, 64.53986, 64.48855, 64.43699, 64.38518, 64.33311, 64.28081, 
    64.22826, 64.17546, 64.12243, 64.06915, 64.01563, 63.96188, 63.90789, 
    63.85367, 63.79921, 63.74453, 63.68961, 63.63446, 63.57909, 63.5235, 
    63.46768, 63.41163, 63.35537, 63.29889, 63.24219, 63.18527, 63.12814, 
    63.07079, 63.01323,
  56.99611, 57.06828, 57.14034, 57.2123, 57.28413, 57.35586, 57.42747, 
    57.49897, 57.57035, 57.64162, 57.71277, 57.7838, 57.85471, 57.92551, 
    57.99618, 58.06673, 58.13716, 58.20747, 58.27765, 58.34771, 58.41764, 
    58.48745, 58.55713, 58.62667, 58.6961, 58.76539, 58.83455, 58.90357, 
    58.97247, 59.04123, 59.10985, 59.17834, 59.24669, 59.3149, 59.38298, 
    59.45091, 59.51871, 59.58636, 59.65387, 59.72123, 59.78845, 59.85553, 
    59.92245, 59.98923, 60.05586, 60.12234, 60.18867, 60.25485, 60.32087, 
    60.38674, 60.45245, 60.51801, 60.5834, 60.64864, 60.71372, 60.77864, 
    60.84339, 60.90799, 60.97241, 61.03667, 61.10077, 61.16469, 61.22845, 
    61.29203, 61.35545, 61.41869, 61.48176, 61.54465, 61.60736, 61.6699, 
    61.73226, 61.79444, 61.85644, 61.91825, 61.97988, 62.04132, 62.10258, 
    62.16365, 62.22454, 62.28522, 62.34573, 62.40603, 62.46614, 62.52606, 
    62.58577, 62.64529, 62.70461, 62.76373, 62.82265, 62.88136, 62.93987, 
    62.99817, 63.05626, 63.11414, 63.17181, 63.22927, 63.28652, 63.34355, 
    63.40036, 63.45696, 63.51334, 63.56949, 63.62542, 63.68113, 63.73662, 
    63.79187, 63.8469, 63.9017, 63.95627, 64.0106, 64.0647, 64.11857, 
    64.1722, 64.22559, 64.27873, 64.33163, 64.3843, 64.43671, 64.48888, 
    64.54081, 64.59248, 64.6439, 64.69507, 64.74598, 64.79664, 64.84704, 
    64.89718, 64.94706, 64.99667, 65.04603, 65.09512, 65.14394, 65.19248, 
    65.24076, 65.28877, 65.33651, 65.38396, 65.43114, 65.47805, 65.52467, 
    65.57101, 65.61707, 65.66283, 65.70832, 65.75352, 65.79842, 65.84303, 
    65.88735, 65.93137, 65.97511, 66.01853, 66.06166, 66.10448, 66.147, 
    66.18922, 66.23113, 66.27273, 66.31403, 66.355, 66.39567, 66.43601, 
    66.47605, 66.51576, 66.55515, 66.59423, 66.63298, 66.6714, 66.7095, 
    66.74726, 66.7847, 66.82181, 66.85858, 66.89502, 66.93111, 66.96688, 
    67.0023, 67.03738, 67.07212, 67.10651, 67.14056, 67.17426, 67.20761, 
    67.24061, 67.27325, 67.30555, 67.33749, 67.36906, 67.40028, 67.43114, 
    67.46165, 67.49178, 67.52155, 67.55096, 67.57999, 67.60866, 67.63696, 
    67.66489, 67.69244, 67.71961, 67.74641, 67.77283, 67.79888, 67.82455, 
    67.84983, 67.87473, 67.89925, 67.92338, 67.94712, 67.97047, 67.99344, 
    68.01601, 68.03819, 68.05998, 68.08138, 68.10238, 68.12298, 68.14319, 
    68.16299, 68.1824, 68.20141, 68.22001, 68.2382, 68.256, 68.27339, 
    68.29038, 68.30695, 68.32313, 68.33888, 68.35423, 68.36918, 68.38371, 
    68.39782, 68.41152, 68.4248, 68.43768, 68.45013, 68.46217, 68.4738, 
    68.485, 68.49579, 68.50616, 68.51611, 68.52563, 68.53474, 68.54343, 
    68.55169, 68.55953, 68.56695, 68.57394, 68.58051, 68.58665, 68.59238, 
    68.59767, 68.60255, 68.60699, 68.61102, 68.61461, 68.61777, 68.62051, 
    68.62283, 68.62472, 68.62617, 68.62721, 68.62782, 68.628, 68.62775, 
    68.62708, 68.62598, 68.62445, 68.62249, 68.62011, 68.6173, 68.61407, 
    68.6104, 68.60632, 68.60181, 68.59686, 68.5915, 68.58572, 68.5795, 
    68.57286, 68.5658, 68.55832, 68.55041, 68.54208, 68.53333, 68.52415, 
    68.51456, 68.50455, 68.49411, 68.48326, 68.47198, 68.4603, 68.4482, 
    68.43567, 68.42273, 68.40938, 68.39561, 68.38143, 68.36684, 68.35184, 
    68.33642, 68.32059, 68.30436, 68.28772, 68.27067, 68.25322, 68.23536, 
    68.21709, 68.19843, 68.17936, 68.15989, 68.14001, 68.11975, 68.09908, 
    68.07802, 68.05656, 68.03471, 68.01247, 67.98983, 67.9668, 67.94339, 
    67.91959, 67.89539, 67.87082, 67.84586, 67.82051, 67.79479, 67.76868, 
    67.7422, 67.71534, 67.6881, 67.66049, 67.63251, 67.60415, 67.57542, 
    67.54633, 67.51687, 67.48704, 67.45685, 67.42628, 67.39537, 67.36409, 
    67.33246, 67.30046, 67.26811, 67.23541, 67.20236, 67.16895, 67.1352, 
    67.1011, 67.06665, 67.03186, 66.99672, 66.96124, 66.92543, 66.88927, 
    66.85278, 66.81596, 66.7788, 66.74131, 66.70349, 66.66534, 66.62687, 
    66.58807, 66.54894, 66.5095, 66.46973, 66.42966, 66.38925, 66.34854, 
    66.30751, 66.26617, 66.22453, 66.18256, 66.1403, 66.09772, 66.05486, 
    66.01168, 65.96821, 65.92443, 65.88036, 65.836, 65.79134, 65.74638, 
    65.70114, 65.65562, 65.6098, 65.5637, 65.51731, 65.47065, 65.4237, 
    65.37647, 65.32897, 65.2812, 65.23315, 65.18482, 65.13623, 65.08736, 
    65.03824, 64.98885, 64.93919, 64.88927, 64.83908, 64.78864, 64.73795, 
    64.68699, 64.63578, 64.58432, 64.53261, 64.48065, 64.42844, 64.37598, 
    64.32328, 64.27034, 64.21716, 64.16373, 64.11006, 64.05616, 64.00202, 
    63.94765, 63.89305, 63.83821, 63.78315, 63.72786, 63.67234, 63.61659, 
    63.56062, 63.50443, 63.44802, 63.39139, 63.33455, 63.27748, 63.2202, 
    63.16271, 63.105,
  57.07566, 57.14794, 57.22011, 57.29218, 57.36412, 57.43596, 57.50769, 
    57.5793, 57.65079, 57.72218, 57.79344, 57.86459, 57.93562, 58.00652, 
    58.07731, 58.14798, 58.21853, 58.28896, 58.35925, 58.42943, 58.49948, 
    58.56941, 58.63921, 58.70888, 58.77842, 58.84783, 58.91711, 58.98626, 
    59.05527, 59.12416, 59.19291, 59.26152, 59.32999, 59.39833, 59.46653, 
    59.5346, 59.60252, 59.6703, 59.73793, 59.80542, 59.87277, 59.93998, 
    60.00703, 60.07394, 60.1407, 60.20731, 60.27377, 60.34007, 60.40623, 
    60.47223, 60.53807, 60.60376, 60.66929, 60.73466, 60.79988, 60.86493, 
    60.92982, 60.99454, 61.05911, 61.1235, 61.18774, 61.2518, 61.31569, 
    61.37942, 61.44297, 61.50635, 61.56956, 61.63259, 61.69544, 61.75812, 
    61.82062, 61.88294, 61.94508, 62.00703, 62.0688, 62.13039, 62.19179, 
    62.253, 62.31403, 62.37486, 62.4355, 62.49595, 62.55621, 62.61626, 
    62.67613, 62.73579, 62.79526, 62.85452, 62.91358, 62.97244, 63.03109, 
    63.08954, 63.14778, 63.20581, 63.26363, 63.32124, 63.37863, 63.43581, 
    63.49277, 63.54951, 63.60604, 63.66234, 63.71842, 63.77428, 63.82991, 
    63.88532, 63.94049, 63.99545, 64.05016, 64.10464, 64.1589, 64.21291, 
    64.26669, 64.32022, 64.37352, 64.42657, 64.47939, 64.53195, 64.58427, 
    64.63634, 64.68816, 64.73974, 64.79105, 64.84212, 64.89293, 64.94347, 
    64.99377, 65.04379, 65.09356, 65.14306, 65.1923, 65.24126, 65.28996, 
    65.33839, 65.38655, 65.43443, 65.48204, 65.52937, 65.57642, 65.62318, 
    65.66968, 65.71587, 65.7618, 65.80743, 65.85277, 65.89782, 65.94257, 
    65.98704, 66.0312, 66.07508, 66.11865, 66.16192, 66.20489, 66.24755, 
    66.28991, 66.33196, 66.3737, 66.41514, 66.45625, 66.49706, 66.53755, 
    66.57772, 66.61758, 66.6571, 66.69631, 66.7352, 66.77376, 66.81199, 
    66.84989, 66.88746, 66.9247, 66.96161, 66.99818, 67.03441, 67.0703, 
    67.10585, 67.14106, 67.17593, 67.21045, 67.24462, 67.27844, 67.31192, 
    67.34504, 67.37781, 67.41022, 67.44228, 67.47398, 67.50532, 67.53629, 
    67.56691, 67.59716, 67.62704, 67.65656, 67.68571, 67.71449, 67.7429, 
    67.77094, 67.79859, 67.82588, 67.85278, 67.87931, 67.90546, 67.93123, 
    67.95661, 67.98161, 68.00622, 68.03045, 68.05428, 68.07774, 68.10079, 
    68.12346, 68.14573, 68.16761, 68.18909, 68.21017, 68.23087, 68.25115, 
    68.27103, 68.29053, 68.30961, 68.32829, 68.34657, 68.36443, 68.3819, 
    68.39895, 68.4156, 68.43183, 68.44766, 68.46307, 68.47807, 68.49266, 
    68.50684, 68.5206, 68.53394, 68.54687, 68.55938, 68.57146, 68.58314, 
    68.59439, 68.60522, 68.61564, 68.62563, 68.63519, 68.64434, 68.65306, 
    68.66136, 68.66924, 68.67668, 68.68371, 68.69031, 68.69648, 68.70222, 
    68.70754, 68.71244, 68.7169, 68.72094, 68.72455, 68.72773, 68.73048, 
    68.73281, 68.7347, 68.73617, 68.73721, 68.73782, 68.738, 68.73775, 
    68.73708, 68.73597, 68.73443, 68.73247, 68.73007, 68.72726, 68.72401, 
    68.72033, 68.71622, 68.71169, 68.70673, 68.70135, 68.69553, 68.68929, 
    68.68262, 68.67554, 68.66801, 68.66007, 68.65171, 68.64292, 68.63371, 
    68.62408, 68.61402, 68.60354, 68.59264, 68.58132, 68.56958, 68.55743, 
    68.54485, 68.53186, 68.51845, 68.50462, 68.49039, 68.47573, 68.46066, 
    68.44518, 68.42929, 68.41299, 68.39628, 68.37916, 68.36163, 68.3437, 
    68.32536, 68.30662, 68.28747, 68.26792, 68.24797, 68.22762, 68.20686, 
    68.18571, 68.16417, 68.14223, 68.1199, 68.09717, 68.07405, 68.05054, 
    68.02664, 68.00235, 67.97768, 67.95262, 67.92718, 67.90135, 67.87514, 
    67.84856, 67.82159, 67.79424, 67.76653, 67.73843, 67.70997, 67.68113, 
    67.65192, 67.62234, 67.5924, 67.56209, 67.53142, 67.50038, 67.46899, 
    67.43723, 67.40512, 67.37265, 67.33982, 67.30665, 67.27312, 67.23923, 
    67.20501, 67.17043, 67.13551, 67.10025, 67.06464, 67.02869, 66.99241, 
    66.95579, 66.91883, 66.88154, 66.84392, 66.80596, 66.76768, 66.72907, 
    66.69013, 66.65087, 66.61129, 66.57139, 66.53117, 66.49063, 66.44978, 
    66.40861, 66.36713, 66.32533, 66.28323, 66.24082, 66.19811, 66.1551, 
    66.11178, 66.06816, 66.02424, 65.98003, 65.93552, 65.89071, 65.84561, 
    65.80022, 65.75455, 65.70859, 65.66234, 65.61581, 65.56899, 65.5219, 
    65.47453, 65.42688, 65.37895, 65.33075, 65.28228, 65.23354, 65.18452, 
    65.13525, 65.0857, 65.0359, 64.98582, 64.93549, 64.8849, 64.83406, 
    64.78295, 64.7316, 64.67999, 64.62813, 64.57601, 64.52365, 64.47105, 
    64.4182, 64.3651, 64.31177, 64.25819, 64.20438, 64.15033, 64.09604, 
    64.04152, 63.98677, 63.93178, 63.87657, 63.82113, 63.76546, 63.70956, 
    63.65345, 63.59711, 63.54055, 63.48377, 63.42678, 63.36956, 63.31214, 
    63.2545, 63.19664,
  57.15505, 57.22744, 57.29972, 57.3719, 57.44396, 57.51591, 57.58775, 
    57.65947, 57.73108, 57.80258, 57.87395, 57.94522, 58.01636, 58.08739, 
    58.15829, 58.22908, 58.29974, 58.37029, 58.4407, 58.511, 58.58117, 
    58.65121, 58.72113, 58.79092, 58.86058, 58.93012, 58.99952, 59.06879, 
    59.13793, 59.20694, 59.27581, 59.34455, 59.41315, 59.48161, 59.54994, 
    59.61813, 59.68617, 59.75408, 59.82184, 59.88946, 59.95694, 60.02427, 
    60.09146, 60.15849, 60.22538, 60.29213, 60.35872, 60.42515, 60.49144, 
    60.55757, 60.62355, 60.68937, 60.75504, 60.82054, 60.88589, 60.95108, 
    61.0161, 61.08096, 61.14566, 61.2102, 61.27456, 61.33876, 61.40279, 
    61.46666, 61.53035, 61.59386, 61.65721, 61.72038, 61.78338, 61.8462, 
    61.90884, 61.97129, 62.03357, 62.09567, 62.15759, 62.21931, 62.28086, 
    62.34221, 62.40338, 62.46436, 62.52514, 62.58574, 62.64614, 62.70634, 
    62.76635, 62.82616, 62.88577, 62.94518, 63.00439, 63.06339, 63.12219, 
    63.18079, 63.23917, 63.29735, 63.35532, 63.41307, 63.47061, 63.52794, 
    63.58505, 63.64194, 63.69861, 63.75507, 63.8113, 63.86731, 63.92308, 
    63.97864, 64.03397, 64.08907, 64.14394, 64.19857, 64.25297, 64.30713, 
    64.36106, 64.41475, 64.46819, 64.5214, 64.57436, 64.62708, 64.67955, 
    64.73177, 64.78374, 64.83546, 64.88693, 64.93815, 64.98911, 65.0398, 
    65.09025, 65.14043, 65.19034, 65.23999, 65.28938, 65.3385, 65.38734, 
    65.43593, 65.48423, 65.53226, 65.58002, 65.62749, 65.67469, 65.72161, 
    65.76825, 65.8146, 65.86066, 65.90644, 65.95193, 65.99712, 66.04203, 
    66.08664, 66.13095, 66.17497, 66.21869, 66.2621, 66.30521, 66.34802, 
    66.39053, 66.43272, 66.4746, 66.51617, 66.55743, 66.59838, 66.63902, 
    66.67932, 66.71931, 66.75899, 66.79833, 66.83736, 66.87605, 66.91441, 
    66.95245, 66.99016, 67.02753, 67.06457, 67.10127, 67.13763, 67.17366, 
    67.20934, 67.24468, 67.27967, 67.31432, 67.34863, 67.38257, 67.41617, 
    67.44942, 67.48231, 67.51485, 67.54703, 67.57884, 67.61031, 67.6414, 
    67.67213, 67.7025, 67.7325, 67.76213, 67.7914, 67.82028, 67.8488, 
    67.87695, 67.90472, 67.93211, 67.95912, 67.98576, 68.012, 68.03787, 
    68.06335, 68.08846, 68.11317, 68.13749, 68.16142, 68.18497, 68.20812, 
    68.23088, 68.25324, 68.27521, 68.29678, 68.31795, 68.33872, 68.35909, 
    68.37907, 68.39863, 68.41779, 68.43655, 68.4549, 68.47285, 68.49038, 
    68.50751, 68.52422, 68.54053, 68.55642, 68.5719, 68.58697, 68.60162, 
    68.61584, 68.62967, 68.64307, 68.65604, 68.66861, 68.68076, 68.69247, 
    68.70377, 68.71465, 68.72511, 68.73515, 68.74475, 68.75394, 68.7627, 
    68.77103, 68.77894, 68.78642, 68.79347, 68.8001, 68.8063, 68.81207, 
    68.81741, 68.82233, 68.82681, 68.83086, 68.83449, 68.83768, 68.84045, 
    68.84278, 68.84469, 68.84616, 68.84721, 68.84782, 68.848, 68.84775, 
    68.84707, 68.84595, 68.84441, 68.84245, 68.84004, 68.83721, 68.83395, 
    68.83025, 68.82613, 68.82158, 68.8166, 68.81119, 68.80535, 68.79908, 
    68.79239, 68.78526, 68.77772, 68.76974, 68.76134, 68.75251, 68.74326, 
    68.73358, 68.72349, 68.71296, 68.70202, 68.69065, 68.67886, 68.66665, 
    68.65402, 68.64098, 68.62751, 68.61362, 68.59933, 68.58461, 68.56948, 
    68.55393, 68.53798, 68.52161, 68.50482, 68.48763, 68.47003, 68.45203, 
    68.43361, 68.41479, 68.39556, 68.37593, 68.3559, 68.33546, 68.31463, 
    68.2934, 68.27176, 68.24973, 68.2273, 68.20448, 68.18127, 68.15767, 
    68.13367, 68.10928, 68.08451, 68.05935, 68.03381, 68.00788, 67.98157, 
    67.95487, 67.9278, 67.90035, 67.87252, 67.84431, 67.81574, 67.78679, 
    67.75747, 67.72778, 67.69772, 67.6673, 67.63651, 67.60535, 67.57384, 
    67.54196, 67.50972, 67.47713, 67.44418, 67.41088, 67.37723, 67.34322, 
    67.30886, 67.27416, 67.23911, 67.20372, 67.16798, 67.1319, 67.09549, 
    67.05873, 67.02164, 66.98421, 66.94646, 66.90837, 66.86995, 66.8312, 
    66.79213, 66.75273, 66.71301, 66.67297, 66.63261, 66.59193, 66.55093, 
    66.50962, 66.468, 66.42606, 66.38382, 66.34127, 66.29842, 66.25526, 
    66.21179, 66.16803, 66.12396, 66.07961, 66.03494, 65.99, 65.94476, 
    65.89922, 65.85339, 65.80728, 65.76089, 65.71421, 65.66724, 65.62, 
    65.57248, 65.52468, 65.47661, 65.42826, 65.37964, 65.33075, 65.28159, 
    65.23215, 65.18246, 65.13251, 65.08228, 65.03181, 64.98106, 64.93006, 
    64.87881, 64.8273, 64.77554, 64.72353, 64.67126, 64.61876, 64.566, 
    64.513, 64.45975, 64.40627, 64.35255, 64.29858, 64.24438, 64.18994, 
    64.13527, 64.08037, 64.02523, 63.96987, 63.91428, 63.85846, 63.80242, 
    63.74615, 63.68966, 63.63295, 63.57603, 63.51888, 63.46152, 63.40395, 
    63.34616, 63.28816,
  57.23429, 57.30679, 57.37918, 57.45147, 57.52364, 57.5957, 57.66765, 
    57.73949, 57.81121, 57.88282, 57.95432, 58.02569, 58.09695, 58.16809, 
    58.23911, 58.31002, 58.3808, 58.45146, 58.522, 58.59241, 58.6627, 
    58.73286, 58.8029, 58.87281, 58.9426, 59.01225, 59.08178, 59.15117, 
    59.22043, 59.28956, 59.35856, 59.42742, 59.49615, 59.56474, 59.63319, 
    59.7015, 59.76968, 59.83771, 59.9056, 59.97335, 60.04095, 60.10841, 
    60.17573, 60.2429, 60.30992, 60.37679, 60.44351, 60.51008, 60.5765, 
    60.64277, 60.70887, 60.77483, 60.84063, 60.90627, 60.97175, 61.03708, 
    61.10223, 61.16723, 61.23207, 61.29674, 61.36124, 61.42558, 61.48975, 
    61.55375, 61.61758, 61.68124, 61.74472, 61.80803, 61.87117, 61.93413, 
    61.99691, 62.05951, 62.12193, 62.18417, 62.24623, 62.3081, 62.36979, 
    62.43128, 62.4926, 62.55371, 62.61465, 62.67538, 62.73593, 62.79628, 
    62.85643, 62.91639, 62.97615, 63.0357, 63.09506, 63.15421, 63.21316, 
    63.2719, 63.33043, 63.38876, 63.44687, 63.50478, 63.56247, 63.61994, 
    63.6772, 63.73424, 63.79107, 63.84767, 63.90405, 63.96021, 64.01614, 
    64.07185, 64.12732, 64.18257, 64.23759, 64.29237, 64.34692, 64.40124, 
    64.45531, 64.50916, 64.56275, 64.61611, 64.66923, 64.72209, 64.77472, 
    64.82709, 64.87921, 64.93108, 64.9827, 65.03407, 65.08518, 65.13603, 
    65.18662, 65.23695, 65.28702, 65.33682, 65.38636, 65.43563, 65.48463, 
    65.53336, 65.58181, 65.63, 65.6779, 65.72552, 65.77287, 65.81995, 
    65.86673, 65.91322, 65.95944, 66.00536, 66.051, 66.09634, 66.1414, 
    66.18616, 66.23061, 66.27478, 66.31864, 66.36221, 66.40546, 66.44841, 
    66.49106, 66.53339, 66.57542, 66.61714, 66.65855, 66.69963, 66.7404, 
    66.78085, 66.82098, 66.86079, 66.90028, 66.93944, 66.97827, 67.01678, 
    67.05495, 67.0928, 67.1303, 67.16747, 67.20431, 67.24081, 67.27696, 
    67.31277, 67.34824, 67.38337, 67.41814, 67.45257, 67.48665, 67.52037, 
    67.55375, 67.58676, 67.61942, 67.65173, 67.68366, 67.71524, 67.74646, 
    67.77731, 67.80779, 67.83791, 67.86766, 67.89703, 67.92604, 67.95467, 
    67.98293, 68.0108, 68.0383, 68.06542, 68.09216, 68.11852, 68.14449, 
    68.17007, 68.19527, 68.22009, 68.24451, 68.26854, 68.29218, 68.31542, 
    68.33827, 68.36073, 68.38279, 68.40444, 68.4257, 68.44656, 68.46702, 
    68.48707, 68.50672, 68.52596, 68.54479, 68.56322, 68.58125, 68.59885, 
    68.61605, 68.63284, 68.64921, 68.66517, 68.68072, 68.69584, 68.71056, 
    68.72485, 68.73872, 68.75218, 68.76522, 68.77783, 68.79003, 68.8018, 
    68.81315, 68.82407, 68.83458, 68.84465, 68.8543, 68.86353, 68.87233, 
    68.8807, 68.88864, 68.89615, 68.90324, 68.90989, 68.91611, 68.92191, 
    68.92728, 68.93221, 68.93672, 68.94079, 68.94444, 68.94764, 68.95042, 
    68.95276, 68.95467, 68.95615, 68.9572, 68.95782, 68.958, 68.95775, 
    68.95706, 68.95595, 68.9544, 68.95242, 68.95, 68.94716, 68.94389, 
    68.94018, 68.93604, 68.93147, 68.92646, 68.92103, 68.91516, 68.90887, 
    68.90215, 68.89499, 68.88741, 68.8794, 68.87096, 68.8621, 68.85281, 
    68.84309, 68.83295, 68.82238, 68.81139, 68.79996, 68.78813, 68.77587, 
    68.76318, 68.75008, 68.73656, 68.72262, 68.70825, 68.69347, 68.67828, 
    68.66267, 68.64664, 68.63021, 68.61336, 68.59609, 68.57842, 68.56033, 
    68.54185, 68.52294, 68.50364, 68.48392, 68.46381, 68.44329, 68.42237, 
    68.40105, 68.37933, 68.3572, 68.33469, 68.31178, 68.28847, 68.26476, 
    68.24067, 68.21619, 68.19131, 68.16605, 68.1404, 68.11437, 68.08796, 
    68.06116, 68.03398, 68.00642, 67.97848, 67.95016, 67.92148, 67.89241, 
    67.86298, 67.83317, 67.80299, 67.77245, 67.74155, 67.71027, 67.67863, 
    67.64664, 67.61428, 67.58157, 67.54849, 67.51506, 67.48129, 67.44715, 
    67.41267, 67.37783, 67.34265, 67.30713, 67.27126, 67.23505, 67.1985, 
    67.16161, 67.12439, 67.08683, 67.04893, 67.01071, 66.97215, 66.93327, 
    66.89406, 66.85452, 66.81466, 66.77448, 66.73397, 66.69315, 66.65202, 
    66.61057, 66.56879, 66.52672, 66.48434, 66.44164, 66.39864, 66.35533, 
    66.31172, 66.26781, 66.2236, 66.17909, 66.13429, 66.0892, 66.0438, 
    65.99812, 65.95215, 65.90589, 65.85934, 65.81252, 65.7654, 65.71801, 
    65.67034, 65.62239, 65.57417, 65.52567, 65.4769, 65.42786, 65.37854, 
    65.32896, 65.27912, 65.22901, 65.17863, 65.12801, 65.07711, 65.02596, 
    64.97456, 64.9229, 64.87099, 64.81882, 64.76641, 64.71375, 64.66084, 
    64.60769, 64.55429, 64.50066, 64.44678, 64.39266, 64.33831, 64.28372, 
    64.2289, 64.17384, 64.11856, 64.06305, 64.0073, 63.95134, 63.89515, 
    63.83873, 63.78209, 63.72523, 63.66816, 63.61086, 63.55335, 63.49563, 
    63.43769, 63.37954,
  57.31336, 57.38597, 57.45848, 57.53088, 57.60316, 57.67533, 57.7474, 
    57.81935, 57.89119, 57.96291, 58.03452, 58.10601, 58.17738, 58.24864, 
    58.31978, 58.3908, 58.4617, 58.53247, 58.60313, 58.67366, 58.74407, 
    58.81436, 58.88452, 58.95455, 59.02445, 59.09423, 59.16388, 59.23339, 
    59.30278, 59.37203, 59.44115, 59.51014, 59.57899, 59.64771, 59.71629, 
    59.78473, 59.85302, 59.92118, 59.9892, 60.05708, 60.12482, 60.19241, 
    60.25985, 60.32715, 60.3943, 60.4613, 60.52816, 60.59486, 60.66141, 
    60.72781, 60.79405, 60.86014, 60.92607, 60.99185, 61.05746, 61.12292, 
    61.18822, 61.25336, 61.31833, 61.38314, 61.44778, 61.51225, 61.57656, 
    61.6407, 61.70467, 61.76847, 61.83209, 61.89554, 61.95882, 62.02192, 
    62.08484, 62.14758, 62.21015, 62.27253, 62.33473, 62.39674, 62.45857, 
    62.52022, 62.58167, 62.64294, 62.70401, 62.7649, 62.82559, 62.88608, 
    62.94638, 63.00648, 63.06639, 63.12609, 63.1856, 63.2449, 63.30399, 
    63.36288, 63.42156, 63.48003, 63.5383, 63.59635, 63.65419, 63.71181, 
    63.76923, 63.82642, 63.88339, 63.94014, 63.99667, 64.05298, 64.10906, 
    64.16492, 64.22055, 64.27595, 64.33112, 64.38605, 64.44076, 64.49522, 
    64.54945, 64.60345, 64.6572, 64.71071, 64.76397, 64.81699, 64.86977, 
    64.92229, 64.97457, 65.0266, 65.07837, 65.12988, 65.18114, 65.23215, 
    65.28289, 65.33337, 65.38359, 65.43355, 65.48324, 65.53266, 65.58181, 
    65.63069, 65.6793, 65.72763, 65.77569, 65.82346, 65.87096, 65.91818, 
    65.96511, 66.01176, 66.05813, 66.1042, 66.14999, 66.19548, 66.24068, 
    66.28558, 66.33019, 66.3745, 66.41851, 66.46222, 66.50562, 66.54872, 
    66.59151, 66.634, 66.67617, 66.71803, 66.75957, 66.8008, 66.84171, 
    66.88231, 66.92258, 66.96253, 67.00216, 67.04146, 67.08043, 67.11907, 
    67.15739, 67.19537, 67.23301, 67.27032, 67.30728, 67.34391, 67.3802, 
    67.41615, 67.45174, 67.487, 67.52191, 67.55647, 67.59067, 67.62453, 
    67.65802, 67.69116, 67.72395, 67.75637, 67.78844, 67.82014, 67.85147, 
    67.88244, 67.91305, 67.94328, 67.97314, 68.00263, 68.03175, 68.06049, 
    68.08886, 68.11685, 68.14446, 68.17169, 68.19853, 68.225, 68.25108, 
    68.27676, 68.30206, 68.32697, 68.35149, 68.37563, 68.39936, 68.4227, 
    68.44565, 68.46819, 68.49034, 68.51209, 68.53343, 68.55438, 68.57492, 
    68.59505, 68.61478, 68.63411, 68.65302, 68.67153, 68.68962, 68.70731, 
    68.72458, 68.74144, 68.75788, 68.7739, 68.78952, 68.80471, 68.81949, 
    68.83384, 68.84778, 68.86129, 68.87438, 68.88705, 68.8993, 68.91113, 
    68.92252, 68.93349, 68.94404, 68.95416, 68.96385, 68.97311, 68.98195, 
    68.99036, 68.99834, 69.00588, 69.013, 69.01968, 69.02593, 69.03175, 
    69.03715, 69.0421, 69.04662, 69.05071, 69.05437, 69.05759, 69.06039, 
    69.06274, 69.06466, 69.06615, 69.0672, 69.06782, 69.068, 69.06775, 
    69.06706, 69.06594, 69.06438, 69.06239, 69.05997, 69.05711, 69.05383, 
    69.05009, 69.04594, 69.04134, 69.03632, 69.03086, 69.02498, 69.01865, 
    69.0119, 69.00471, 68.9971, 68.98906, 68.98058, 68.97168, 68.96235, 
    68.95259, 68.9424, 68.93179, 68.92075, 68.90928, 68.89739, 68.88508, 
    68.87234, 68.85918, 68.8456, 68.8316, 68.81718, 68.80234, 68.78708, 
    68.7714, 68.7553, 68.7388, 68.72188, 68.70454, 68.68679, 68.66863, 
    68.65006, 68.63108, 68.61169, 68.5919, 68.5717, 68.55109, 68.53008, 
    68.50867, 68.48686, 68.46465, 68.44204, 68.41904, 68.39563, 68.37183, 
    68.34764, 68.32306, 68.29809, 68.27273, 68.24697, 68.22083, 68.19431, 
    68.1674, 68.14012, 68.11245, 68.0844, 68.05598, 68.02718, 67.99799, 
    67.96844, 67.93852, 67.90823, 67.87757, 67.84654, 67.81515, 67.78339, 
    67.75127, 67.71879, 67.68594, 67.65275, 67.61919, 67.58528, 67.55103, 
    67.51641, 67.48145, 67.44614, 67.41048, 67.37448, 67.33814, 67.30146, 
    67.26443, 67.22707, 67.18938, 67.15134, 67.11298, 67.07429, 67.03526, 
    66.99591, 66.95624, 66.91624, 66.87591, 66.83527, 66.7943, 66.75302, 
    66.71143, 66.66952, 66.6273, 66.58476, 66.54192, 66.49878, 66.45532, 
    66.41157, 66.36752, 66.32316, 66.2785, 66.23355, 66.1883, 66.14276, 
    66.09693, 66.05081, 66.0044, 65.95771, 65.91073, 65.86346, 65.81593, 
    65.7681, 65.72, 65.67162, 65.62298, 65.57405, 65.52486, 65.4754, 
    65.42567, 65.37566, 65.32541, 65.27488, 65.2241, 65.17306, 65.12175, 
    65.0702, 65.01838, 64.96632, 64.914, 64.86143, 64.80862, 64.75556, 
    64.70226, 64.64871, 64.59492, 64.54089, 64.48663, 64.43212, 64.37738, 
    64.32241, 64.2672, 64.21177, 64.15611, 64.10021, 64.04409, 63.98775, 
    63.93118, 63.87439, 63.81738, 63.76016, 63.70271, 63.64505, 63.58718, 
    63.52909, 63.4708,
  57.39228, 57.465, 57.53762, 57.61013, 57.68253, 57.75481, 57.82698, 
    57.89905, 57.971, 58.04284, 58.11456, 58.18616, 58.25766, 58.32903, 
    58.40028, 58.47142, 58.54244, 58.61333, 58.68411, 58.75476, 58.82529, 
    58.89569, 58.96597, 59.03613, 59.10615, 59.17605, 59.24582, 59.31546, 
    59.38497, 59.45435, 59.52359, 59.5927, 59.66168, 59.73052, 59.79922, 
    59.86779, 59.93622, 60.00451, 60.07265, 60.14066, 60.20853, 60.27625, 
    60.34382, 60.41125, 60.47853, 60.54567, 60.61265, 60.67949, 60.74617, 
    60.8127, 60.87908, 60.9453, 61.01137, 61.07728, 61.14303, 61.20862, 
    61.27406, 61.33933, 61.40444, 61.46938, 61.53416, 61.59878, 61.66322, 
    61.7275, 61.79161, 61.85555, 61.91932, 61.98291, 62.04632, 62.10956, 
    62.17263, 62.23551, 62.29822, 62.36074, 62.42309, 62.48524, 62.54722, 
    62.60901, 62.67061, 62.73202, 62.79324, 62.85427, 62.9151, 62.97575, 
    63.03619, 63.09644, 63.15649, 63.21635, 63.276, 63.33545, 63.39469, 
    63.45373, 63.51256, 63.57118, 63.62959, 63.6878, 63.74578, 63.80356, 
    63.86112, 63.91846, 63.97559, 64.03249, 64.08917, 64.14563, 64.20187, 
    64.25787, 64.31366, 64.36921, 64.42453, 64.47962, 64.53448, 64.5891, 
    64.64348, 64.69762, 64.75153, 64.80518, 64.8586, 64.91178, 64.96471, 
    65.01739, 65.06982, 65.12199, 65.17392, 65.22559, 65.277, 65.32816, 
    65.37905, 65.42969, 65.48006, 65.53017, 65.58001, 65.62959, 65.67889, 
    65.72792, 65.77668, 65.82516, 65.87337, 65.9213, 65.96895, 66.01632, 
    66.06341, 66.11021, 66.15672, 66.20294, 66.24888, 66.29452, 66.33987, 
    66.38493, 66.42968, 66.47414, 66.5183, 66.56215, 66.60571, 66.64895, 
    66.69189, 66.73451, 66.77683, 66.81883, 66.86053, 66.9019, 66.94296, 
    66.9837, 67.02411, 67.0642, 67.10397, 67.1434, 67.18252, 67.2213, 
    67.25975, 67.29787, 67.33565, 67.37309, 67.41019, 67.44696, 67.48338, 
    67.51946, 67.55519, 67.59058, 67.62562, 67.6603, 67.69464, 67.72862, 
    67.76225, 67.79552, 67.82842, 67.86097, 67.89316, 67.92498, 67.95644, 
    67.98753, 68.01825, 68.04861, 68.07858, 68.10819, 68.13743, 68.16628, 
    68.19476, 68.22286, 68.25058, 68.27792, 68.30487, 68.33144, 68.35762, 
    68.38342, 68.40882, 68.43384, 68.45846, 68.48268, 68.50652, 68.52995, 
    68.55299, 68.57563, 68.59787, 68.61971, 68.64114, 68.66218, 68.68281, 
    68.70303, 68.72284, 68.74224, 68.76124, 68.77982, 68.79799, 68.81575, 
    68.83309, 68.85002, 68.86653, 68.88263, 68.89831, 68.91357, 68.92841, 
    68.94282, 68.95682, 68.97039, 68.98354, 68.99626, 69.00857, 69.02044, 
    69.03188, 69.04291, 69.0535, 69.06366, 69.07339, 69.0827, 69.09158, 
    69.10002, 69.10803, 69.11561, 69.12276, 69.12947, 69.13575, 69.14159, 
    69.14701, 69.15199, 69.15653, 69.16064, 69.16431, 69.16755, 69.17035, 
    69.17271, 69.17464, 69.17614, 69.17719, 69.17782, 69.178, 69.17775, 
    69.17706, 69.17593, 69.17437, 69.17237, 69.16994, 69.16707, 69.16376, 
    69.16002, 69.15584, 69.15123, 69.14618, 69.1407, 69.13479, 69.12843, 
    69.12165, 69.11444, 69.10679, 69.09871, 69.0902, 69.08126, 69.07188, 
    69.06208, 69.05185, 69.04119, 69.03011, 69.01859, 69.00665, 68.99428, 
    68.98149, 68.96827, 68.95463, 68.94057, 68.92609, 68.91118, 68.89586, 
    68.88011, 68.86395, 68.84737, 68.83038, 68.81297, 68.79514, 68.77691, 
    68.75826, 68.7392, 68.71973, 68.69985, 68.67957, 68.65887, 68.63778, 
    68.61628, 68.59438, 68.57207, 68.54938, 68.52628, 68.50277, 68.47887, 
    68.45459, 68.4299, 68.40483, 68.37936, 68.35351, 68.32726, 68.30064, 
    68.27362, 68.24622, 68.21844, 68.19028, 68.16174, 68.13283, 68.10354, 
    68.07387, 68.04383, 68.01342, 67.98264, 67.95148, 67.91998, 67.88809, 
    67.85585, 67.82324, 67.79028, 67.75695, 67.72327, 67.68923, 67.65484, 
    67.6201, 67.58501, 67.54957, 67.51378, 67.47765, 67.44117, 67.40435, 
    67.36719, 67.32969, 67.29185, 67.25369, 67.21519, 67.17635, 67.13719, 
    67.09769, 67.05788, 67.01774, 66.97727, 66.93649, 66.89538, 66.85395, 
    66.81221, 66.77016, 66.72779, 66.68511, 66.64213, 66.59883, 66.55524, 
    66.51133, 66.46712, 66.42262, 66.37782, 66.33272, 66.28732, 66.24163, 
    66.19565, 66.14938, 66.10282, 66.05598, 66.00884, 65.96143, 65.91373, 
    65.86576, 65.81751, 65.76898, 65.72018, 65.6711, 65.62176, 65.57214, 
    65.52226, 65.47211, 65.4217, 65.37102, 65.32008, 65.26888, 65.21743, 
    65.16572, 65.11375, 65.06154, 65.00907, 64.95635, 64.90338, 64.85017, 
    64.79671, 64.74301, 64.68907, 64.63489, 64.58047, 64.52581, 64.47092, 
    64.41579, 64.36044, 64.30485, 64.24903, 64.19299, 64.13672, 64.08022, 
    64.02351, 63.96656, 63.90941, 63.85203, 63.79444, 63.73663, 63.6786, 
    63.62037, 63.56192,
  57.47104, 57.54387, 57.6166, 57.68922, 57.76173, 57.83413, 57.90641, 
    57.97859, 58.05065, 58.1226, 58.19444, 58.26616, 58.33777, 58.40926, 
    58.48063, 58.55188, 58.62302, 58.69403, 58.76493, 58.8357, 58.90635, 
    58.97687, 59.04727, 59.11755, 59.18769, 59.25771, 59.32761, 59.39737, 
    59.467, 59.5365, 59.60587, 59.67511, 59.74421, 59.81318, 59.88201, 
    59.9507, 60.01926, 60.08767, 60.15595, 60.22409, 60.29208, 60.35993, 
    60.42763, 60.49519, 60.56261, 60.62987, 60.69699, 60.76395, 60.83077, 
    60.89744, 60.96395, 61.0303, 61.09651, 61.16255, 61.22844, 61.29417, 
    61.35974, 61.42515, 61.49039, 61.55548, 61.6204, 61.68515, 61.74974, 
    61.81416, 61.8784, 61.94248, 62.00639, 62.07012, 62.13368, 62.19706, 
    62.26027, 62.3233, 62.38615, 62.44881, 62.5113, 62.5736, 62.63572, 
    62.69765, 62.7594, 62.82096, 62.88232, 62.9435, 63.00449, 63.06527, 
    63.12587, 63.18626, 63.24646, 63.30647, 63.36626, 63.42586, 63.48525, 
    63.54444, 63.60342, 63.66219, 63.72076, 63.77911, 63.83725, 63.89518, 
    63.95288, 64.01038, 64.06766, 64.12471, 64.18154, 64.23816, 64.29454, 
    64.35071, 64.40664, 64.46234, 64.51781, 64.57306, 64.62807, 64.68284, 
    64.73737, 64.79167, 64.84573, 64.89954, 64.95312, 65.00645, 65.05952, 
    65.11236, 65.16495, 65.21728, 65.26936, 65.32118, 65.37275, 65.42406, 
    65.47511, 65.52589, 65.57642, 65.62669, 65.67667, 65.7264, 65.77586, 
    65.82504, 65.87396, 65.92259, 65.97095, 66.01904, 66.06684, 66.11436, 
    66.1616, 66.20855, 66.25522, 66.30159, 66.34768, 66.39347, 66.43897, 
    66.48418, 66.52908, 66.57368, 66.618, 66.66199, 66.7057, 66.74909, 
    66.79218, 66.83495, 66.87741, 66.91956, 66.9614, 67.00292, 67.04412, 
    67.085, 67.12556, 67.16579, 67.2057, 67.24529, 67.28454, 67.32346, 
    67.36205, 67.4003, 67.43822, 67.4758, 67.51305, 67.54994, 67.5865, 
    67.62271, 67.65858, 67.6941, 67.72927, 67.76409, 67.79855, 67.83266, 
    67.86642, 67.89981, 67.93285, 67.96552, 67.99783, 68.02978, 68.06136, 
    68.09258, 68.12341, 68.15388, 68.18399, 68.21371, 68.24306, 68.27203, 
    68.30063, 68.32883, 68.35667, 68.38412, 68.41118, 68.43785, 68.46414, 
    68.49004, 68.51555, 68.54066, 68.56538, 68.58971, 68.61365, 68.63718, 
    68.66031, 68.68304, 68.70538, 68.72731, 68.74883, 68.76995, 68.79066, 
    68.81097, 68.83087, 68.85036, 68.86943, 68.88809, 68.90634, 68.92417, 
    68.94159, 68.9586, 68.97517, 68.99134, 69.00709, 69.02241, 69.03732, 
    69.0518, 69.06585, 69.07948, 69.09269, 69.10547, 69.11782, 69.12975, 
    69.14124, 69.15231, 69.16295, 69.17316, 69.18294, 69.19228, 69.20119, 
    69.20967, 69.21772, 69.22533, 69.23251, 69.23926, 69.24557, 69.25143, 
    69.25687, 69.26187, 69.26643, 69.27056, 69.27425, 69.2775, 69.28032, 
    69.28269, 69.28463, 69.28613, 69.28719, 69.28781, 69.288, 69.28774, 
    69.28706, 69.28592, 69.28436, 69.28235, 69.2799, 69.27702, 69.2737, 
    69.26994, 69.26575, 69.26111, 69.25604, 69.25053, 69.2446, 69.23822, 
    69.23141, 69.22416, 69.21648, 69.20836, 69.19981, 69.19083, 69.18142, 
    69.17157, 69.16129, 69.15059, 69.13945, 69.12789, 69.1159, 69.10347, 
    69.09062, 69.07735, 69.06365, 69.04953, 69.03498, 69.02001, 69.00462, 
    68.98882, 68.97258, 68.95593, 68.93887, 68.92138, 68.90348, 68.88517, 
    68.86644, 68.8473, 68.82775, 68.80779, 68.78741, 68.76664, 68.74545, 
    68.72387, 68.70187, 68.67947, 68.65668, 68.63348, 68.60989, 68.58589, 
    68.5615, 68.53672, 68.51154, 68.48597, 68.46001, 68.43366, 68.40692, 
    68.3798, 68.35229, 68.3244, 68.29613, 68.26747, 68.23844, 68.20904, 
    68.17925, 68.14909, 68.11856, 68.08766, 68.05639, 68.02475, 67.99274, 
    67.96038, 67.92764, 67.89455, 67.8611, 67.82729, 67.79312, 67.75861, 
    67.72373, 67.68851, 67.65293, 67.61701, 67.58074, 67.54413, 67.50717, 
    67.46988, 67.43224, 67.39427, 67.35596, 67.31732, 67.27835, 67.23904, 
    67.19941, 67.15945, 67.11916, 67.07855, 67.03762, 66.99638, 66.9548, 
    66.91292, 66.87072, 66.8282, 66.78538, 66.74225, 66.69881, 66.65506, 
    66.61101, 66.56665, 66.522, 66.47704, 66.43179, 66.38625, 66.34041, 
    66.29427, 66.24786, 66.20114, 66.15414, 66.10686, 66.0593, 66.01145, 
    65.96333, 65.91492, 65.86624, 65.81728, 65.76806, 65.71856, 65.66879, 
    65.61875, 65.56844, 65.51788, 65.46705, 65.41595, 65.36461, 65.313, 
    65.26113, 65.20901, 65.15665, 65.10402, 65.05115, 64.99802, 64.94466, 
    64.89105, 64.8372, 64.7831, 64.72877, 64.67419, 64.61938, 64.56434, 
    64.50906, 64.45354, 64.3978, 64.34184, 64.28564, 64.22922, 64.17257, 
    64.1157, 64.05861, 64.0013, 63.94377, 63.88602, 63.82807, 63.76989, 
    63.71151, 63.65291,
  57.54963, 57.62258, 57.69542, 57.76815, 57.84077, 57.91328, 57.98568, 
    58.05797, 58.13015, 58.20221, 58.27416, 58.346, 58.41772, 58.48933, 
    58.56081, 58.63219, 58.70344, 58.77457, 58.84558, 58.91647, 58.98724, 
    59.05789, 59.12841, 59.1988, 59.26907, 59.33922, 59.40923, 59.47912, 
    59.54887, 59.6185, 59.688, 59.75735, 59.82658, 59.89568, 59.96463, 
    60.03345, 60.10214, 60.17068, 60.23909, 60.30735, 60.37547, 60.44345, 
    60.51129, 60.57898, 60.64652, 60.71392, 60.78117, 60.84827, 60.91522, 
    60.98202, 61.04866, 61.11516, 61.1815, 61.24768, 61.3137, 61.37957, 
    61.44527, 61.51082, 61.5762, 61.64143, 61.70648, 61.77137, 61.8361, 
    61.90066, 61.96505, 62.02927, 62.09332, 62.15719, 62.22089, 62.28442, 
    62.34776, 62.41093, 62.47393, 62.53674, 62.59937, 62.66182, 62.72408, 
    62.78616, 62.84805, 62.90976, 62.97127, 63.03259, 63.09372, 63.15466, 
    63.2154, 63.27595, 63.33629, 63.39644, 63.45639, 63.51614, 63.57568, 
    63.63501, 63.69415, 63.75307, 63.81178, 63.87029, 63.92858, 63.98666, 
    64.04452, 64.10217, 64.15959, 64.2168, 64.27379, 64.33055, 64.38709, 
    64.44341, 64.4995, 64.55535, 64.61098, 64.66637, 64.72153, 64.77647, 
    64.83115, 64.8856, 64.93982, 64.99379, 65.04752, 65.101, 65.15424, 
    65.20722, 65.25996, 65.31245, 65.36468, 65.41666, 65.46838, 65.51984, 
    65.57105, 65.62199, 65.67268, 65.72309, 65.77324, 65.82312, 65.87273, 
    65.92207, 65.97114, 66.01993, 66.06844, 66.11668, 66.16463, 66.2123, 
    66.2597, 66.3068, 66.35361, 66.40015, 66.44638, 66.49233, 66.53798, 
    66.58334, 66.6284, 66.67315, 66.71761, 66.76176, 66.8056, 66.84915, 
    66.89238, 66.9353, 66.97791, 67.02021, 67.06219, 67.10386, 67.1452, 
    67.18623, 67.22694, 67.26731, 67.30737, 67.34708, 67.38648, 67.42554, 
    67.46427, 67.50267, 67.54073, 67.57845, 67.61583, 67.65286, 67.68956, 
    67.72591, 67.76191, 67.79756, 67.83286, 67.86781, 67.90241, 67.93665, 
    67.97054, 68.00406, 68.03722, 68.07002, 68.10246, 68.13453, 68.16624, 
    68.19757, 68.22853, 68.25912, 68.28934, 68.31918, 68.34866, 68.37774, 
    68.40645, 68.43478, 68.46272, 68.49027, 68.51745, 68.54423, 68.57063, 
    68.59663, 68.62225, 68.64746, 68.67229, 68.69672, 68.72074, 68.74438, 
    68.76761, 68.79044, 68.81286, 68.83488, 68.8565, 68.87771, 68.89851, 
    68.9189, 68.93888, 68.95845, 68.97761, 68.99635, 69.01467, 69.03259, 
    69.05008, 69.06715, 69.08381, 69.10004, 69.11585, 69.13124, 69.14621, 
    69.16075, 69.17487, 69.18856, 69.20183, 69.21466, 69.22707, 69.23904, 
    69.2506, 69.26171, 69.2724, 69.28265, 69.29247, 69.30186, 69.31081, 
    69.31933, 69.32741, 69.33505, 69.34226, 69.34904, 69.35538, 69.36127, 
    69.36674, 69.37176, 69.37634, 69.38049, 69.38419, 69.38746, 69.39028, 
    69.39267, 69.39462, 69.39612, 69.39719, 69.39781, 69.39799, 69.39774, 
    69.39705, 69.39591, 69.39433, 69.39232, 69.38986, 69.38697, 69.38364, 
    69.37986, 69.37564, 69.37099, 69.3659, 69.36037, 69.3544, 69.348, 
    69.34116, 69.33388, 69.32616, 69.31801, 69.30942, 69.3004, 69.29095, 
    69.28106, 69.27074, 69.25998, 69.24879, 69.23718, 69.22514, 69.21266, 
    69.19975, 69.18642, 69.17267, 69.15848, 69.14387, 69.12884, 69.11338, 
    69.0975, 69.0812, 69.06448, 69.04734, 69.02978, 69.0118, 68.99341, 
    68.9746, 68.95538, 68.93575, 68.9157, 68.89525, 68.87438, 68.8531, 
    68.83143, 68.80934, 68.78685, 68.76396, 68.74066, 68.71697, 68.69288, 
    68.66839, 68.6435, 68.61822, 68.59254, 68.56647, 68.54002, 68.51318, 
    68.48594, 68.45832, 68.43032, 68.40193, 68.37316, 68.34402, 68.31449, 
    68.28459, 68.25431, 68.22366, 68.19263, 68.16124, 68.12948, 68.09735, 
    68.06486, 68.032, 67.99878, 67.96519, 67.93126, 67.89696, 67.86231, 
    67.8273, 67.79195, 67.75624, 67.72018, 67.68378, 67.64703, 67.60994, 
    67.5725, 67.53473, 67.49662, 67.45817, 67.41939, 67.38027, 67.34083, 
    67.30105, 67.26095, 67.22052, 67.17976, 67.13869, 67.09729, 67.05557, 
    67.01354, 66.9712, 66.92854, 66.88557, 66.84229, 66.79869, 66.75479, 
    66.71059, 66.66609, 66.62128, 66.57618, 66.53078, 66.48508, 66.43909, 
    66.39281, 66.34623, 66.29937, 66.25222, 66.20478, 66.15707, 66.10906, 
    66.06078, 66.01223, 65.96339, 65.91428, 65.8649, 65.81525, 65.76532, 
    65.71513, 65.66467, 65.61395, 65.56297, 65.51172, 65.46021, 65.40845, 
    65.35643, 65.30416, 65.25163, 65.19885, 65.14583, 65.09255, 65.03903, 
    64.98527, 64.93126, 64.87701, 64.82252, 64.76779, 64.71283, 64.65763, 
    64.6022, 64.54653, 64.49064, 64.43452, 64.37817, 64.32159, 64.26479, 
    64.20776, 64.15052, 64.09306, 64.03538, 63.97749, 63.91937, 63.86105, 
    63.80251, 63.74376,
  57.62807, 57.70112, 57.77407, 57.84691, 57.91964, 57.99227, 58.06478, 
    58.13718, 58.20947, 58.28165, 58.35372, 58.42567, 58.49751, 58.56923, 
    58.64084, 58.71233, 58.7837, 58.85495, 58.92608, 58.99709, 59.06798, 
    59.13874, 59.20938, 59.2799, 59.35029, 59.42056, 59.4907, 59.56071, 
    59.63058, 59.70034, 59.76995, 59.83944, 59.90879, 59.97802, 60.0471, 
    60.11605, 60.18486, 60.25353, 60.32206, 60.39046, 60.45871, 60.52682, 
    60.59479, 60.66261, 60.73029, 60.79781, 60.8652, 60.93243, 60.99951, 
    61.06644, 61.13323, 61.19985, 61.26633, 61.33265, 61.3988, 61.46481, 
    61.53065, 61.59634, 61.66186, 61.72722, 61.79242, 61.85744, 61.92231, 
    61.98701, 62.05154, 62.1159, 62.18009, 62.24411, 62.30795, 62.37162, 
    62.43511, 62.49842, 62.56156, 62.62452, 62.68729, 62.74989, 62.8123, 
    62.87452, 62.93656, 62.99841, 63.06007, 63.12154, 63.18282, 63.2439, 
    63.30479, 63.36549, 63.42598, 63.48628, 63.54638, 63.60627, 63.66597, 
    63.72545, 63.78474, 63.84381, 63.90268, 63.96133, 64.01978, 64.078, 
    64.13602, 64.19382, 64.2514, 64.30876, 64.3659, 64.42282, 64.47952, 
    64.53598, 64.59222, 64.64823, 64.70402, 64.75957, 64.81488, 64.86996, 
    64.92481, 64.97942, 65.03378, 65.08791, 65.14179, 65.19543, 65.24882, 
    65.30196, 65.35486, 65.4075, 65.45988, 65.51202, 65.5639, 65.61552, 
    65.66688, 65.71798, 65.76881, 65.81939, 65.86969, 65.91972, 65.96949, 
    66.01899, 66.06821, 66.11716, 66.16582, 66.21421, 66.26232, 66.31015, 
    66.3577, 66.40495, 66.45193, 66.4986, 66.545, 66.59109, 66.63689, 
    66.6824, 66.72761, 66.77252, 66.81713, 66.86143, 66.90543, 66.94912, 
    66.9925, 67.03558, 67.07834, 67.12078, 67.16291, 67.20472, 67.24622, 
    67.28738, 67.32823, 67.36876, 67.40895, 67.44882, 67.48836, 67.52757, 
    67.56644, 67.60497, 67.64317, 67.68103, 67.71854, 67.75572, 67.79255, 
    67.82904, 67.86517, 67.90096, 67.9364, 67.97148, 68.00621, 68.04058, 
    68.07459, 68.10825, 68.14154, 68.17447, 68.20703, 68.23923, 68.27106, 
    68.30251, 68.3336, 68.36432, 68.39465, 68.42462, 68.4542, 68.48341, 
    68.51223, 68.54067, 68.56873, 68.5964, 68.62368, 68.65057, 68.67708, 
    68.70319, 68.7289, 68.75423, 68.77916, 68.80369, 68.82782, 68.85155, 
    68.87488, 68.8978, 68.92032, 68.94244, 68.96414, 68.98544, 69.00632, 
    69.02681, 69.04688, 69.06653, 69.08576, 69.10458, 69.12299, 69.14098, 
    69.15855, 69.1757, 69.19242, 69.20872, 69.22461, 69.24007, 69.2551, 
    69.26971, 69.28388, 69.29763, 69.31095, 69.32384, 69.33631, 69.34834, 
    69.35994, 69.3711, 69.38184, 69.39214, 69.402, 69.41143, 69.42042, 
    69.42898, 69.4371, 69.44477, 69.45202, 69.45882, 69.46519, 69.47111, 
    69.47659, 69.48164, 69.48624, 69.49041, 69.49413, 69.49741, 69.50024, 
    69.50265, 69.5046, 69.50611, 69.50719, 69.50781, 69.508, 69.50774, 
    69.50704, 69.50591, 69.50432, 69.5023, 69.49982, 69.49692, 69.49357, 
    69.48978, 69.48554, 69.48087, 69.47575, 69.4702, 69.46421, 69.45777, 
    69.4509, 69.44359, 69.43584, 69.42765, 69.41903, 69.40997, 69.40047, 
    69.39053, 69.38017, 69.36937, 69.35813, 69.34647, 69.33437, 69.32184, 
    69.30888, 69.29549, 69.28167, 69.26742, 69.25275, 69.23765, 69.22212, 
    69.20618, 69.1898, 69.17301, 69.15579, 69.13816, 69.12011, 69.10164, 
    69.08275, 69.06345, 69.04372, 69.0236, 69.00305, 68.98209, 68.96073, 
    68.93896, 68.91679, 68.8942, 68.87121, 68.84782, 68.82403, 68.79984, 
    68.77524, 68.75025, 68.72486, 68.69908, 68.67291, 68.64635, 68.61939, 
    68.59205, 68.56432, 68.53619, 68.5077, 68.47881, 68.44955, 68.41991, 
    68.38988, 68.35948, 68.32871, 68.29756, 68.26604, 68.23416, 68.2019, 
    68.16929, 68.1363, 68.10295, 68.06924, 68.03517, 68.00074, 67.96596, 
    67.93082, 67.89532, 67.85948, 67.82329, 67.78675, 67.74986, 67.71263, 
    67.67506, 67.63715, 67.59889, 67.56031, 67.52139, 67.48212, 67.44254, 
    67.40262, 67.36237, 67.32179, 67.28089, 67.23967, 67.19813, 67.15627, 
    67.11409, 67.07159, 67.02879, 66.98566, 66.94223, 66.89849, 66.85445, 
    66.81009, 66.76543, 66.72048, 66.67522, 66.62967, 66.58382, 66.53767, 
    66.49124, 66.44451, 66.3975, 66.3502, 66.3026, 66.25473, 66.20658, 
    66.15814, 66.10943, 66.06044, 66.01118, 65.96164, 65.91183, 65.86175, 
    65.8114, 65.76079, 65.70992, 65.65878, 65.60737, 65.55571, 65.50379, 
    65.45161, 65.39919, 65.3465, 65.29357, 65.24039, 65.18696, 65.13329, 
    65.07936, 65.0252, 64.97079, 64.91615, 64.86127, 64.80614, 64.75079, 
    64.69521, 64.63939, 64.58334, 64.52706, 64.47056, 64.41383, 64.35688, 
    64.2997, 64.2423, 64.18469, 64.12685, 64.06881, 64.01054, 63.95207, 
    63.89338, 63.83448,
  57.70634, 57.7795, 57.85256, 57.92551, 57.99836, 58.07109, 58.14372, 
    58.21624, 58.28864, 58.36094, 58.43312, 58.50518, 58.57714, 58.64898, 
    58.7207, 58.7923, 58.86379, 58.93516, 59.00641, 59.07754, 59.14855, 
    59.21943, 59.2902, 59.36084, 59.43135, 59.50174, 59.572, 59.64213, 
    59.71214, 59.78201, 59.85175, 59.92137, 59.99085, 60.06019, 60.12941, 
    60.19848, 60.26742, 60.33622, 60.40488, 60.47341, 60.54179, 60.61003, 
    60.67813, 60.74608, 60.81389, 60.88155, 60.94907, 61.01643, 61.08365, 
    61.15071, 61.21763, 61.28439, 61.351, 61.41745, 61.48375, 61.54989, 
    61.61588, 61.6817, 61.74736, 61.81286, 61.87819, 61.94336, 62.00837, 
    62.07321, 62.13788, 62.20238, 62.26671, 62.33087, 62.39486, 62.45867, 
    62.5223, 62.58577, 62.64905, 62.71215, 62.77507, 62.83781, 62.90036, 
    62.96273, 63.02492, 63.08691, 63.14872, 63.21034, 63.27177, 63.333, 
    63.39404, 63.45488, 63.51553, 63.57598, 63.63623, 63.69627, 63.75611, 
    63.81575, 63.87519, 63.93441, 63.99343, 64.05224, 64.11083, 64.16922, 
    64.22739, 64.28534, 64.34307, 64.40059, 64.45788, 64.51495, 64.5718, 
    64.62843, 64.68482, 64.74099, 64.79692, 64.85263, 64.9081, 64.96334, 
    65.01834, 65.0731, 65.12762, 65.18191, 65.23595, 65.28974, 65.34328, 
    65.39658, 65.44964, 65.50243, 65.55498, 65.60727, 65.6593, 65.71108, 
    65.7626, 65.81385, 65.86485, 65.91557, 65.96603, 66.01623, 66.06615, 
    66.1158, 66.16518, 66.21428, 66.2631, 66.31165, 66.35991, 66.4079, 
    66.4556, 66.50301, 66.55013, 66.59697, 66.64351, 66.68976, 66.73572, 
    66.78138, 66.82674, 66.8718, 66.91656, 66.96101, 67.00517, 67.049, 
    67.09254, 67.13577, 67.17867, 67.22127, 67.26354, 67.3055, 67.34715, 
    67.38846, 67.42946, 67.47012, 67.51047, 67.55048, 67.59016, 67.62951, 
    67.66852, 67.7072, 67.74554, 67.78354, 67.8212, 67.85851, 67.89548, 
    67.93211, 67.96838, 68.0043, 68.03987, 68.07509, 68.10995, 68.14445, 
    68.1786, 68.21239, 68.24581, 68.27886, 68.31155, 68.34388, 68.37583, 
    68.40742, 68.43863, 68.46947, 68.49992, 68.53001, 68.55971, 68.58904, 
    68.61797, 68.64653, 68.6747, 68.70248, 68.72987, 68.75688, 68.78349, 
    68.80972, 68.83554, 68.86096, 68.88599, 68.91063, 68.93486, 68.95869, 
    68.98212, 69.00513, 69.02775, 69.04996, 69.07176, 69.09315, 69.11413, 
    69.13469, 69.15485, 69.17458, 69.1939, 69.21281, 69.23129, 69.24936, 
    69.267, 69.28423, 69.30103, 69.3174, 69.33335, 69.34888, 69.36398, 
    69.37864, 69.39288, 69.40669, 69.42007, 69.43303, 69.44554, 69.45763, 
    69.46928, 69.48049, 69.49127, 69.50162, 69.51153, 69.521, 69.53003, 
    69.53862, 69.54678, 69.55449, 69.56177, 69.5686, 69.57499, 69.58094, 
    69.58646, 69.59152, 69.59615, 69.60033, 69.60406, 69.60736, 69.61021, 
    69.61262, 69.61459, 69.6161, 69.61718, 69.61781, 69.618, 69.61774, 
    69.61704, 69.61589, 69.6143, 69.61227, 69.60979, 69.60687, 69.6035, 
    69.59969, 69.59544, 69.59075, 69.58561, 69.58003, 69.57401, 69.56755, 
    69.56065, 69.5533, 69.54552, 69.53729, 69.52863, 69.51952, 69.50999, 
    69.50001, 69.48959, 69.47874, 69.46746, 69.45574, 69.44359, 69.43101, 
    69.41799, 69.40454, 69.39066, 69.37635, 69.36161, 69.34644, 69.33086, 
    69.31483, 69.29839, 69.28152, 69.26424, 69.24653, 69.22839, 69.20985, 
    69.19087, 69.17149, 69.15169, 69.13147, 69.11083, 69.08979, 69.06834, 
    69.04647, 69.0242, 69.00152, 68.97844, 68.95495, 68.93105, 68.90676, 
    68.88206, 68.85697, 68.83148, 68.80559, 68.77931, 68.75263, 68.72557, 
    68.69811, 68.67027, 68.64204, 68.61342, 68.58442, 68.55504, 68.52528, 
    68.49513, 68.46461, 68.43372, 68.40244, 68.3708, 68.33879, 68.30641, 
    68.27366, 68.24055, 68.20707, 68.17323, 68.13902, 68.10446, 68.06954, 
    68.03427, 67.99864, 67.96266, 67.92634, 67.88966, 67.85263, 67.81526, 
    67.77755, 67.73949, 67.7011, 67.66237, 67.62331, 67.5839, 67.54417, 
    67.5041, 67.46371, 67.42299, 67.38194, 67.34058, 67.29889, 67.25687, 
    67.21455, 67.17191, 67.12894, 67.08568, 67.04209, 66.9982, 66.954, 
    66.9095, 66.86469, 66.81959, 66.77418, 66.72847, 66.68246, 66.63617, 
    66.58958, 66.54269, 66.49553, 66.44807, 66.40032, 66.35229, 66.30399, 
    66.25539, 66.20653, 66.15739, 66.10796, 66.05827, 66.00831, 65.95807, 
    65.90757, 65.8568, 65.80576, 65.75446, 65.70291, 65.65109, 65.59901, 
    65.54668, 65.4941, 65.44126, 65.38817, 65.33483, 65.28124, 65.22741, 
    65.17333, 65.11902, 65.06445, 65.00965, 64.95461, 64.89935, 64.84383, 
    64.78809, 64.73212, 64.67591, 64.61948, 64.56282, 64.50594, 64.44883, 
    64.3915, 64.33395, 64.27618, 64.2182, 64.16, 64.10158, 64.04295, 
    63.98411, 63.92506,
  57.78444, 57.85772, 57.93089, 58.00395, 58.0769, 58.14975, 58.22249, 
    58.29512, 58.36764, 58.44005, 58.51234, 58.58453, 58.6566, 58.72855, 
    58.80039, 58.87212, 58.94372, 59.01521, 59.08658, 59.15783, 59.22895, 
    59.29996, 59.37085, 59.44161, 59.51224, 59.58275, 59.65314, 59.72339, 
    59.79352, 59.86352, 59.93339, 60.00313, 60.07273, 60.14221, 60.21155, 
    60.28075, 60.34982, 60.41875, 60.48754, 60.55619, 60.62471, 60.69308, 
    60.7613, 60.82939, 60.89733, 60.96513, 61.03277, 61.10027, 61.16763, 
    61.23483, 61.30188, 61.36877, 61.43552, 61.50211, 61.56854, 61.63482, 
    61.70094, 61.7669, 61.8327, 61.89834, 61.96381, 62.02913, 62.09427, 
    62.15925, 62.22407, 62.28871, 62.35318, 62.41748, 62.48161, 62.54557, 
    62.60935, 62.67295, 62.73638, 62.79963, 62.86269, 62.92558, 62.98828, 
    63.0508, 63.11313, 63.17527, 63.23723, 63.299, 63.36057, 63.42196, 
    63.48314, 63.54414, 63.60493, 63.66553, 63.72593, 63.78613, 63.84612, 
    63.90591, 63.9655, 64.02488, 64.08405, 64.14301, 64.20176, 64.26029, 
    64.31861, 64.37672, 64.43461, 64.49228, 64.54973, 64.60696, 64.66396, 
    64.72073, 64.77729, 64.83361, 64.8897, 64.94556, 65.00119, 65.05659, 
    65.11174, 65.16666, 65.22134, 65.27578, 65.32998, 65.38393, 65.43763, 
    65.49109, 65.5443, 65.59725, 65.64996, 65.7024, 65.75459, 65.80653, 
    65.8582, 65.90961, 65.96076, 66.01165, 66.06226, 66.11262, 66.1627, 
    66.2125, 66.26204, 66.31129, 66.36028, 66.40897, 66.4574, 66.50554, 
    66.55339, 66.60096, 66.64824, 66.69523, 66.74193, 66.78834, 66.83444, 
    66.88026, 66.92577, 66.97099, 67.0159, 67.06051, 67.10481, 67.1488, 
    67.19249, 67.23586, 67.27892, 67.32166, 67.3641, 67.4062, 67.44799, 
    67.48946, 67.5306, 67.57141, 67.6119, 67.65206, 67.69189, 67.73138, 
    67.77054, 67.80936, 67.84784, 67.88599, 67.92378, 67.96124, 67.99834, 
    68.03511, 68.07152, 68.10758, 68.14329, 68.17864, 68.21364, 68.24828, 
    68.28255, 68.31647, 68.35002, 68.38321, 68.41603, 68.44848, 68.48056, 
    68.51227, 68.5436, 68.57456, 68.60515, 68.63535, 68.66518, 68.69462, 
    68.72367, 68.75234, 68.78063, 68.80853, 68.83604, 68.86315, 68.88988, 
    68.9162, 68.94213, 68.96767, 68.99281, 69.01754, 69.04187, 69.0658, 
    69.08932, 69.11245, 69.13516, 69.15746, 69.17935, 69.20084, 69.2219, 
    69.24255, 69.26279, 69.28262, 69.30202, 69.32101, 69.33958, 69.35772, 
    69.37543, 69.39274, 69.40961, 69.42606, 69.44208, 69.45767, 69.47284, 
    69.48757, 69.50188, 69.51575, 69.52919, 69.5422, 69.55477, 69.5669, 
    69.57861, 69.58987, 69.6007, 69.61109, 69.62105, 69.63055, 69.63963, 
    69.64826, 69.65646, 69.6642, 69.67151, 69.67838, 69.6848, 69.69077, 
    69.69631, 69.7014, 69.70605, 69.71024, 69.714, 69.71732, 69.72018, 
    69.7226, 69.72457, 69.7261, 69.72717, 69.72781, 69.728, 69.72774, 
    69.72704, 69.72588, 69.72429, 69.72224, 69.71976, 69.71682, 69.71344, 
    69.70961, 69.70534, 69.70062, 69.69547, 69.68986, 69.68381, 69.67732, 
    69.67039, 69.66301, 69.65519, 69.64693, 69.63822, 69.62908, 69.6195, 
    69.60948, 69.59902, 69.58812, 69.57678, 69.56502, 69.55281, 69.54017, 
    69.52709, 69.51358, 69.49964, 69.48527, 69.47047, 69.45523, 69.43958, 
    69.42348, 69.40697, 69.39003, 69.37267, 69.35487, 69.33666, 69.31803, 
    69.29898, 69.27951, 69.25962, 69.23932, 69.2186, 69.19746, 69.17592, 
    69.15396, 69.13159, 69.10882, 69.08563, 69.06204, 69.03805, 69.01366, 
    68.98885, 68.96365, 68.93806, 68.91206, 68.88567, 68.85889, 68.83171, 
    68.80414, 68.77618, 68.74783, 68.7191, 68.68999, 68.66048, 68.6306, 
    68.60033, 68.56969, 68.53867, 68.50728, 68.47551, 68.44337, 68.41086, 
    68.37798, 68.34474, 68.31113, 68.27715, 68.24282, 68.20812, 68.17307, 
    68.13766, 68.1019, 68.06578, 68.02932, 67.9925, 67.95534, 67.91782, 
    67.87997, 67.84177, 67.80324, 67.76437, 67.72516, 67.68561, 67.64573, 
    67.60552, 67.56498, 67.52411, 67.48292, 67.44141, 67.39957, 67.35741, 
    67.31493, 67.27213, 67.22902, 67.1856, 67.14187, 67.09782, 67.05347, 
    67.00882, 66.96386, 66.91859, 66.87303, 66.82717, 66.78101, 66.73456, 
    66.68781, 66.64078, 66.59345, 66.54584, 66.49794, 66.44976, 66.40129, 
    66.35255, 66.30352, 66.25422, 66.20464, 66.15479, 66.10467, 66.05428, 
    66.00362, 65.95269, 65.9015, 65.85004, 65.79833, 65.74635, 65.69412, 
    65.64163, 65.58889, 65.5359, 65.48265, 65.42915, 65.37541, 65.32142, 
    65.26719, 65.21271, 65.15799, 65.10303, 65.04784, 64.99241, 64.93674, 
    64.88084, 64.82471, 64.76836, 64.71177, 64.65495, 64.59792, 64.54066, 
    64.48317, 64.42547, 64.36755, 64.3094, 64.25105, 64.19247, 64.1337, 
    64.0747, 64.0155,
  57.86238, 57.93576, 58.00904, 58.08222, 58.15528, 58.22824, 58.3011, 
    58.37384, 58.44647, 58.519, 58.59141, 58.66371, 58.73589, 58.80796, 
    58.87992, 58.95176, 59.02349, 59.09509, 59.16658, 59.23795, 59.3092, 
    59.38033, 59.45133, 59.52221, 59.59297, 59.6636, 59.73411, 59.80449, 
    59.87474, 59.94487, 60.01486, 60.08473, 60.15446, 60.22406, 60.29353, 
    60.36286, 60.43205, 60.50111, 60.57003, 60.63882, 60.70746, 60.77596, 
    60.84432, 60.91254, 60.98061, 61.04854, 61.11632, 61.18396, 61.25144, 
    61.31878, 61.38596, 61.453, 61.51988, 61.58661, 61.65318, 61.71959, 
    61.78585, 61.85195, 61.91789, 61.98367, 62.04928, 62.11473, 62.18002, 
    62.24514, 62.3101, 62.37488, 62.4395, 62.50394, 62.56822, 62.63232, 
    62.69624, 62.75999, 62.82356, 62.88696, 62.95017, 63.0132, 63.07605, 
    63.13871, 63.20119, 63.26348, 63.32559, 63.3875, 63.44923, 63.51076, 
    63.5721, 63.63324, 63.69419, 63.75494, 63.81549, 63.87584, 63.93599, 
    63.99593, 64.05567, 64.1152, 64.17452, 64.23363, 64.29254, 64.35123, 
    64.40971, 64.46796, 64.52601, 64.58383, 64.64144, 64.69882, 64.75598, 
    64.81291, 64.86962, 64.9261, 64.98235, 65.03837, 65.09415, 65.1497, 
    65.20502, 65.26009, 65.31493, 65.36953, 65.42388, 65.47799, 65.53185, 
    65.58547, 65.63883, 65.69195, 65.74481, 65.79742, 65.84977, 65.90186, 
    65.95369, 66.00526, 66.05657, 66.10761, 66.15839, 66.20889, 66.25913, 
    66.3091, 66.35879, 66.4082, 66.45734, 66.5062, 66.55478, 66.60307, 
    66.65108, 66.69881, 66.74625, 66.7934, 66.84025, 66.88681, 66.93307, 
    66.97904, 67.02471, 67.07008, 67.11515, 67.15991, 67.20437, 67.24851, 
    67.29235, 67.33588, 67.37909, 67.42198, 67.46456, 67.50682, 67.54876, 
    67.59037, 67.63166, 67.67263, 67.71326, 67.75357, 67.79354, 67.83318, 
    67.87248, 67.91145, 67.95007, 67.98836, 68.0263, 68.0639, 68.10114, 
    68.13805, 68.1746, 68.2108, 68.24664, 68.28214, 68.31726, 68.35204, 
    68.38644, 68.42049, 68.45418, 68.4875, 68.52045, 68.55303, 68.58524, 
    68.61707, 68.64854, 68.67962, 68.71033, 68.74065, 68.77059, 68.80016, 
    68.82933, 68.85812, 68.88652, 68.91454, 68.94215, 68.96938, 68.99622, 
    69.02266, 69.0487, 69.07434, 69.09958, 69.12442, 69.14886, 69.17289, 
    69.19651, 69.21973, 69.24254, 69.26494, 69.28693, 69.30849, 69.32966, 
    69.3504, 69.37073, 69.39063, 69.41013, 69.42919, 69.44784, 69.46606, 
    69.48386, 69.50124, 69.51818, 69.53471, 69.5508, 69.56646, 69.58169, 
    69.59649, 69.61086, 69.62479, 69.63829, 69.65136, 69.66399, 69.67618, 
    69.68793, 69.69925, 69.71013, 69.72057, 69.73056, 69.74011, 69.74923, 
    69.7579, 69.76613, 69.77391, 69.78125, 69.78815, 69.7946, 69.80061, 
    69.80617, 69.81128, 69.81595, 69.82017, 69.82394, 69.82726, 69.83014, 
    69.83257, 69.83456, 69.83609, 69.83717, 69.83781, 69.838, 69.83774, 
    69.83703, 69.83588, 69.83427, 69.83221, 69.82972, 69.82677, 69.82337, 
    69.81953, 69.81524, 69.8105, 69.80531, 69.79968, 69.79361, 69.78709, 
    69.78012, 69.77271, 69.76485, 69.75656, 69.74782, 69.73863, 69.729, 
    69.71894, 69.70844, 69.69749, 69.6861, 69.67428, 69.66202, 69.64931, 
    69.63618, 69.62261, 69.60861, 69.59418, 69.57931, 69.56401, 69.54828, 
    69.53212, 69.51553, 69.49851, 69.48107, 69.4632, 69.44492, 69.4262, 
    69.40707, 69.38751, 69.36754, 69.34715, 69.32634, 69.30511, 69.28348, 
    69.26142, 69.23896, 69.21609, 69.1928, 69.16911, 69.14502, 69.12052, 
    69.09562, 69.07031, 69.04461, 69.0185, 68.992, 68.9651, 68.93781, 
    68.91013, 68.88206, 68.85359, 68.82475, 68.7955, 68.76588, 68.73588, 
    68.70549, 68.67473, 68.64359, 68.61206, 68.58017, 68.5479, 68.51526, 
    68.48225, 68.44888, 68.41513, 68.38103, 68.34656, 68.31173, 68.27654, 
    68.241, 68.20509, 68.16884, 68.13223, 68.09528, 68.05797, 68.02032, 
    67.98232, 67.94398, 67.9053, 67.86629, 67.82693, 67.78724, 67.74722, 
    67.70686, 67.66617, 67.62515, 67.58381, 67.54214, 67.50016, 67.45785, 
    67.41522, 67.37228, 67.32901, 67.28544, 67.24155, 67.19736, 67.15285, 
    67.10804, 67.06293, 67.01751, 66.97179, 66.92578, 66.87946, 66.83286, 
    66.78596, 66.73876, 66.69128, 66.64351, 66.59545, 66.54711, 66.49849, 
    66.44958, 66.40041, 66.35094, 66.30121, 66.25121, 66.20092, 66.15038, 
    66.09956, 66.04847, 65.99712, 65.94551, 65.89364, 65.8415, 65.78911, 
    65.73647, 65.68356, 65.63041, 65.577, 65.52335, 65.46945, 65.4153, 
    65.36091, 65.30627, 65.2514, 65.19629, 65.14094, 65.08535, 65.02953, 
    64.97347, 64.91718, 64.86066, 64.80392, 64.74696, 64.68976, 64.63234, 
    64.5747, 64.51685, 64.45876, 64.40047, 64.34196, 64.28323, 64.2243, 
    64.16515, 64.1058,
  57.94014, 58.01364, 58.08703, 58.16032, 58.2335, 58.30657, 58.37954, 
    58.45239, 58.52514, 58.59778, 58.6703, 58.74272, 58.81502, 58.88721, 
    58.95928, 59.03124, 59.10308, 59.17481, 59.24641, 59.31791, 59.38927, 
    59.46052, 59.53165, 59.60265, 59.67353, 59.74429, 59.81492, 59.88542, 
    59.9558, 60.02605, 60.09617, 60.16616, 60.23602, 60.30574, 60.37534, 
    60.4448, 60.51412, 60.58331, 60.65236, 60.72128, 60.79005, 60.85868, 
    60.92717, 60.99552, 61.06373, 61.13179, 61.1997, 61.26748, 61.33509, 
    61.40257, 61.46989, 61.53706, 61.60408, 61.67094, 61.73765, 61.8042, 
    61.8706, 61.93684, 62.00291, 62.06883, 62.13459, 62.20018, 62.26561, 
    62.33088, 62.39597, 62.4609, 62.52566, 62.59025, 62.65467, 62.71891, 
    62.78298, 62.84687, 62.91059, 62.97413, 63.03749, 63.10067, 63.16367, 
    63.22648, 63.2891, 63.35155, 63.4138, 63.47586, 63.53774, 63.59942, 
    63.66091, 63.72221, 63.7833, 63.8442, 63.90491, 63.96541, 64.02571, 
    64.08581, 64.1457, 64.20538, 64.26486, 64.32413, 64.38319, 64.44203, 
    64.50066, 64.55907, 64.61727, 64.67525, 64.73302, 64.79055, 64.84787, 
    64.90496, 64.96182, 65.01846, 65.07487, 65.13104, 65.18699, 65.2427, 
    65.29816, 65.3534, 65.4084, 65.46315, 65.51766, 65.57193, 65.62595, 
    65.67973, 65.73325, 65.78652, 65.83955, 65.89231, 65.94482, 65.99707, 
    66.04906, 66.10079, 66.15226, 66.20346, 66.25439, 66.30506, 66.35545, 
    66.40558, 66.45543, 66.505, 66.5543, 66.60332, 66.65205, 66.70051, 
    66.74868, 66.79656, 66.84415, 66.89146, 66.93847, 66.98519, 67.03161, 
    67.07774, 67.12356, 67.16908, 67.2143, 67.25922, 67.30383, 67.34813, 
    67.39212, 67.4358, 67.47916, 67.52222, 67.56494, 67.60735, 67.64944, 
    67.69121, 67.73265, 67.77376, 67.81454, 67.855, 67.89512, 67.93491, 
    67.97435, 68.01347, 68.05223, 68.09066, 68.12875, 68.16649, 68.20388, 
    68.24092, 68.27761, 68.31395, 68.34993, 68.38556, 68.42083, 68.45573, 
    68.49028, 68.52447, 68.55828, 68.59174, 68.62482, 68.65752, 68.68987, 
    68.72182, 68.75341, 68.78462, 68.81545, 68.8459, 68.87597, 68.90565, 
    68.93495, 68.96386, 68.99238, 69.02051, 69.04824, 69.07558, 69.10253, 
    69.12908, 69.15523, 69.18098, 69.20633, 69.23127, 69.25581, 69.27995, 
    69.30367, 69.32699, 69.34989, 69.37239, 69.39447, 69.41614, 69.43739, 
    69.45822, 69.47864, 69.49863, 69.5182, 69.53736, 69.55608, 69.57439, 
    69.59227, 69.60972, 69.62674, 69.64333, 69.6595, 69.67523, 69.69053, 
    69.7054, 69.71983, 69.73383, 69.74738, 69.76051, 69.77319, 69.78544, 
    69.79725, 69.80862, 69.81954, 69.83002, 69.84007, 69.84967, 69.85883, 
    69.86753, 69.8758, 69.88362, 69.89099, 69.89792, 69.9044, 69.91044, 
    69.91602, 69.92116, 69.92584, 69.93008, 69.93388, 69.93722, 69.94011, 
    69.94255, 69.94453, 69.94608, 69.94717, 69.94781, 69.948, 69.94774, 
    69.94703, 69.94586, 69.94425, 69.94219, 69.93968, 69.93671, 69.9333, 
    69.92944, 69.92513, 69.92037, 69.91517, 69.90951, 69.9034, 69.89686, 
    69.88985, 69.88242, 69.87452, 69.86619, 69.85741, 69.84818, 69.83851, 
    69.8284, 69.81784, 69.80685, 69.79541, 69.78353, 69.77122, 69.75846, 
    69.74527, 69.73164, 69.71758, 69.70307, 69.68814, 69.67277, 69.65697, 
    69.64074, 69.62408, 69.60699, 69.58947, 69.57153, 69.55315, 69.53436, 
    69.51514, 69.4955, 69.47543, 69.45496, 69.43405, 69.41273, 69.39101, 
    69.36886, 69.3463, 69.32333, 69.29994, 69.27615, 69.25195, 69.22736, 
    69.20235, 69.17693, 69.15112, 69.12491, 69.09829, 69.07128, 69.04388, 
    69.01608, 68.98789, 68.95931, 68.93034, 68.90099, 68.87124, 68.84111, 
    68.8106, 68.77971, 68.74844, 68.7168, 68.68477, 68.65237, 68.61961, 
    68.58646, 68.55296, 68.51908, 68.48484, 68.45024, 68.41528, 68.37995, 
    68.34426, 68.30823, 68.27183, 68.23508, 68.19798, 68.16054, 68.12275, 
    68.08461, 68.04612, 68.0073, 67.96813, 67.92863, 67.88879, 67.84862, 
    67.80811, 67.76728, 67.72611, 67.68462, 67.64281, 67.60067, 67.5582, 
    67.51543, 67.47233, 67.42892, 67.38519, 67.34115, 67.2968, 67.25214, 
    67.20718, 67.1619, 67.11633, 67.07046, 67.02428, 66.97781, 66.93105, 
    66.884, 66.83665, 66.789, 66.74107, 66.69286, 66.64436, 66.59558, 
    66.54652, 66.49718, 66.44756, 66.39767, 66.3475, 66.29707, 66.24635, 
    66.19538, 66.14413, 66.09263, 66.04086, 65.98882, 65.93653, 65.88398, 
    65.83118, 65.77811, 65.7248, 65.67123, 65.61742, 65.56336, 65.50906, 
    65.45451, 65.39971, 65.34468, 65.28941, 65.2339, 65.17815, 65.12218, 
    65.06596, 65.00952, 64.95284, 64.89594, 64.83882, 64.78146, 64.72389, 
    64.6661, 64.60809, 64.54985, 64.4914, 64.43273, 64.37386, 64.31477, 
    64.25546, 64.19595,
  58.01775, 58.09135, 58.16485, 58.23825, 58.31154, 58.38473, 58.45781, 
    58.53078, 58.60364, 58.67639, 58.74903, 58.82156, 58.89398, 58.96628, 
    59.03848, 59.11055, 59.18251, 59.25436, 59.32608, 59.39769, 59.46918, 
    59.54055, 59.6118, 59.68292, 59.75393, 59.82481, 59.89556, 59.96619, 
    60.03669, 60.10706, 60.17731, 60.24743, 60.31741, 60.38726, 60.45699, 
    60.52657, 60.59603, 60.66534, 60.73453, 60.80357, 60.87247, 60.94124, 
    61.00986, 61.07834, 61.14668, 61.21488, 61.28292, 61.35083, 61.41858, 
    61.48619, 61.55365, 61.62096, 61.68811, 61.75511, 61.82196, 61.88865, 
    61.95518, 62.02156, 62.08778, 62.15384, 62.21974, 62.28547, 62.35104, 
    62.41645, 62.48169, 62.54676, 62.61166, 62.6764, 62.74096, 62.80535, 
    62.86956, 62.9336, 62.99747, 63.06115, 63.12466, 63.18798, 63.25113, 
    63.31409, 63.37687, 63.43946, 63.50186, 63.56408, 63.6261, 63.68793, 
    63.74957, 63.81102, 63.87227, 63.93332, 63.99417, 64.05483, 64.11528, 
    64.17553, 64.23558, 64.29542, 64.35505, 64.41447, 64.47369, 64.53268, 
    64.59147, 64.65005, 64.7084, 64.76653, 64.82446, 64.88215, 64.93962, 
    64.99687, 65.05389, 65.11069, 65.16725, 65.22359, 65.27969, 65.33556, 
    65.39118, 65.44658, 65.50173, 65.55665, 65.61132, 65.66575, 65.71992, 
    65.77386, 65.82755, 65.88097, 65.93416, 65.98708, 66.03975, 66.09216, 
    66.14431, 66.19621, 66.24783, 66.29919, 66.35029, 66.40112, 66.45167, 
    66.50195, 66.55196, 66.60169, 66.65115, 66.70033, 66.74922, 66.79784, 
    66.84616, 66.8942, 66.94196, 66.98942, 67.03659, 67.08347, 67.13004, 
    67.17632, 67.22231, 67.26799, 67.31337, 67.35844, 67.40321, 67.44766, 
    67.49181, 67.53564, 67.57915, 67.62236, 67.66524, 67.7078, 67.75005, 
    67.79196, 67.83355, 67.87482, 67.91575, 67.95635, 67.99662, 68.03655, 
    68.07615, 68.1154, 68.15432, 68.19289, 68.23112, 68.269, 68.30654, 
    68.34373, 68.38056, 68.41704, 68.45316, 68.48893, 68.52433, 68.55938, 
    68.59406, 68.62838, 68.66233, 68.69592, 68.72913, 68.76197, 68.79443, 
    68.82653, 68.85825, 68.88958, 68.92053, 68.95111, 68.9813, 69.01111, 
    69.04052, 69.06955, 69.09819, 69.12643, 69.15429, 69.18174, 69.2088, 
    69.23547, 69.26173, 69.28758, 69.31304, 69.33809, 69.36273, 69.38697, 
    69.4108, 69.43422, 69.45722, 69.47981, 69.50199, 69.52375, 69.5451, 
    69.56602, 69.58652, 69.60661, 69.62627, 69.64551, 69.66431, 69.6827, 
    69.70065, 69.71819, 69.73528, 69.75195, 69.76819, 69.78399, 69.79935, 
    69.81429, 69.82879, 69.84285, 69.85647, 69.86965, 69.88239, 69.8947, 
    69.90656, 69.91798, 69.92896, 69.93948, 69.94958, 69.95921, 69.96841, 
    69.97717, 69.98547, 69.99332, 70.00073, 70.00769, 70.0142, 70.02026, 
    70.02587, 70.03104, 70.03574, 70.04, 70.04381, 70.04716, 70.05007, 
    70.05252, 70.05452, 70.05607, 70.05717, 70.05781, 70.058, 70.05774, 
    70.05702, 70.05585, 70.05424, 70.05216, 70.04964, 70.04666, 70.04324, 
    70.03936, 70.03503, 70.03025, 70.02502, 70.01933, 70.0132, 70.00662, 
    69.99959, 69.99211, 69.98418, 69.97581, 69.96699, 69.95772, 69.94801, 
    69.93785, 69.92725, 69.9162, 69.90471, 69.89278, 69.88041, 69.8676, 
    69.85434, 69.84065, 69.82652, 69.81196, 69.79695, 69.78152, 69.76565, 
    69.74934, 69.7326, 69.71544, 69.69785, 69.67982, 69.66137, 69.64249, 
    69.62318, 69.60346, 69.58331, 69.56274, 69.54175, 69.52034, 69.49851, 
    69.47626, 69.45361, 69.43054, 69.40706, 69.38316, 69.35886, 69.33415, 
    69.30904, 69.28352, 69.2576, 69.23127, 69.20455, 69.17743, 69.14991, 
    69.12199, 69.09368, 69.06499, 69.0359, 69.00642, 68.97655, 68.9463, 
    68.91566, 68.88465, 68.85325, 68.82148, 68.78932, 68.7568, 68.7239, 
    68.69063, 68.65698, 68.62298, 68.5886, 68.55386, 68.51875, 68.48329, 
    68.44747, 68.41129, 68.37476, 68.33787, 68.30063, 68.26304, 68.2251, 
    68.18681, 68.14819, 68.10921, 68.06991, 68.03026, 67.99027, 67.94995, 
    67.90929, 67.86831, 67.827, 67.78535, 67.74339, 67.70109, 67.65848, 
    67.61555, 67.5723, 67.52872, 67.48484, 67.44065, 67.39614, 67.35133, 
    67.30621, 67.26078, 67.21506, 67.16902, 67.1227, 67.07607, 67.02914, 
    66.98193, 66.93443, 66.88663, 66.83854, 66.79017, 66.74151, 66.69257, 
    66.64335, 66.59385, 66.54407, 66.49402, 66.44369, 66.39309, 66.34222, 
    66.29108, 66.23969, 66.18801, 66.13608, 66.08389, 66.03143, 65.97873, 
    65.92576, 65.87254, 65.81907, 65.76534, 65.71137, 65.65715, 65.60268, 
    65.54798, 65.49303, 65.43784, 65.3824, 65.32674, 65.27083, 65.21469, 
    65.15832, 65.10172, 65.04488, 64.98783, 64.93054, 64.87304, 64.81531, 
    64.75735, 64.69918, 64.64079, 64.58218, 64.52337, 64.46433, 64.40509, 
    64.34563, 64.28596,
  58.09518, 58.16889, 58.2425, 58.31601, 58.38942, 58.46272, 58.5359, 
    58.60899, 58.68196, 58.75483, 58.82759, 58.90023, 58.97277, 59.04519, 
    59.1175, 59.18969, 59.26177, 59.33373, 59.40558, 59.47731, 59.54892, 
    59.62041, 59.69178, 59.76302, 59.83415, 59.90515, 59.97603, 60.04678, 
    60.11741, 60.18791, 60.25828, 60.32853, 60.39864, 60.46862, 60.53847, 
    60.60818, 60.67776, 60.74721, 60.81652, 60.8857, 60.95473, 61.02363, 
    61.09238, 61.161, 61.22947, 61.2978, 61.36598, 61.43402, 61.50191, 
    61.56965, 61.63725, 61.70469, 61.77198, 61.83912, 61.90611, 61.97294, 
    62.03961, 62.10613, 62.17249, 62.23869, 62.30473, 62.3706, 62.43631, 
    62.50186, 62.56725, 62.63246, 62.69751, 62.76238, 62.82709, 62.89162, 
    62.95599, 63.02017, 63.08418, 63.14801, 63.21167, 63.27514, 63.33844, 
    63.40155, 63.46447, 63.52721, 63.58977, 63.65213, 63.71431, 63.77629, 
    63.83808, 63.89968, 63.96108, 64.02229, 64.0833, 64.1441, 64.20471, 
    64.26511, 64.32532, 64.38531, 64.4451, 64.50468, 64.56404, 64.6232, 
    64.68214, 64.74087, 64.79939, 64.85767, 64.91575, 64.9736, 65.03123, 
    65.08865, 65.14582, 65.20277, 65.2595, 65.31599, 65.37225, 65.42828, 
    65.48407, 65.53963, 65.59494, 65.65002, 65.70484, 65.75943, 65.81377, 
    65.86787, 65.92171, 65.9753, 66.02865, 66.08173, 66.13456, 66.18713, 
    66.23945, 66.2915, 66.34328, 66.39481, 66.44606, 66.49705, 66.54777, 
    66.59821, 66.64838, 66.69827, 66.74789, 66.79723, 66.84628, 66.89506, 
    66.94354, 66.99174, 67.03966, 67.08728, 67.13461, 67.18164, 67.22838, 
    67.27482, 67.32096, 67.3668, 67.41233, 67.45756, 67.50248, 67.5471, 
    67.59139, 67.63538, 67.67905, 67.72241, 67.76545, 67.80817, 67.85056, 
    67.89263, 67.93437, 67.97578, 68.01687, 68.05762, 68.09804, 68.13812, 
    68.17786, 68.21727, 68.25634, 68.29506, 68.33343, 68.37146, 68.40913, 
    68.44646, 68.48344, 68.52006, 68.55633, 68.59223, 68.62778, 68.66296, 
    68.69778, 68.73223, 68.76632, 68.80003, 68.83338, 68.86636, 68.89896, 
    68.93118, 68.96302, 68.99448, 69.02557, 69.05627, 69.08659, 69.11652, 
    69.14605, 69.1752, 69.20396, 69.23232, 69.26029, 69.28786, 69.31504, 
    69.34181, 69.36819, 69.39415, 69.41972, 69.44488, 69.46963, 69.49397, 
    69.5179, 69.54142, 69.56452, 69.58721, 69.60949, 69.63135, 69.65278, 
    69.6738, 69.69439, 69.71456, 69.73431, 69.75363, 69.77253, 69.79099, 
    69.80903, 69.82664, 69.84381, 69.86055, 69.87686, 69.89274, 69.90817, 
    69.92317, 69.93774, 69.95186, 69.96555, 69.97878, 69.99158, 70.00394, 
    70.01586, 70.02734, 70.03836, 70.04894, 70.05907, 70.06876, 70.078, 
    70.08679, 70.09513, 70.10303, 70.11047, 70.11745, 70.124, 70.13009, 
    70.13573, 70.14091, 70.14564, 70.14992, 70.15374, 70.15711, 70.16003, 
    70.1625, 70.16451, 70.16606, 70.16716, 70.16781, 70.168, 70.16773, 
    70.16702, 70.16585, 70.16422, 70.16214, 70.1596, 70.15661, 70.15317, 
    70.14927, 70.14492, 70.14012, 70.13486, 70.12915, 70.12299, 70.11638, 
    70.10932, 70.10181, 70.09384, 70.08543, 70.07657, 70.06726, 70.0575, 
    70.04729, 70.03664, 70.02555, 70.01401, 70.00202, 69.98959, 69.97672, 
    69.96341, 69.94965, 69.93546, 69.92083, 69.90576, 69.89025, 69.87431, 
    69.85793, 69.84113, 69.82388, 69.80621, 69.7881, 69.76957, 69.7506, 
    69.73122, 69.7114, 69.69116, 69.6705, 69.64942, 69.62791, 69.606, 
    69.58365, 69.5609, 69.53773, 69.51414, 69.49014, 69.46574, 69.44093, 
    69.4157, 69.39008, 69.36404, 69.3376, 69.31077, 69.28353, 69.25589, 
    69.22786, 69.19943, 69.17062, 69.1414, 69.1118, 69.08182, 69.05144, 
    69.02068, 68.98953, 68.95801, 68.92611, 68.89382, 68.86117, 68.82813, 
    68.79473, 68.76096, 68.72681, 68.6923, 68.65742, 68.62218, 68.58657, 
    68.55061, 68.51429, 68.47762, 68.44058, 68.4032, 68.36546, 68.32738, 
    68.28896, 68.25018, 68.21106, 68.1716, 68.13181, 68.09167, 68.0512, 
    68.01039, 67.96925, 67.92779, 67.88599, 67.84387, 67.80143, 67.75866, 
    67.71558, 67.67217, 67.62845, 67.58441, 67.54006, 67.4954, 67.45042, 
    67.40515, 67.35957, 67.31368, 67.26749, 67.22101, 67.17422, 67.12714, 
    67.07977, 67.0321, 66.98414, 66.93589, 66.88736, 66.83855, 66.78944, 
    66.74006, 66.6904, 66.64046, 66.59025, 66.53976, 66.489, 66.43797, 
    66.38667, 66.33511, 66.28328, 66.23119, 66.17883, 66.12622, 66.07335, 
    66.02023, 65.96684, 65.91321, 65.85933, 65.80519, 65.75082, 65.69619, 
    65.64132, 65.5862, 65.53085, 65.47527, 65.41943, 65.36337, 65.30708, 
    65.25054, 65.19378, 65.1368, 65.07957, 65.02213, 64.96447, 64.90658, 
    64.84847, 64.79015, 64.7316, 64.67284, 64.61385, 64.55466, 64.49526, 
    64.43565, 64.37583,
  58.17243, 58.24626, 58.31998, 58.3936, 58.46712, 58.54053, 58.61383, 
    58.68703, 58.76012, 58.8331, 58.90597, 58.97873, 59.05138, 59.12392, 
    59.19635, 59.26866, 59.34086, 59.41294, 59.48491, 59.55675, 59.62848, 
    59.7001, 59.77158, 59.84296, 59.9142, 59.98533, 60.05633, 60.12721, 
    60.19796, 60.26859, 60.33908, 60.40945, 60.47969, 60.5498, 60.61978, 
    60.68962, 60.75933, 60.82891, 60.89835, 60.96766, 61.03682, 61.10585, 
    61.17474, 61.24348, 61.31209, 61.38055, 61.44887, 61.51704, 61.58507, 
    61.65295, 61.72068, 61.78826, 61.85569, 61.92297, 61.99009, 62.05706, 
    62.12387, 62.19053, 62.25703, 62.32337, 62.38955, 62.45557, 62.52142, 
    62.58711, 62.65264, 62.718, 62.78319, 62.84821, 62.91306, 62.97775, 
    63.04225, 63.10659, 63.17074, 63.23472, 63.29852, 63.36215, 63.42559, 
    63.48885, 63.55192, 63.61481, 63.67752, 63.74004, 63.80236, 63.8645, 
    63.92644, 63.98819, 64.04974, 64.11111, 64.17226, 64.23323, 64.29399, 
    64.35455, 64.4149, 64.47505, 64.535, 64.59473, 64.65426, 64.71357, 
    64.77267, 64.83156, 64.89023, 64.94868, 65.00691, 65.06492, 65.12271, 
    65.18027, 65.23762, 65.29473, 65.35161, 65.40826, 65.46468, 65.52087, 
    65.57682, 65.63254, 65.68801, 65.74325, 65.79824, 65.85299, 65.90749, 
    65.96175, 66.01575, 66.0695, 66.12301, 66.17625, 66.22925, 66.28198, 
    66.33446, 66.38667, 66.43862, 66.4903, 66.54172, 66.59287, 66.64375, 
    66.69435, 66.74468, 66.79474, 66.84452, 66.89402, 66.94324, 66.99216, 
    67.04082, 67.08918, 67.13725, 67.18503, 67.23252, 67.27972, 67.32661, 
    67.37321, 67.41951, 67.46551, 67.5112, 67.55659, 67.60167, 67.64644, 
    67.6909, 67.73504, 67.77887, 67.82238, 67.86557, 67.90844, 67.95099, 
    67.99321, 68.03511, 68.07668, 68.11791, 68.15881, 68.19939, 68.23962, 
    68.27951, 68.31906, 68.35828, 68.39714, 68.43567, 68.47384, 68.51167, 
    68.54913, 68.58625, 68.62302, 68.65942, 68.69547, 68.73116, 68.76648, 
    68.80144, 68.83603, 68.87025, 68.90411, 68.93758, 68.97069, 69.00343, 
    69.03577, 69.06775, 69.09934, 69.13055, 69.16138, 69.19183, 69.22188, 
    69.25153, 69.28081, 69.30968, 69.33817, 69.36626, 69.39394, 69.42123, 
    69.44812, 69.47461, 69.50069, 69.52636, 69.55163, 69.57648, 69.60094, 
    69.62497, 69.64859, 69.6718, 69.69459, 69.71696, 69.73891, 69.76044, 
    69.78155, 69.80224, 69.82249, 69.84233, 69.86174, 69.88072, 69.89927, 
    69.91739, 69.93507, 69.95232, 69.96914, 69.98553, 70.00147, 70.01698, 
    70.03204, 70.04668, 70.06086, 70.07461, 70.08791, 70.10077, 70.11319, 
    70.12516, 70.13668, 70.14776, 70.15839, 70.16857, 70.1783, 70.18758, 
    70.19641, 70.2048, 70.21272, 70.2202, 70.22723, 70.2338, 70.23991, 
    70.24557, 70.25078, 70.25554, 70.25983, 70.26368, 70.26707, 70.27, 
    70.27247, 70.27449, 70.27605, 70.27716, 70.27781, 70.278, 70.27773, 
    70.27702, 70.27583, 70.2742, 70.27211, 70.26956, 70.26656, 70.2631, 
    70.25919, 70.25481, 70.24998, 70.24471, 70.23898, 70.23278, 70.22614, 
    70.21905, 70.21149, 70.2035, 70.19505, 70.18614, 70.17679, 70.16698, 
    70.15674, 70.14603, 70.13489, 70.12329, 70.11125, 70.09877, 70.08584, 
    70.07246, 70.05865, 70.04439, 70.02969, 70.01455, 69.99898, 69.98296, 
    69.96651, 69.94962, 69.9323, 69.91455, 69.89636, 69.87775, 69.8587, 
    69.83923, 69.81932, 69.799, 69.77824, 69.75706, 69.73547, 69.71345, 
    69.69101, 69.66815, 69.64488, 69.62119, 69.59709, 69.57259, 69.54766, 
    69.52233, 69.49659, 69.47044, 69.44389, 69.41695, 69.3896, 69.36184, 
    69.33369, 69.30515, 69.27621, 69.24687, 69.21715, 69.18703, 69.15653, 
    69.12564, 69.09438, 69.06272, 69.03069, 68.99827, 68.96548, 68.93231, 
    68.89877, 68.86486, 68.83058, 68.79593, 68.76092, 68.72553, 68.68979, 
    68.65369, 68.61723, 68.58041, 68.54323, 68.50571, 68.46783, 68.4296, 
    68.39102, 68.3521, 68.31283, 68.27322, 68.23328, 68.19299, 68.15237, 
    68.11141, 68.07012, 68.0285, 67.98656, 67.94428, 67.90168, 67.85876, 
    67.81551, 67.77196, 67.72807, 67.68388, 67.63937, 67.59456, 67.54943, 
    67.50399, 67.45825, 67.41221, 67.36586, 67.31921, 67.27227, 67.22503, 
    67.17749, 67.12966, 67.08154, 67.03314, 66.98444, 66.93547, 66.88621, 
    66.83666, 66.78684, 66.73674, 66.68637, 66.63572, 66.58479, 66.53361, 
    66.48215, 66.43042, 66.37843, 66.32617, 66.27366, 66.22089, 66.16785, 
    66.11456, 66.06102, 66.00723, 65.95318, 65.89889, 65.84435, 65.78956, 
    65.73453, 65.67925, 65.62374, 65.56799, 65.512, 65.45578, 65.39932, 
    65.34263, 65.28571, 65.22856, 65.17119, 65.11359, 65.05576, 64.99771, 
    64.93945, 64.88096, 64.82226, 64.76334, 64.7042, 64.64485, 64.5853, 
    64.52553, 64.46555,
  58.24952, 58.32346, 58.39729, 58.47102, 58.54465, 58.61817, 58.69159, 
    58.7649, 58.8381, 58.9112, 58.98418, 59.05706, 59.12983, 59.20248, 
    59.27503, 59.34746, 59.41977, 59.49197, 59.56406, 59.63603, 59.70788, 
    59.77961, 59.85122, 59.92271, 59.99409, 60.06533, 60.13646, 60.20746, 
    60.27834, 60.34909, 60.41971, 60.49021, 60.56058, 60.63081, 60.70092, 
    60.77089, 60.84073, 60.91044, 60.98001, 61.04945, 61.11874, 61.1879, 
    61.25692, 61.32581, 61.39454, 61.46314, 61.53159, 61.5999, 61.66806, 
    61.73608, 61.80394, 61.87166, 61.93923, 62.00665, 62.07391, 62.14101, 
    62.20797, 62.27477, 62.34141, 62.40789, 62.47421, 62.54037, 62.60637, 
    62.6722, 62.73787, 62.80338, 62.86871, 62.93388, 62.99888, 63.06371, 
    63.12836, 63.19284, 63.25714, 63.32127, 63.38522, 63.44899, 63.51258, 
    63.57599, 63.63922, 63.70226, 63.76511, 63.82778, 63.89026, 63.95255, 
    64.01465, 64.07655, 64.13826, 64.19978, 64.26109, 64.3222, 64.38312, 
    64.44383, 64.50435, 64.56465, 64.62475, 64.68464, 64.74432, 64.80379, 
    64.86305, 64.9221, 64.98093, 65.03954, 65.09792, 65.1561, 65.21404, 
    65.27177, 65.32927, 65.38654, 65.44359, 65.5004, 65.55698, 65.61333, 
    65.66944, 65.72532, 65.78095, 65.83635, 65.8915, 65.94641, 66.00108, 
    66.0555, 66.10966, 66.16358, 66.21725, 66.27066, 66.32381, 66.37671, 
    66.42934, 66.48172, 66.53384, 66.58568, 66.63726, 66.68857, 66.73962, 
    66.79038, 66.84087, 66.89109, 66.94103, 66.99069, 67.04008, 67.08917, 
    67.13798, 67.1865, 67.23473, 67.28268, 67.33033, 67.37769, 67.42474, 
    67.4715, 67.51796, 67.56412, 67.60997, 67.65552, 67.70075, 67.74568, 
    67.7903, 67.8346, 67.87859, 67.92226, 67.9656, 68.00863, 68.05133, 
    68.09371, 68.13576, 68.17748, 68.21887, 68.25993, 68.30064, 68.34103, 
    68.38107, 68.42078, 68.46014, 68.49916, 68.53783, 68.57615, 68.61412, 
    68.65173, 68.689, 68.72591, 68.76246, 68.79865, 68.83447, 68.86993, 
    68.90503, 68.93977, 68.97412, 69.00811, 69.04173, 69.07497, 69.10783, 
    69.14032, 69.17242, 69.20415, 69.23549, 69.26645, 69.29701, 69.32719, 
    69.35698, 69.38638, 69.41537, 69.44398, 69.47218, 69.49999, 69.5274, 
    69.5544, 69.58099, 69.60719, 69.63297, 69.65835, 69.68332, 69.70787, 
    69.73201, 69.75574, 69.77905, 69.80193, 69.8244, 69.84645, 69.86808, 
    69.88928, 69.91006, 69.93041, 69.95033, 69.96983, 69.98889, 70.00752, 
    70.02573, 70.04349, 70.06082, 70.07771, 70.09417, 70.11019, 70.12577, 
    70.14091, 70.1556, 70.16985, 70.18366, 70.19703, 70.20995, 70.22242, 
    70.23444, 70.24603, 70.25715, 70.26783, 70.27805, 70.28783, 70.29716, 
    70.30603, 70.31445, 70.32242, 70.32993, 70.33698, 70.34358, 70.34973, 
    70.35542, 70.36066, 70.36543, 70.36975, 70.37361, 70.37701, 70.37996, 
    70.38245, 70.38448, 70.38604, 70.38715, 70.3878, 70.388, 70.38773, 
    70.38701, 70.38583, 70.38419, 70.38208, 70.37952, 70.3765, 70.37303, 
    70.36909, 70.36471, 70.35986, 70.35455, 70.34879, 70.34258, 70.3359, 
    70.32877, 70.32119, 70.31315, 70.30466, 70.29572, 70.28632, 70.27647, 
    70.26617, 70.25542, 70.24422, 70.23257, 70.22047, 70.20793, 70.19495, 
    70.18151, 70.16763, 70.15331, 70.13854, 70.12333, 70.10768, 70.0916, 
    70.07507, 70.05811, 70.04071, 70.02287, 70.00461, 69.98591, 69.96677, 
    69.94721, 69.92722, 69.9068, 69.88596, 69.86469, 69.84299, 69.82088, 
    69.79834, 69.77538, 69.75201, 69.72822, 69.70401, 69.6794, 69.65437, 
    69.62892, 69.60307, 69.57681, 69.55016, 69.52309, 69.49561, 69.46774, 
    69.43948, 69.41081, 69.38175, 69.35229, 69.32244, 69.29221, 69.26157, 
    69.23056, 69.19916, 69.16737, 69.13521, 69.10266, 69.06974, 69.03644, 
    69.00276, 68.96871, 68.9343, 68.89951, 68.86435, 68.82883, 68.79295, 
    68.7567, 68.72009, 68.68313, 68.64581, 68.60814, 68.57011, 68.53173, 
    68.49301, 68.45394, 68.41452, 68.37476, 68.33466, 68.29423, 68.25346, 
    68.21235, 68.17091, 68.12913, 68.08703, 68.0446, 68.00185, 67.95876, 
    67.91537, 67.87165, 67.82761, 67.78326, 67.73859, 67.69362, 67.64833, 
    67.60274, 67.55684, 67.51063, 67.46413, 67.41732, 67.37021, 67.32281, 
    67.27512, 67.22713, 67.17885, 67.13028, 67.08142, 67.03228, 66.98286, 
    66.93315, 66.88317, 66.83291, 66.78237, 66.73156, 66.68047, 66.62912, 
    66.5775, 66.5256, 66.47345, 66.42104, 66.36835, 66.31542, 66.26222, 
    66.20878, 66.15507, 66.10111, 66.04691, 65.99245, 65.93774, 65.8828, 
    65.82761, 65.77217, 65.71649, 65.66058, 65.60443, 65.54805, 65.49142, 
    65.43458, 65.37749, 65.32019, 65.26266, 65.2049, 65.14691, 65.08871, 
    65.03027, 64.97163, 64.91277, 64.85369, 64.7944, 64.73489, 64.67518, 
    64.61526, 64.55512,
  58.32643, 58.40048, 58.47442, 58.54827, 58.62201, 58.69564, 58.76917, 
    58.84259, 58.91591, 58.98912, 59.06223, 59.13522, 59.2081, 59.28087, 
    59.35353, 59.42608, 59.49851, 59.57084, 59.64304, 59.71513, 59.7871, 
    59.85895, 59.93069, 60.0023, 60.0738, 60.14517, 60.21642, 60.28754, 
    60.35855, 60.42942, 60.50017, 60.57079, 60.64129, 60.71165, 60.78189, 
    60.85199, 60.92196, 60.99179, 61.0615, 61.13107, 61.20049, 61.26979, 
    61.33894, 61.40795, 61.47683, 61.54556, 61.61414, 61.68259, 61.75089, 
    61.81903, 61.88704, 61.9549, 62.0226, 62.09015, 62.15755, 62.2248, 
    62.2919, 62.35884, 62.42562, 62.49224, 62.5587, 62.62501, 62.69115, 
    62.75713, 62.82294, 62.88859, 62.95407, 63.01938, 63.08453, 63.1495, 
    63.2143, 63.27893, 63.34338, 63.40766, 63.47176, 63.53568, 63.59942, 
    63.66298, 63.72636, 63.78955, 63.85255, 63.91537, 63.978, 64.04044, 
    64.1027, 64.16476, 64.22662, 64.28828, 64.34975, 64.41103, 64.4721, 
    64.53297, 64.59364, 64.6541, 64.71436, 64.7744, 64.83424, 64.89387, 
    64.95329, 65.01249, 65.07147, 65.13025, 65.1888, 65.24712, 65.30524, 
    65.36312, 65.42078, 65.47822, 65.53542, 65.59239, 65.64914, 65.70565, 
    65.76192, 65.81796, 65.87376, 65.92932, 65.98463, 66.03971, 66.09454, 
    66.14912, 66.20345, 66.25753, 66.31136, 66.36493, 66.41825, 66.47131, 
    66.52411, 66.57664, 66.62892, 66.68094, 66.73268, 66.78416, 66.83536, 
    66.88629, 66.93695, 66.98733, 67.03744, 67.08726, 67.1368, 67.18606, 
    67.23503, 67.28371, 67.33212, 67.38022, 67.42803, 67.47555, 67.52277, 
    67.56969, 67.61631, 67.66263, 67.70864, 67.75435, 67.79974, 67.84483, 
    67.8896, 67.93407, 67.97821, 68.02203, 68.06554, 68.10873, 68.15159, 
    68.19412, 68.23633, 68.2782, 68.31975, 68.36095, 68.40183, 68.44237, 
    68.48256, 68.52242, 68.56193, 68.6011, 68.63992, 68.67838, 68.7165, 
    68.75426, 68.79167, 68.82873, 68.86542, 68.90176, 68.93772, 68.97333, 
    69.00857, 69.04343, 69.07793, 69.11206, 69.14581, 69.17919, 69.2122, 
    69.24481, 69.27705, 69.30891, 69.34038, 69.37146, 69.40215, 69.43246, 
    69.46237, 69.49189, 69.52101, 69.54974, 69.57806, 69.60599, 69.63351, 
    69.66064, 69.68735, 69.71365, 69.73955, 69.76504, 69.79012, 69.81477, 
    69.83902, 69.86285, 69.88626, 69.90925, 69.93182, 69.95396, 69.97569, 
    69.99699, 70.01786, 70.0383, 70.05831, 70.0779, 70.09705, 70.11576, 
    70.13405, 70.15189, 70.1693, 70.18627, 70.2028, 70.21889, 70.23454, 
    70.24976, 70.26452, 70.27883, 70.29271, 70.30614, 70.31911, 70.33164, 
    70.34373, 70.35535, 70.36654, 70.37727, 70.38754, 70.39736, 70.40673, 
    70.41564, 70.4241, 70.43211, 70.43965, 70.44675, 70.45338, 70.45955, 
    70.46527, 70.47053, 70.47533, 70.47966, 70.48354, 70.48696, 70.48992, 
    70.49242, 70.49445, 70.49603, 70.49715, 70.4978, 70.498, 70.49773, 
    70.497, 70.49581, 70.49416, 70.49205, 70.48948, 70.48645, 70.48296, 
    70.479, 70.47459, 70.46973, 70.46439, 70.4586, 70.45235, 70.44566, 
    70.43849, 70.43087, 70.4228, 70.41427, 70.40528, 70.39584, 70.38595, 
    70.3756, 70.3648, 70.35355, 70.34184, 70.32969, 70.31709, 70.30404, 
    70.29054, 70.2766, 70.26221, 70.24738, 70.2321, 70.21638, 70.20022, 
    70.18362, 70.16658, 70.1491, 70.13118, 70.11283, 70.09405, 70.07483, 
    70.05518, 70.0351, 70.01459, 69.99364, 69.97228, 69.95049, 69.92828, 
    69.90564, 69.88258, 69.85911, 69.83521, 69.8109, 69.78617, 69.76103, 
    69.73548, 69.70952, 69.68315, 69.65637, 69.62919, 69.6016, 69.57361, 
    69.54522, 69.51643, 69.48725, 69.45766, 69.4277, 69.39732, 69.36657, 
    69.33543, 69.30389, 69.27198, 69.23968, 69.207, 69.17394, 69.1405, 
    69.10669, 69.0725, 69.03795, 69.00301, 68.96772, 68.93206, 68.89603, 
    68.85964, 68.82289, 68.78578, 68.74831, 68.71049, 68.67233, 68.6338, 
    68.59492, 68.5557, 68.51614, 68.47623, 68.43597, 68.39539, 68.35446, 
    68.31319, 68.2716, 68.22968, 68.18742, 68.14483, 68.10192, 68.05869, 
    68.01513, 67.97125, 67.92706, 67.88255, 67.83772, 67.79258, 67.74714, 
    67.70138, 67.65532, 67.60896, 67.56229, 67.51532, 67.46805, 67.42049, 
    67.37263, 67.32448, 67.27604, 67.2273, 67.17828, 67.12898, 67.0794, 
    67.02953, 66.97938, 66.92896, 66.87825, 66.82728, 66.77603, 66.72451, 
    66.67273, 66.62067, 66.56835, 66.51578, 66.46294, 66.40983, 66.35648, 
    66.30286, 66.24899, 66.19487, 66.1405, 66.08588, 66.03101, 65.9759, 
    65.92055, 65.86495, 65.80911, 65.75304, 65.69672, 65.64017, 65.5834, 
    65.52639, 65.46915, 65.41167, 65.35398, 65.29606, 65.23792, 65.17955, 
    65.12096, 65.06216, 65.00314, 64.9439, 64.88445, 64.82479, 64.76492, 
    64.70483, 64.64455,
  58.40317, 58.47733, 58.55138, 58.62534, 58.69918, 58.77293, 58.84658, 
    58.92011, 58.99355, 59.06687, 59.14009, 59.2132, 59.28619, 59.35909, 
    59.43186, 59.50453, 59.57708, 59.64952, 59.72184, 59.79405, 59.86614, 
    59.93812, 60.00998, 60.08171, 60.15333, 60.22483, 60.2962, 60.36745, 
    60.43858, 60.50958, 60.58046, 60.6512, 60.72182, 60.79232, 60.86268, 
    60.93291, 61.00301, 61.07298, 61.14281, 61.21251, 61.28207, 61.35149, 
    61.42078, 61.48993, 61.55894, 61.6278, 61.69652, 61.7651, 61.83353, 
    61.90182, 61.96997, 62.03796, 62.1058, 62.1735, 62.24104, 62.30843, 
    62.37566, 62.44274, 62.50966, 62.57643, 62.64303, 62.70948, 62.77576, 
    62.84188, 62.90784, 62.97364, 63.03926, 63.10472, 63.17001, 63.23513, 
    63.30008, 63.36486, 63.42946, 63.49389, 63.55813, 63.6222, 63.68609, 
    63.74981, 63.81333, 63.87667, 63.93983, 64.00281, 64.06559, 64.12818, 
    64.19059, 64.2528, 64.31482, 64.37664, 64.43826, 64.49969, 64.56092, 
    64.62195, 64.68277, 64.74339, 64.8038, 64.86401, 64.92401, 64.9838, 
    65.04337, 65.10274, 65.16188, 65.22081, 65.27953, 65.33801, 65.39629, 
    65.45433, 65.51215, 65.56975, 65.62711, 65.68425, 65.74116, 65.79783, 
    65.85426, 65.91047, 65.96643, 66.02215, 66.07763, 66.13287, 66.18786, 
    66.24261, 66.2971, 66.35134, 66.40533, 66.45908, 66.51256, 66.56578, 
    66.61874, 66.67145, 66.72389, 66.77607, 66.82797, 66.87962, 66.93098, 
    66.98208, 67.03291, 67.08345, 67.13372, 67.18371, 67.23341, 67.28284, 
    67.33197, 67.38082, 67.42938, 67.47765, 67.52563, 67.5733, 67.62069, 
    67.66777, 67.71455, 67.76103, 67.80721, 67.85307, 67.89864, 67.94389, 
    67.98882, 68.03344, 68.07774, 68.12173, 68.16539, 68.20873, 68.25175, 
    68.29444, 68.33681, 68.37884, 68.42053, 68.4619, 68.50293, 68.54362, 
    68.58397, 68.62398, 68.66364, 68.70296, 68.74193, 68.78055, 68.81881, 
    68.85673, 68.89428, 68.93148, 68.96832, 69.0048, 69.04091, 69.07666, 
    69.11204, 69.14705, 69.18169, 69.21596, 69.24985, 69.28336, 69.3165, 
    69.34925, 69.38162, 69.41361, 69.44521, 69.47643, 69.50725, 69.53768, 
    69.56772, 69.59737, 69.62661, 69.65546, 69.68391, 69.71195, 69.73959, 
    69.76683, 69.79366, 69.82008, 69.84609, 69.87169, 69.89687, 69.92165, 
    69.946, 69.96993, 69.99345, 70.01654, 70.03921, 70.06145, 70.08327, 
    70.10467, 70.12563, 70.14617, 70.16628, 70.18594, 70.20518, 70.22398, 
    70.24235, 70.26028, 70.27776, 70.29482, 70.31142, 70.32759, 70.34331, 
    70.35859, 70.37342, 70.3878, 70.40174, 70.41523, 70.42827, 70.44086, 
    70.453, 70.46468, 70.47591, 70.48669, 70.49702, 70.50689, 70.5163, 
    70.52525, 70.53375, 70.54179, 70.54938, 70.5565, 70.56316, 70.56937, 
    70.57511, 70.58039, 70.58521, 70.58958, 70.59348, 70.59691, 70.59988, 
    70.60239, 70.60444, 70.60603, 70.60715, 70.6078, 70.608, 70.60773, 
    70.607, 70.6058, 70.60415, 70.60203, 70.59944, 70.5964, 70.59289, 
    70.58891, 70.58448, 70.57959, 70.57423, 70.56842, 70.56214, 70.5554, 
    70.54821, 70.54055, 70.53244, 70.52387, 70.51484, 70.50536, 70.49541, 
    70.48502, 70.47417, 70.46287, 70.45111, 70.4389, 70.42624, 70.41312, 
    70.39957, 70.38556, 70.3711, 70.3562, 70.34085, 70.32506, 70.30882, 
    70.29214, 70.27503, 70.25747, 70.23947, 70.22104, 70.20217, 70.18286, 
    70.16312, 70.14295, 70.12234, 70.10132, 70.07986, 70.05797, 70.03565, 
    70.01292, 69.98975, 69.96617, 69.94218, 69.91776, 69.89292, 69.86767, 
    69.842, 69.81593, 69.78944, 69.76255, 69.73525, 69.70754, 69.67944, 
    69.65092, 69.62201, 69.5927, 69.563, 69.5329, 69.5024, 69.47151, 
    69.44024, 69.40858, 69.37653, 69.34409, 69.31128, 69.27808, 69.24451, 
    69.21056, 69.17623, 69.14153, 69.10647, 69.07103, 69.03522, 68.99905, 
    68.96252, 68.92562, 68.88837, 68.85075, 68.81278, 68.77446, 68.73579, 
    68.69676, 68.65739, 68.61767, 68.57761, 68.53721, 68.49646, 68.45538, 
    68.41396, 68.37221, 68.33012, 68.28771, 68.24497, 68.2019, 68.15851, 
    68.11479, 68.07076, 68.0264, 67.98173, 67.93674, 67.89145, 67.84584, 
    67.79993, 67.7537, 67.70718, 67.66035, 67.61321, 67.56578, 67.51806, 
    67.47003, 67.42172, 67.37312, 67.32422, 67.27504, 67.22557, 67.17582, 
    67.12579, 67.07547, 67.02488, 66.97401, 66.92287, 66.87147, 66.81979, 
    66.76783, 66.71561, 66.66313, 66.61039, 66.55738, 66.50411, 66.45059, 
    66.39681, 66.34278, 66.2885, 66.23396, 66.17918, 66.12415, 66.06887, 
    66.01335, 65.9576, 65.90159, 65.84535, 65.78888, 65.73217, 65.67522, 
    65.61806, 65.56065, 65.50302, 65.44516, 65.38708, 65.32877, 65.27025, 
    65.2115, 65.15254, 65.09336, 65.03397, 64.97436, 64.91454, 64.8545, 
    64.79427, 64.73382,
  58.47972, 58.55399, 58.62816, 58.70222, 58.77619, 58.85005, 58.92381, 
    58.99746, 59.071, 59.14444, 59.21777, 59.291, 59.36411, 59.43712, 
    59.51001, 59.5828, 59.65547, 59.72803, 59.80047, 59.8728, 59.94501, 
    60.01711, 60.08909, 60.16095, 60.23269, 60.30431, 60.3758, 60.44718, 
    60.51843, 60.58956, 60.66056, 60.73144, 60.80219, 60.87281, 60.9433, 
    61.01366, 61.08389, 61.15399, 61.22395, 61.29378, 61.36348, 61.43303, 
    61.50245, 61.57173, 61.64087, 61.70987, 61.77873, 61.84745, 61.91602, 
    61.98444, 62.05272, 62.12085, 62.18883, 62.25666, 62.32434, 62.39187, 
    62.45925, 62.52647, 62.59353, 62.66044, 62.72719, 62.79378, 62.86021, 
    62.92648, 62.99258, 63.05852, 63.12429, 63.1899, 63.25533, 63.3206, 
    63.3857, 63.45062, 63.51537, 63.57994, 63.64434, 63.70856, 63.77261, 
    63.83647, 63.90015, 63.96364, 64.02695, 64.09008, 64.15302, 64.21577, 
    64.27832, 64.34069, 64.40286, 64.46484, 64.52662, 64.5882, 64.64959, 
    64.71078, 64.77176, 64.83253, 64.8931, 64.95347, 65.01363, 65.07358, 
    65.13331, 65.19283, 65.25214, 65.31123, 65.3701, 65.42876, 65.48718, 
    65.54539, 65.60338, 65.66113, 65.71867, 65.77596, 65.83303, 65.88987, 
    65.94647, 66.00283, 66.05896, 66.11485, 66.17049, 66.22589, 66.28105, 
    66.33596, 66.39062, 66.44503, 66.49918, 66.55309, 66.60674, 66.66013, 
    66.71326, 66.76613, 66.81873, 66.87108, 66.92315, 66.97495, 67.02649, 
    67.07775, 67.12874, 67.17945, 67.22988, 67.28004, 67.32991, 67.3795, 
    67.4288, 67.47781, 67.52654, 67.57497, 67.62311, 67.67095, 67.7185, 
    67.76575, 67.81269, 67.85934, 67.90568, 67.95171, 67.99743, 68.04284, 
    68.08793, 68.13271, 68.17718, 68.22132, 68.26514, 68.30865, 68.35182, 
    68.39468, 68.43719, 68.47939, 68.52124, 68.56276, 68.60394, 68.64479, 
    68.6853, 68.72546, 68.76527, 68.80474, 68.84386, 68.88263, 68.92105, 
    68.95911, 68.99682, 69.03416, 69.07114, 69.10777, 69.14403, 69.17992, 
    69.21545, 69.2506, 69.28538, 69.31979, 69.35381, 69.38747, 69.42074, 
    69.45363, 69.48614, 69.51826, 69.55, 69.58134, 69.6123, 69.64285, 
    69.67302, 69.70279, 69.73216, 69.76114, 69.7897, 69.81787, 69.84563, 
    69.87299, 69.89994, 69.92648, 69.9526, 69.97831, 70.0036, 70.02848, 
    70.05295, 70.07699, 70.1006, 70.1238, 70.14658, 70.16892, 70.19084, 
    70.21233, 70.23339, 70.25401, 70.27421, 70.29398, 70.3133, 70.33218, 
    70.35064, 70.36864, 70.38622, 70.40334, 70.42003, 70.43627, 70.45206, 
    70.46741, 70.48232, 70.49677, 70.51077, 70.52432, 70.53742, 70.55006, 
    70.56226, 70.57401, 70.58529, 70.59612, 70.60649, 70.6164, 70.62586, 
    70.63486, 70.6434, 70.65148, 70.6591, 70.66625, 70.67295, 70.67918, 
    70.68495, 70.69026, 70.69511, 70.69949, 70.7034, 70.70686, 70.70984, 
    70.71236, 70.71442, 70.71601, 70.71714, 70.7178, 70.718, 70.71773, 
    70.717, 70.71579, 70.71413, 70.712, 70.7094, 70.70634, 70.70281, 
    70.69882, 70.69437, 70.68945, 70.68407, 70.67823, 70.67192, 70.66515, 
    70.65792, 70.65023, 70.64208, 70.63347, 70.6244, 70.61487, 70.60488, 
    70.59444, 70.58353, 70.57217, 70.56036, 70.5481, 70.53538, 70.5222, 
    70.50858, 70.49451, 70.47999, 70.46501, 70.44959, 70.43373, 70.41742, 
    70.40067, 70.38347, 70.36583, 70.34775, 70.32922, 70.31027, 70.29088, 
    70.27105, 70.25079, 70.23009, 70.20896, 70.1874, 70.16541, 70.143, 
    70.12016, 70.09689, 70.07321, 70.0491, 70.02457, 69.99963, 69.97427, 
    69.94849, 69.9223, 69.8957, 69.86869, 69.84127, 69.81345, 69.78522, 
    69.75658, 69.72755, 69.69811, 69.66827, 69.63805, 69.60742, 69.57641, 
    69.545, 69.51321, 69.48103, 69.44846, 69.4155, 69.38217, 69.34846, 
    69.31437, 69.2799, 69.24506, 69.20985, 69.17427, 69.13832, 69.10201, 
    69.06532, 69.02827, 68.99088, 68.95311, 68.91499, 68.87653, 68.8377, 
    68.79852, 68.759, 68.71912, 68.67891, 68.63835, 68.59745, 68.55621, 
    68.51464, 68.47273, 68.43049, 68.38792, 68.34502, 68.30179, 68.25824, 
    68.21436, 68.17017, 68.12565, 68.08082, 68.03568, 67.99021, 67.94444, 
    67.89837, 67.85198, 67.80529, 67.75829, 67.711, 67.66341, 67.61552, 
    67.56733, 67.51885, 67.47008, 67.42102, 67.37167, 67.32204, 67.27213, 
    67.22192, 67.17145, 67.12069, 67.06966, 67.01836, 66.96677, 66.91493, 
    66.86282, 66.81043, 66.75778, 66.70487, 66.6517, 66.59827, 66.54458, 
    66.49064, 66.43644, 66.38199, 66.32729, 66.27234, 66.21715, 66.16171, 
    66.10602, 66.05009, 65.99393, 65.93753, 65.88089, 65.82402, 65.76691, 
    65.70958, 65.65202, 65.59422, 65.5362, 65.47796, 65.41949, 65.3608, 
    65.3019, 65.24277, 65.18343, 65.12388, 65.06411, 65.00413, 64.94394, 
    64.88354, 64.82294,
  58.55611, 58.63049, 58.70476, 58.77894, 58.85302, 58.92699, 59.00085, 
    59.07462, 59.14828, 59.22184, 59.29528, 59.36862, 59.44185, 59.51498, 
    59.58799, 59.66089, 59.73368, 59.80636, 59.87892, 59.95137, 60.0237, 
    60.09592, 60.16802, 60.24001, 60.31187, 60.38361, 60.45523, 60.52673, 
    60.59811, 60.66936, 60.74049, 60.8115, 60.88237, 60.95312, 61.02374, 
    61.09423, 61.16459, 61.23482, 61.30492, 61.37488, 61.4447, 61.51439, 
    61.58395, 61.65336, 61.72263, 61.79177, 61.86076, 61.92962, 61.99832, 
    62.06688, 62.1353, 62.20357, 62.27169, 62.33966, 62.40748, 62.47515, 
    62.54267, 62.61003, 62.67724, 62.74429, 62.81118, 62.87791, 62.94448, 
    63.01089, 63.07714, 63.14323, 63.20915, 63.2749, 63.34048, 63.4059, 
    63.47115, 63.53622, 63.60112, 63.66584, 63.73039, 63.79476, 63.85896, 
    63.92297, 63.9868, 64.05045, 64.11391, 64.17719, 64.24028, 64.30318, 
    64.3659, 64.42842, 64.49075, 64.55288, 64.61482, 64.67656, 64.73811, 
    64.79945, 64.86059, 64.92152, 64.98225, 65.04278, 65.1031, 65.1632, 
    65.2231, 65.28278, 65.34225, 65.4015, 65.46053, 65.51935, 65.57794, 
    65.63631, 65.69446, 65.75238, 65.81007, 65.86753, 65.92477, 65.98177, 
    66.03853, 66.09506, 66.15135, 66.20741, 66.26321, 66.31878, 66.3741, 
    66.42918, 66.484, 66.53858, 66.5929, 66.64697, 66.70078, 66.75434, 
    66.80764, 66.86067, 66.91345, 66.96596, 67.0182, 67.07017, 67.12187, 
    67.1733, 67.22446, 67.27533, 67.32594, 67.37625, 67.42629, 67.47604, 
    67.52551, 67.57469, 67.62358, 67.67218, 67.72049, 67.76849, 67.81621, 
    67.86362, 67.91073, 67.95753, 68.00404, 68.05023, 68.09612, 68.14169, 
    68.18695, 68.23189, 68.27652, 68.32082, 68.36481, 68.40847, 68.45181, 
    68.49482, 68.5375, 68.57984, 68.62186, 68.66354, 68.70488, 68.74588, 
    68.78654, 68.82685, 68.86682, 68.90645, 68.94572, 68.98464, 69.02321, 
    69.06142, 69.09927, 69.13677, 69.1739, 69.21068, 69.24708, 69.28312, 
    69.31879, 69.35408, 69.38901, 69.42355, 69.45773, 69.49152, 69.52493, 
    69.55795, 69.5906, 69.62286, 69.65472, 69.6862, 69.71729, 69.74798, 
    69.77827, 69.80817, 69.83767, 69.86677, 69.89546, 69.92375, 69.95164, 
    69.97911, 70.00617, 70.03283, 70.05907, 70.08489, 70.1103, 70.13529, 
    70.15986, 70.18401, 70.20773, 70.23103, 70.25391, 70.27636, 70.29838, 
    70.31996, 70.34112, 70.36184, 70.38213, 70.40198, 70.42139, 70.44037, 
    70.4589, 70.477, 70.49464, 70.51186, 70.52862, 70.54493, 70.5608, 
    70.57622, 70.59119, 70.60571, 70.61978, 70.6334, 70.64656, 70.65926, 
    70.67152, 70.68331, 70.69466, 70.70554, 70.71596, 70.72592, 70.73542, 
    70.74446, 70.75304, 70.76116, 70.76881, 70.77601, 70.78274, 70.78899, 
    70.79479, 70.80013, 70.805, 70.80939, 70.81333, 70.8168, 70.8198, 
    70.82233, 70.8244, 70.826, 70.82714, 70.8278, 70.828, 70.82773, 70.82699, 
    70.82578, 70.82411, 70.82197, 70.81936, 70.81628, 70.81274, 70.80873, 
    70.80426, 70.79932, 70.79391, 70.78804, 70.7817, 70.7749, 70.76763, 
    70.75991, 70.75172, 70.74306, 70.73395, 70.72437, 70.71434, 70.70384, 
    70.69289, 70.68148, 70.66961, 70.65729, 70.64451, 70.63127, 70.61758, 
    70.60345, 70.58885, 70.57381, 70.55832, 70.54238, 70.52599, 70.50916, 
    70.49188, 70.47417, 70.456, 70.43739, 70.41835, 70.39886, 70.37894, 
    70.35859, 70.3378, 70.31657, 70.29492, 70.27283, 70.25032, 70.22738, 
    70.20401, 70.18021, 70.156, 70.13136, 70.10631, 70.08083, 70.05495, 
    70.02864, 70.00192, 69.97479, 69.94725, 69.9193, 69.89095, 69.86219, 
    69.83303, 69.80347, 69.77351, 69.74315, 69.71239, 69.68125, 69.64971, 
    69.61778, 69.58546, 69.55276, 69.51967, 69.4862, 69.45235, 69.41811, 
    69.38351, 69.34853, 69.31317, 69.27744, 69.24135, 69.20489, 69.16806, 
    69.13087, 69.09332, 69.0554, 69.01714, 68.97851, 68.93953, 68.9002, 
    68.86053, 68.8205, 68.78013, 68.73942, 68.69836, 68.65697, 68.61523, 
    68.57317, 68.53077, 68.48804, 68.44498, 68.40159, 68.35787, 68.31384, 
    68.26948, 68.2248, 68.17981, 68.1345, 68.08887, 68.04295, 67.9967, 
    67.95015, 67.9033, 67.85614, 67.80868, 67.76092, 67.71287, 67.66451, 
    67.61587, 67.56693, 67.51771, 67.46819, 67.4184, 67.36831, 67.31795, 
    67.2673, 67.21638, 67.16518, 67.11371, 67.06197, 67.00995, 66.95766, 
    66.90512, 66.8523, 66.79922, 66.74589, 66.69229, 66.63844, 66.58433, 
    66.52996, 66.47535, 66.42048, 66.36536, 66.31001, 66.2544, 66.19855, 
    66.14246, 66.08614, 66.02957, 65.97276, 65.91573, 65.85846, 65.80096, 
    65.74323, 65.68527, 65.62709, 65.56869, 65.51006, 65.45121, 65.39214, 
    65.33286, 65.27335, 65.21364, 65.15371, 65.09357, 65.03322, 64.97266, 
    64.9119,
  58.63231, 58.7068, 58.78119, 58.85547, 58.92966, 59.00375, 59.07773, 
    59.15161, 59.22538, 59.29905, 59.37261, 59.44607, 59.51942, 59.59266, 
    59.66578, 59.7388, 59.81171, 59.88451, 59.95719, 60.02976, 60.10222, 
    60.17456, 60.24678, 60.31888, 60.39087, 60.46274, 60.53448, 60.60611, 
    60.67761, 60.74899, 60.82025, 60.89138, 60.96238, 61.03326, 61.10401, 
    61.17463, 61.24512, 61.31548, 61.3857, 61.4558, 61.52575, 61.59558, 
    61.66526, 61.73481, 61.80422, 61.87349, 61.94262, 62.01161, 62.08045, 
    62.14915, 62.2177, 62.28611, 62.35437, 62.42249, 62.49045, 62.55826, 
    62.62592, 62.69342, 62.76077, 62.82796, 62.895, 62.96187, 63.02859, 
    63.09515, 63.16154, 63.22777, 63.29383, 63.35974, 63.42547, 63.49103, 
    63.55642, 63.62165, 63.6867, 63.75157, 63.81627, 63.88079, 63.94514, 
    64.0093, 64.07329, 64.13708, 64.20071, 64.26414, 64.32738, 64.39044, 
    64.45331, 64.51599, 64.57848, 64.64076, 64.70286, 64.76476, 64.82646, 
    64.88795, 64.94926, 65.01035, 65.07124, 65.13193, 65.19241, 65.25267, 
    65.31273, 65.37257, 65.4322, 65.49162, 65.55081, 65.60979, 65.66854, 
    65.72708, 65.78539, 65.84348, 65.90133, 65.95896, 66.01636, 66.07352, 
    66.13045, 66.18714, 66.2436, 66.29982, 66.3558, 66.41153, 66.46702, 
    66.52225, 66.57725, 66.632, 66.68649, 66.74072, 66.7947, 66.84843, 
    66.90189, 66.95509, 67.00803, 67.06071, 67.11312, 67.16526, 67.21712, 
    67.26872, 67.32005, 67.37109, 67.42186, 67.47234, 67.52255, 67.57247, 
    67.62211, 67.67146, 67.72051, 67.76928, 67.81775, 67.86592, 67.9138, 
    67.96138, 68.00866, 68.05563, 68.10229, 68.14865, 68.1947, 68.24044, 
    68.28586, 68.33097, 68.37576, 68.42023, 68.46438, 68.5082, 68.5517, 
    68.59486, 68.6377, 68.68021, 68.72238, 68.76422, 68.80573, 68.84688, 
    68.8877, 68.92817, 68.96829, 69.00807, 69.0475, 69.08658, 69.1253, 
    69.16366, 69.20167, 69.23931, 69.2766, 69.31351, 69.35007, 69.38625, 
    69.42207, 69.4575, 69.49257, 69.52726, 69.56158, 69.5955, 69.62906, 
    69.66222, 69.69501, 69.72739, 69.7594, 69.79102, 69.82223, 69.85305, 
    69.88348, 69.91351, 69.94313, 69.97236, 70.00117, 70.02959, 70.05759, 
    70.08519, 70.11237, 70.13914, 70.1655, 70.19144, 70.21696, 70.24206, 
    70.26674, 70.291, 70.31483, 70.33823, 70.36121, 70.38377, 70.40588, 
    70.42757, 70.44882, 70.46964, 70.49002, 70.50996, 70.52946, 70.54853, 
    70.56715, 70.58533, 70.60307, 70.62035, 70.63719, 70.65358, 70.66953, 
    70.68502, 70.70006, 70.71465, 70.72878, 70.74246, 70.75569, 70.76846, 
    70.78077, 70.79262, 70.80401, 70.81494, 70.82542, 70.83543, 70.84498, 
    70.85406, 70.86268, 70.87083, 70.87853, 70.88576, 70.89252, 70.89881, 
    70.90463, 70.91, 70.91489, 70.91931, 70.92326, 70.92675, 70.92976, 
    70.93231, 70.93439, 70.936, 70.93713, 70.9378, 70.938, 70.93773, 
    70.93698, 70.93578, 70.93409, 70.93194, 70.92932, 70.92622, 70.92267, 
    70.91864, 70.91415, 70.90918, 70.90375, 70.89784, 70.89148, 70.88464, 
    70.87734, 70.86958, 70.86135, 70.85265, 70.8435, 70.83388, 70.82379, 
    70.81325, 70.80224, 70.79077, 70.77885, 70.76646, 70.75362, 70.74033, 
    70.72658, 70.71237, 70.69771, 70.68259, 70.66703, 70.65102, 70.63456, 
    70.61765, 70.60029, 70.58248, 70.56423, 70.54555, 70.52641, 70.50684, 
    70.48682, 70.46638, 70.44549, 70.42417, 70.40241, 70.38023, 70.35761, 
    70.33456, 70.31109, 70.28719, 70.26286, 70.23812, 70.21295, 70.18736, 
    70.16135, 70.13493, 70.1081, 70.08085, 70.05319, 70.02512, 69.99664, 
    69.96776, 69.93848, 69.90878, 69.87869, 69.84821, 69.81732, 69.78604, 
    69.75436, 69.7223, 69.68984, 69.65701, 69.62378, 69.59016, 69.55618, 
    69.5218, 69.48705, 69.45192, 69.41642, 69.38055, 69.34431, 69.30769, 
    69.27072, 69.23338, 69.19568, 69.15762, 69.11919, 69.08041, 69.04129, 
    69.0018, 68.96197, 68.92179, 68.88126, 68.84039, 68.79918, 68.75763, 
    68.71574, 68.67351, 68.63095, 68.58806, 68.54484, 68.50129, 68.45741, 
    68.41322, 68.3687, 68.32385, 68.27869, 68.23322, 68.18744, 68.14134, 
    68.09493, 68.04822, 68.0012, 67.95387, 67.90625, 67.85832, 67.8101, 
    67.76158, 67.71277, 67.66367, 67.61427, 67.5646, 67.51463, 67.46438, 
    67.41385, 67.36304, 67.31194, 67.26058, 67.20894, 67.15703, 67.10484, 
    67.0524, 66.99968, 66.94669, 66.89345, 66.83994, 66.78618, 66.73216, 
    66.67788, 66.62335, 66.56857, 66.51353, 66.45825, 66.40273, 66.34695, 
    66.29094, 66.23469, 66.17819, 66.12146, 66.06449, 66.00729, 65.94986, 
    65.8922, 65.8343, 65.77618, 65.71783, 65.65926, 65.60047, 65.54146, 
    65.48223, 65.42278, 65.36312, 65.30324, 65.24315, 65.18285, 65.12234, 
    65.06162, 65.0007,
  58.70833, 58.78293, 58.85743, 58.93183, 59.00613, 59.08032, 59.15442, 
    59.22841, 59.3023, 59.37608, 59.44976, 59.52333, 59.59679, 59.67015, 
    59.7434, 59.81654, 59.88956, 59.96248, 60.03528, 60.10797, 60.18055, 
    60.25301, 60.32536, 60.39758, 60.46969, 60.54168, 60.61355, 60.6853, 
    60.75693, 60.82844, 60.89982, 60.97108, 61.04221, 61.11322, 61.1841, 
    61.25484, 61.32547, 61.39595, 61.46631, 61.53654, 61.60663, 61.67658, 
    61.7464, 61.81609, 61.88563, 61.95504, 62.0243, 62.09343, 62.16241, 
    62.23124, 62.29993, 62.36848, 62.43688, 62.50513, 62.57323, 62.64119, 
    62.70898, 62.77663, 62.84412, 62.91146, 62.97864, 63.04566, 63.11252, 
    63.17922, 63.24577, 63.31214, 63.37835, 63.4444, 63.51028, 63.57599, 
    63.64154, 63.70691, 63.77211, 63.83713, 63.90198, 63.96666, 64.03115, 
    64.09547, 64.15961, 64.22356, 64.28734, 64.35092, 64.41432, 64.47754, 
    64.54056, 64.60339, 64.66604, 64.72849, 64.79074, 64.85279, 64.91465, 
    64.97631, 65.03777, 65.09902, 65.16007, 65.22092, 65.28156, 65.34199, 
    65.40221, 65.46221, 65.522, 65.58158, 65.64094, 65.70008, 65.759, 
    65.8177, 65.87617, 65.93442, 65.99244, 66.05024, 66.1078, 66.16513, 
    66.22223, 66.27908, 66.33571, 66.39209, 66.44823, 66.50414, 66.55979, 
    66.6152, 66.67036, 66.72527, 66.77993, 66.83434, 66.88849, 66.94238, 
    66.99601, 67.04939, 67.10249, 67.15533, 67.20791, 67.26022, 67.31226, 
    67.36402, 67.41551, 67.46673, 67.51766, 67.56832, 67.61869, 67.66879, 
    67.71858, 67.7681, 67.81733, 67.86626, 67.9149, 67.96324, 68.01128, 
    68.05903, 68.10648, 68.15361, 68.20045, 68.24697, 68.29318, 68.33909, 
    68.38467, 68.42995, 68.4749, 68.51953, 68.56384, 68.60783, 68.65149, 
    68.69482, 68.73782, 68.78049, 68.82282, 68.86482, 68.90648, 68.9478, 
    68.98877, 69.0294, 69.06969, 69.10962, 69.1492, 69.18843, 69.2273, 
    69.26582, 69.30398, 69.34177, 69.37921, 69.41628, 69.45298, 69.48931, 
    69.52527, 69.56086, 69.59607, 69.63091, 69.66536, 69.69943, 69.73312, 
    69.76643, 69.79935, 69.83189, 69.86402, 69.89577, 69.92712, 69.95808, 
    69.98863, 70.01879, 70.04855, 70.0779, 70.10684, 70.13538, 70.16351, 
    70.19122, 70.21853, 70.24542, 70.2719, 70.29795, 70.32359, 70.3488, 
    70.37359, 70.39796, 70.4219, 70.44541, 70.46849, 70.49115, 70.51337, 
    70.53515, 70.5565, 70.57742, 70.59789, 70.61793, 70.63752, 70.65667, 
    70.67538, 70.69364, 70.71146, 70.72883, 70.74575, 70.76221, 70.77824, 
    70.7938, 70.80891, 70.82357, 70.83778, 70.85152, 70.86481, 70.87764, 
    70.89001, 70.90192, 70.91336, 70.92435, 70.93487, 70.94493, 70.95452, 
    70.96365, 70.97231, 70.98051, 70.98824, 70.9955, 71.0023, 71.00862, 
    71.01447, 71.01986, 71.02477, 71.02922, 71.03319, 71.03669, 71.03973, 
    71.04228, 71.04437, 71.04598, 71.04713, 71.0478, 71.048, 71.04772, 
    71.04698, 71.04576, 71.04408, 71.04191, 71.03928, 71.03617, 71.03259, 
    71.02854, 71.02402, 71.01904, 71.01358, 71.00765, 71.00125, 70.99438, 
    70.98705, 70.97925, 70.97098, 70.96224, 70.95303, 70.94337, 70.93324, 
    70.92265, 70.91158, 70.90006, 70.88808, 70.87564, 70.86274, 70.84938, 
    70.83556, 70.82128, 70.80656, 70.79137, 70.77573, 70.75964, 70.7431, 
    70.72611, 70.70867, 70.69078, 70.67245, 70.65367, 70.63445, 70.61478, 
    70.59468, 70.57413, 70.55315, 70.53174, 70.50988, 70.48759, 70.46487, 
    70.44172, 70.41814, 70.39413, 70.3697, 70.34484, 70.31956, 70.29385, 
    70.26773, 70.2412, 70.21424, 70.18687, 70.15909, 70.13089, 70.10229, 
    70.07328, 70.04387, 70.01405, 69.98383, 69.95321, 69.92219, 69.89078, 
    69.85896, 69.82677, 69.79417, 69.76119, 69.72782, 69.69407, 69.65993, 
    69.62542, 69.59052, 69.55525, 69.51961, 69.48359, 69.4472, 69.41044, 
    69.37331, 69.33582, 69.29797, 69.25975, 69.22118, 69.18225, 69.14296, 
    69.10332, 69.06333, 69.02299, 68.98232, 68.94128, 68.89991, 68.8582, 
    68.81615, 68.77377, 68.73104, 68.68799, 68.64461, 68.60089, 68.55685, 
    68.5125, 68.46781, 68.42281, 68.37749, 68.33185, 68.2859, 68.23963, 
    68.19305, 68.14618, 68.09899, 68.0515, 68.00371, 67.95561, 67.90723, 
    67.85854, 67.80956, 67.76028, 67.71072, 67.66088, 67.61074, 67.56033, 
    67.50963, 67.45865, 67.40739, 67.35585, 67.30405, 67.25196, 67.19962, 
    67.147, 67.09411, 67.04095, 66.98754, 66.93387, 66.87994, 66.82574, 
    66.7713, 66.71661, 66.66165, 66.60645, 66.551, 66.49531, 66.43937, 
    66.38319, 66.32677, 66.27011, 66.21321, 66.15607, 66.09871, 66.04111, 
    65.98328, 65.92522, 65.86694, 65.80843, 65.74969, 65.69073, 65.63156, 
    65.57217, 65.51256, 65.45274, 65.39269, 65.33244, 65.27198, 65.21131, 
    65.15043, 65.08935,
  58.78417, 58.85888, 58.93349, 59.008, 59.08241, 59.15672, 59.23093, 
    59.30503, 59.37903, 59.45293, 59.52673, 59.60041, 59.67399, 59.74747, 
    59.82083, 59.89409, 59.96723, 60.04027, 60.11319, 60.186, 60.2587, 
    60.33128, 60.40375, 60.4761, 60.54833, 60.62045, 60.69244, 60.76432, 
    60.83607, 60.9077, 60.97921, 61.0506, 61.12186, 61.19299, 61.264, 
    61.33488, 61.40563, 61.47625, 61.54674, 61.6171, 61.68732, 61.75741, 
    61.82736, 61.89718, 61.96686, 62.0364, 62.1058, 62.17506, 62.24418, 
    62.31316, 62.38199, 62.45067, 62.51921, 62.5876, 62.65585, 62.72394, 
    62.79188, 62.85967, 62.9273, 62.99478, 63.06211, 63.12927, 63.19628, 
    63.26313, 63.32981, 63.39634, 63.4627, 63.52889, 63.59492, 63.66078, 
    63.72647, 63.792, 63.85735, 63.92252, 63.98752, 64.05235, 64.117, 
    64.18147, 64.24576, 64.30987, 64.37379, 64.43754, 64.5011, 64.56447, 
    64.62765, 64.69064, 64.75343, 64.81604, 64.87846, 64.94067, 65.00269, 
    65.06451, 65.12612, 65.18754, 65.24875, 65.30975, 65.37055, 65.43114, 
    65.49152, 65.55169, 65.61165, 65.67139, 65.73091, 65.79021, 65.8493, 
    65.90816, 65.9668, 66.02522, 66.0834, 66.14137, 66.1991, 66.25659, 
    66.31386, 66.37088, 66.42767, 66.48422, 66.54053, 66.5966, 66.65243, 
    66.708, 66.76333, 66.81841, 66.87324, 66.92781, 66.98213, 67.03619, 
    67.09, 67.14354, 67.19682, 67.24982, 67.30257, 67.35505, 67.40726, 
    67.4592, 67.51086, 67.56224, 67.61334, 67.66417, 67.71471, 67.76497, 
    67.81494, 67.86463, 67.91402, 67.96313, 68.01193, 68.06045, 68.10866, 
    68.15657, 68.20418, 68.25149, 68.29848, 68.34518, 68.39156, 68.43763, 
    68.48338, 68.52882, 68.57394, 68.61874, 68.66322, 68.70737, 68.75119, 
    68.79469, 68.83784, 68.88068, 68.92317, 68.96533, 69.00715, 69.04862, 
    69.08976, 69.13055, 69.17099, 69.21108, 69.25082, 69.29021, 69.32923, 
    69.3679, 69.40622, 69.44417, 69.48175, 69.51897, 69.55582, 69.5923, 
    69.62841, 69.66415, 69.69951, 69.73449, 69.76909, 69.80331, 69.83714, 
    69.87058, 69.90364, 69.93631, 69.96859, 70.00047, 70.03196, 70.06305, 
    70.09374, 70.12403, 70.15392, 70.1834, 70.21246, 70.24113, 70.26938, 
    70.29722, 70.32465, 70.35166, 70.37825, 70.40443, 70.43018, 70.45551, 
    70.48041, 70.50488, 70.52893, 70.55255, 70.57574, 70.5985, 70.62082, 
    70.64271, 70.66415, 70.68517, 70.70574, 70.72587, 70.74555, 70.76479, 
    70.78359, 70.80194, 70.81984, 70.83729, 70.85429, 70.87084, 70.88693, 
    70.90257, 70.91776, 70.93249, 70.94675, 70.96056, 70.97392, 70.98681, 
    70.99924, 71.01121, 71.02271, 71.03374, 71.04432, 71.05443, 71.06406, 
    71.07324, 71.08195, 71.09018, 71.09795, 71.10525, 71.11207, 71.11842, 
    71.12431, 71.12972, 71.13466, 71.13912, 71.14312, 71.14664, 71.14968, 
    71.15225, 71.15435, 71.15598, 71.15713, 71.1578, 71.158, 71.15772, 
    71.15697, 71.15575, 71.15405, 71.15188, 71.14923, 71.14611, 71.14252, 
    71.13845, 71.13391, 71.1289, 71.12341, 71.11745, 71.11102, 71.10412, 
    71.09675, 71.08891, 71.0806, 71.07182, 71.06258, 71.05286, 71.04268, 
    71.03203, 71.02092, 71.00935, 70.99731, 70.9848, 70.97184, 70.95841, 
    70.94453, 70.93018, 70.91539, 70.90013, 70.88441, 70.86825, 70.85163, 
    70.83456, 70.81704, 70.79906, 70.78065, 70.76178, 70.74247, 70.72271, 
    70.70251, 70.68188, 70.6608, 70.63927, 70.61732, 70.59493, 70.57211, 
    70.54884, 70.52516, 70.50104, 70.47649, 70.45152, 70.42613, 70.40031, 
    70.37407, 70.34741, 70.32034, 70.29285, 70.26494, 70.23663, 70.20789, 
    70.17876, 70.14922, 70.11926, 70.08891, 70.05816, 70.02701, 69.99545, 
    69.96351, 69.93117, 69.89844, 69.86532, 69.83181, 69.79792, 69.76364, 
    69.72898, 69.69394, 69.65852, 69.62273, 69.58656, 69.55002, 69.51311, 
    69.47583, 69.43819, 69.40018, 69.36181, 69.32308, 69.284, 69.24455, 
    69.20476, 69.16461, 69.12412, 69.08327, 69.04209, 69.00056, 68.95869, 
    68.91647, 68.87392, 68.83104, 68.78783, 68.74428, 68.7004, 68.6562, 
    68.61167, 68.56683, 68.52165, 68.47617, 68.43037, 68.38425, 68.33781, 
    68.29108, 68.24403, 68.19667, 68.14901, 68.10105, 68.05279, 68.00423, 
    67.95538, 67.90623, 67.85679, 67.80706, 67.75704, 67.70673, 67.65615, 
    67.60528, 67.55413, 67.5027, 67.451, 67.39902, 67.34677, 67.29425, 
    67.24146, 67.18841, 67.13509, 67.0815, 67.02766, 66.97356, 66.9192, 
    66.86459, 66.80972, 66.7546, 66.69923, 66.64361, 66.58775, 66.53165, 
    66.4753, 66.41871, 66.36188, 66.30481, 66.24751, 66.18998, 66.13221, 
    66.07422, 66.01599, 65.95754, 65.89886, 65.83997, 65.78085, 65.72151, 
    65.66195, 65.60218, 65.54219, 65.48199, 65.42158, 65.36095, 65.30012, 
    65.23908, 65.17783,
  58.85983, 58.93465, 59.00937, 59.08399, 59.15851, 59.23293, 59.30725, 
    59.38147, 59.45559, 59.5296, 59.60351, 59.67731, 59.75101, 59.8246, 
    59.89808, 59.97145, 60.04472, 60.11787, 60.19091, 60.26385, 60.33667, 
    60.40937, 60.48196, 60.55443, 60.62679, 60.69902, 60.77114, 60.84315, 
    60.91503, 60.98679, 61.05842, 61.12994, 61.20132, 61.27259, 61.34372, 
    61.41473, 61.48561, 61.55637, 61.62698, 61.69748, 61.76783, 61.83805, 
    61.90814, 61.97809, 62.04791, 62.11758, 62.18712, 62.25652, 62.32578, 
    62.39489, 62.46386, 62.53268, 62.60136, 62.6699, 62.73828, 62.80651, 
    62.8746, 62.94253, 63.01031, 63.07793, 63.1454, 63.21271, 63.27986, 
    63.34686, 63.41369, 63.48036, 63.54687, 63.61321, 63.67939, 63.7454, 
    63.81124, 63.87691, 63.94241, 64.00774, 64.07289, 64.13787, 64.20267, 
    64.2673, 64.33174, 64.39601, 64.46009, 64.52399, 64.5877, 64.65122, 
    64.71456, 64.77771, 64.84067, 64.90343, 64.966, 65.02837, 65.09055, 
    65.15253, 65.21431, 65.27589, 65.33726, 65.39843, 65.45939, 65.52014, 
    65.58069, 65.64102, 65.70113, 65.76104, 65.82073, 65.8802, 65.93945, 
    65.99847, 66.05728, 66.11586, 66.17422, 66.23235, 66.29024, 66.34791, 
    66.40533, 66.46253, 66.51949, 66.57621, 66.63269, 66.68893, 66.74492, 
    66.80067, 66.85616, 66.91142, 66.96641, 67.02116, 67.07564, 67.12988, 
    67.18385, 67.23756, 67.29101, 67.34419, 67.39711, 67.44975, 67.50214, 
    67.55424, 67.60607, 67.65762, 67.7089, 67.7599, 67.81061, 67.86104, 
    67.91118, 67.96104, 68.0106, 68.05988, 68.10885, 68.15753, 68.20592, 
    68.254, 68.30177, 68.34925, 68.39642, 68.44328, 68.48983, 68.53606, 
    68.58199, 68.62759, 68.67287, 68.71784, 68.76248, 68.8068, 68.85078, 
    68.89445, 68.93777, 68.98077, 69.02343, 69.06575, 69.10773, 69.14937, 
    69.19066, 69.23161, 69.27221, 69.31246, 69.35236, 69.3919, 69.43108, 
    69.46991, 69.50838, 69.54648, 69.58422, 69.62159, 69.65859, 69.69523, 
    69.73148, 69.76736, 69.80287, 69.838, 69.87275, 69.90711, 69.94109, 
    69.97468, 70.00787, 70.04069, 70.0731, 70.10512, 70.13674, 70.16797, 
    70.19879, 70.22922, 70.25923, 70.28884, 70.31804, 70.34683, 70.37521, 
    70.40318, 70.43073, 70.45786, 70.48457, 70.51086, 70.53673, 70.56217, 
    70.58719, 70.61178, 70.63594, 70.65967, 70.68296, 70.70583, 70.72825, 
    70.75024, 70.77179, 70.79289, 70.81356, 70.83379, 70.85356, 70.87289, 
    70.89178, 70.91022, 70.9282, 70.94574, 70.96281, 70.97945, 70.99561, 
    71.01133, 71.02659, 71.04139, 71.05573, 71.0696, 71.08302, 71.09597, 
    71.10846, 71.12048, 71.13204, 71.14314, 71.15376, 71.16392, 71.17361, 
    71.18282, 71.19157, 71.19984, 71.20765, 71.21498, 71.22185, 71.22823, 
    71.23415, 71.23958, 71.24454, 71.24903, 71.25304, 71.25658, 71.25964, 
    71.26223, 71.26434, 71.26597, 71.26712, 71.2678, 71.268, 71.26772, 
    71.26697, 71.26574, 71.26403, 71.26185, 71.25919, 71.25605, 71.25244, 
    71.24835, 71.24379, 71.23875, 71.23324, 71.22725, 71.22079, 71.21386, 
    71.20645, 71.19857, 71.19022, 71.1814, 71.1721, 71.16235, 71.15211, 
    71.14141, 71.13025, 71.11861, 71.10651, 71.09396, 71.08092, 71.06744, 
    71.05349, 71.03908, 71.02421, 71.00887, 70.99309, 70.97684, 70.96014, 
    70.94299, 70.92538, 70.90733, 70.88882, 70.86987, 70.85046, 70.83062, 
    70.81033, 70.78959, 70.76841, 70.74679, 70.72473, 70.70224, 70.67931, 
    70.65594, 70.63214, 70.60792, 70.58326, 70.55817, 70.53266, 70.50673, 
    70.48037, 70.45359, 70.42639, 70.39878, 70.37075, 70.34231, 70.31345, 
    70.28419, 70.25451, 70.22443, 70.19395, 70.16306, 70.13177, 70.10008, 
    70.068, 70.03552, 70.00265, 69.96939, 69.93574, 69.9017, 69.86728, 
    69.83247, 69.79728, 69.76172, 69.72578, 69.68945, 69.65276, 69.61571, 
    69.57828, 69.54048, 69.50232, 69.46379, 69.42491, 69.38567, 69.34607, 
    69.30611, 69.26581, 69.22516, 69.18415, 69.1428, 69.10111, 69.05907, 
    69.0167, 68.97399, 68.93095, 68.88757, 68.84385, 68.79981, 68.75544, 
    68.71075, 68.66573, 68.6204, 68.57475, 68.52877, 68.48249, 68.43589, 
    68.38898, 68.34177, 68.29424, 68.24641, 68.19828, 68.14985, 68.10112, 
    68.0521, 68.00278, 67.95317, 67.90327, 67.85308, 67.8026, 67.75185, 
    67.70081, 67.64949, 67.59789, 67.54601, 67.49387, 67.44144, 67.38876, 
    67.33579, 67.28257, 67.22908, 67.17532, 67.12132, 67.06704, 67.01251, 
    66.95773, 66.90269, 66.8474, 66.79186, 66.73608, 66.68005, 66.62377, 
    66.56725, 66.5105, 66.4535, 66.39626, 66.3388, 66.2811, 66.22317, 66.165, 
    66.10661, 66.048, 65.98916, 65.93009, 65.8708, 65.8113, 65.75158, 
    65.69164, 65.63149, 65.57112, 65.51054, 65.44976, 65.38876, 65.32757, 
    65.26616,
  58.9353, 59.01023, 59.08506, 59.15979, 59.23442, 59.30896, 59.38339, 
    59.45773, 59.53195, 59.60608, 59.6801, 59.75402, 59.82784, 59.90154, 
    59.97514, 60.04864, 60.12202, 60.19529, 60.26846, 60.34151, 60.41444, 
    60.48727, 60.55998, 60.63258, 60.70506, 60.77742, 60.84967, 60.92179, 
    60.9938, 61.06569, 61.13745, 61.20909, 61.28061, 61.352, 61.42326, 
    61.4944, 61.56541, 61.6363, 61.70705, 61.77767, 61.84816, 61.91851, 
    61.98874, 62.05882, 62.12878, 62.19859, 62.26826, 62.3378, 62.40719, 
    62.47644, 62.54555, 62.61452, 62.68333, 62.75201, 62.82053, 62.88891, 
    62.95713, 63.02521, 63.09313, 63.1609, 63.22851, 63.29597, 63.36327, 
    63.4304, 63.49738, 63.5642, 63.63086, 63.69735, 63.76368, 63.82984, 
    63.89583, 63.96165, 64.02731, 64.09278, 64.15809, 64.22322, 64.28818, 
    64.35296, 64.41756, 64.48197, 64.54621, 64.61027, 64.67413, 64.73782, 
    64.80132, 64.86462, 64.92773, 64.99065, 65.05339, 65.11592, 65.17826, 
    65.24039, 65.30234, 65.36407, 65.42561, 65.48694, 65.54807, 65.60898, 
    65.66969, 65.73019, 65.79047, 65.85054, 65.91039, 65.97002, 66.02944, 
    66.08864, 66.14761, 66.20635, 66.26488, 66.32317, 66.38123, 66.43906, 
    66.49667, 66.55403, 66.61116, 66.66805, 66.72469, 66.78111, 66.83727, 
    66.89318, 66.94885, 67.00427, 67.05944, 67.11435, 67.16901, 67.22341, 
    67.27756, 67.33144, 67.38506, 67.43842, 67.49151, 67.54433, 67.59688, 
    67.64915, 67.70116, 67.75288, 67.80433, 67.8555, 67.90638, 67.95699, 
    68.00729, 68.05733, 68.10706, 68.1565, 68.20565, 68.2545, 68.30305, 
    68.35131, 68.39926, 68.44691, 68.49424, 68.54128, 68.58799, 68.6344, 
    68.68049, 68.72626, 68.77171, 68.81684, 68.86165, 68.90614, 68.95029, 
    68.99412, 69.03761, 69.08076, 69.12359, 69.16607, 69.20821, 69.25002, 
    69.29147, 69.33258, 69.37334, 69.41375, 69.45381, 69.49351, 69.53285, 
    69.57184, 69.61046, 69.64872, 69.68661, 69.72414, 69.76129, 69.79808, 
    69.83449, 69.87052, 69.90617, 69.94145, 69.97634, 70.01085, 70.04497, 
    70.0787, 70.11205, 70.145, 70.17755, 70.20972, 70.24148, 70.27283, 
    70.30379, 70.33435, 70.3645, 70.39424, 70.42357, 70.45249, 70.481, 
    70.50909, 70.53676, 70.56401, 70.59084, 70.61726, 70.64324, 70.6688, 
    70.69393, 70.71864, 70.74291, 70.76675, 70.79015, 70.81312, 70.83565, 
    70.85774, 70.87939, 70.9006, 70.92136, 70.94168, 70.96156, 70.98098, 
    70.99995, 71.01848, 71.03654, 71.05416, 71.07133, 71.08804, 71.10429, 
    71.12007, 71.13541, 71.15028, 71.16468, 71.17863, 71.19211, 71.20512, 
    71.21767, 71.22976, 71.24137, 71.25252, 71.2632, 71.27341, 71.28314, 
    71.2924, 71.30119, 71.30951, 71.31735, 71.32472, 71.33161, 71.33804, 
    71.34397, 71.34944, 71.35442, 71.35894, 71.36297, 71.36652, 71.3696, 
    71.3722, 71.37431, 71.37595, 71.37711, 71.3778, 71.378, 71.37772, 
    71.37696, 71.37572, 71.37402, 71.37182, 71.36915, 71.366, 71.36237, 
    71.35825, 71.35367, 71.34861, 71.34306, 71.33705, 71.33056, 71.32359, 
    71.31615, 71.30823, 71.29984, 71.29097, 71.28163, 71.27182, 71.26154, 
    71.25079, 71.23957, 71.22788, 71.21572, 71.20309, 71.19001, 71.17645, 
    71.16244, 71.14796, 71.13301, 71.11761, 71.10175, 71.08542, 71.06864, 
    71.05141, 71.03371, 71.01557, 70.99698, 70.97794, 70.95844, 70.9385, 
    70.91811, 70.89727, 70.876, 70.85428, 70.83212, 70.80952, 70.78648, 
    70.76301, 70.7391, 70.71476, 70.68999, 70.66479, 70.63916, 70.61311, 
    70.58663, 70.55973, 70.53241, 70.50467, 70.47652, 70.44794, 70.41896, 
    70.38956, 70.35976, 70.32954, 70.29893, 70.26791, 70.23648, 70.20465, 
    70.17243, 70.13981, 70.1068, 70.07339, 70.0396, 70.00542, 69.97085, 
    69.9359, 69.90056, 69.86485, 69.82875, 69.79228, 69.75544, 69.71822, 
    69.68064, 69.64269, 69.60438, 69.5657, 69.52666, 69.48725, 69.44749, 
    69.40739, 69.36692, 69.3261, 69.28494, 69.24343, 69.20158, 69.15938, 
    69.11684, 69.07396, 69.03075, 68.98721, 68.94333, 68.89912, 68.85458, 
    68.80972, 68.76454, 68.71904, 68.67322, 68.62708, 68.58062, 68.53385, 
    68.48678, 68.43938, 68.39169, 68.3437, 68.29539, 68.2468, 68.1979, 
    68.1487, 68.09921, 68.04943, 67.99936, 67.949, 67.89835, 67.84742, 
    67.79621, 67.74472, 67.69295, 67.6409, 67.58858, 67.53599, 67.48312, 
    67.42999, 67.37659, 67.32294, 67.26901, 67.21483, 67.16039, 67.10568, 
    67.05073, 66.99552, 66.94006, 66.88435, 66.8284, 66.77219, 66.71575, 
    66.65907, 66.60213, 66.54498, 66.48757, 66.42993, 66.37206, 66.31396, 
    66.25564, 66.19707, 66.1383, 66.07928, 66.02006, 65.96061, 65.90094, 
    65.84105, 65.78094, 65.72063, 65.6601, 65.59936, 65.53841, 65.47726, 
    65.41589, 65.35432,
  59.01059, 59.08562, 59.16056, 59.23541, 59.31015, 59.3848, 59.45935, 
    59.53379, 59.60814, 59.68238, 59.75652, 59.83055, 59.90448, 59.9783, 
    60.05202, 60.12563, 60.19913, 60.27253, 60.34581, 60.41898, 60.49204, 
    60.56499, 60.63782, 60.71054, 60.78314, 60.85563, 60.928, 61.00025, 
    61.07238, 61.1444, 61.21629, 61.28806, 61.3597, 61.43122, 61.50262, 
    61.57389, 61.64503, 61.71604, 61.78693, 61.85768, 61.9283, 61.99879, 
    62.06915, 62.13937, 62.20946, 62.27941, 62.34922, 62.41889, 62.48842, 
    62.55781, 62.62706, 62.69616, 62.76512, 62.83393, 62.9026, 62.97112, 
    63.03949, 63.10771, 63.17577, 63.24368, 63.31144, 63.37904, 63.44649, 
    63.51377, 63.5809, 63.64787, 63.71467, 63.78131, 63.84779, 63.9141, 
    63.98024, 64.04622, 64.11202, 64.17765, 64.24311, 64.3084, 64.3735, 
    64.43844, 64.5032, 64.56777, 64.63216, 64.69637, 64.7604, 64.82424, 
    64.88789, 64.95135, 65.01463, 65.07771, 65.1406, 65.2033, 65.26579, 
    65.32809, 65.3902, 65.4521, 65.51379, 65.57529, 65.63657, 65.69765, 
    65.75853, 65.81919, 65.87964, 65.93987, 65.99989, 66.05969, 66.11928, 
    66.17863, 66.23778, 66.29669, 66.35538, 66.41384, 66.47208, 66.53008, 
    66.58784, 66.64538, 66.70267, 66.75974, 66.81655, 66.87313, 66.92947, 
    66.98555, 67.04139, 67.09698, 67.15232, 67.20741, 67.26225, 67.31682, 
    67.37113, 67.42519, 67.47898, 67.53251, 67.58577, 67.63876, 67.69148, 
    67.74393, 67.79611, 67.84801, 67.89963, 67.95097, 68.00203, 68.0528, 
    68.10329, 68.15349, 68.20339, 68.25301, 68.30233, 68.35136, 68.40008, 
    68.4485, 68.49663, 68.54444, 68.59195, 68.63915, 68.68604, 68.73261, 
    68.77888, 68.82482, 68.87044, 68.91574, 68.96072, 69.00537, 69.04969, 
    69.09368, 69.13734, 69.18066, 69.22366, 69.2663, 69.30861, 69.35058, 
    69.3922, 69.43347, 69.47439, 69.51496, 69.55518, 69.59504, 69.63454, 
    69.67368, 69.71246, 69.75088, 69.78893, 69.82661, 69.86392, 69.90086, 
    69.93742, 69.9736, 70.00941, 70.04483, 70.07987, 70.11452, 70.1488, 
    70.18267, 70.21616, 70.24925, 70.28195, 70.31425, 70.34615, 70.37765, 
    70.40874, 70.43944, 70.46972, 70.49959, 70.52905, 70.55811, 70.58674, 
    70.61495, 70.64275, 70.67013, 70.69708, 70.72362, 70.74972, 70.7754, 
    70.80064, 70.82546, 70.84985, 70.87379, 70.89731, 70.92039, 70.94302, 
    70.96522, 70.98697, 71.00828, 71.02914, 71.04955, 71.06952, 71.08904, 
    71.1081, 71.12672, 71.14487, 71.16257, 71.17982, 71.19661, 71.21294, 
    71.22881, 71.24421, 71.25915, 71.27363, 71.28764, 71.30119, 71.31427, 
    71.32688, 71.33903, 71.35069, 71.3619, 71.37263, 71.38288, 71.39267, 
    71.40198, 71.41081, 71.41917, 71.42705, 71.43446, 71.44138, 71.44783, 
    71.4538, 71.4593, 71.46431, 71.46884, 71.47289, 71.47646, 71.47956, 
    71.48217, 71.4843, 71.48595, 71.48711, 71.48779, 71.488, 71.48772, 
    71.48696, 71.48572, 71.48399, 71.48179, 71.4791, 71.47594, 71.47228, 
    71.46815, 71.46355, 71.45846, 71.45289, 71.44685, 71.44032, 71.43332, 
    71.42583, 71.41788, 71.40945, 71.40054, 71.39115, 71.38129, 71.37096, 
    71.36016, 71.34888, 71.33714, 71.32492, 71.31223, 71.29908, 71.28545, 
    71.27137, 71.25682, 71.2418, 71.22633, 71.21038, 71.19398, 71.17712, 
    71.15981, 71.14203, 71.1238, 71.10512, 71.08598, 71.06639, 71.04636, 
    71.02587, 71.00494, 70.98356, 70.96173, 70.93947, 70.91676, 70.89362, 
    70.87004, 70.84602, 70.82156, 70.79668, 70.77136, 70.74562, 70.71944, 
    70.69285, 70.66582, 70.63838, 70.61052, 70.58224, 70.55354, 70.52442, 
    70.4949, 70.46496, 70.43461, 70.40385, 70.3727, 70.34113, 70.30917, 
    70.2768, 70.24404, 70.21089, 70.17734, 70.1434, 70.10907, 70.07436, 
    70.03925, 70.00377, 69.9679, 69.93166, 69.89503, 69.85804, 69.82067, 
    69.78294, 69.74483, 69.70635, 69.66752, 69.62832, 69.58876, 69.54884, 
    69.50857, 69.46794, 69.42696, 69.38564, 69.34396, 69.30194, 69.25958, 
    69.21688, 69.17384, 69.13046, 69.08675, 69.0427, 68.99833, 68.95363, 
    68.9086, 68.86324, 68.81757, 68.77158, 68.72527, 68.67864, 68.63171, 
    68.58446, 68.5369, 68.48904, 68.44086, 68.3924, 68.34362, 68.29455, 
    68.24518, 68.19552, 68.14557, 68.09532, 68.04479, 67.99397, 67.94287, 
    67.89148, 67.83982, 67.78787, 67.73566, 67.68316, 67.63039, 67.57736, 
    67.52406, 67.47049, 67.41666, 67.36256, 67.3082, 67.25359, 67.19872, 
    67.14359, 67.0882, 67.03258, 66.9767, 66.92057, 66.8642, 66.80759, 
    66.75072, 66.69363, 66.63629, 66.57872, 66.52092, 66.46288, 66.40461, 
    66.34612, 66.28738, 66.22844, 66.16927, 66.10986, 66.05025, 65.99041, 
    65.93036, 65.87009, 65.80961, 65.74892, 65.68801, 65.6269, 65.56557, 
    65.50405, 65.44232,
  59.08569, 59.16083, 59.23589, 59.31084, 59.3857, 59.46045, 59.53511, 
    59.60967, 59.68413, 59.75848, 59.83274, 59.90689, 59.98093, 60.05487, 
    60.12871, 60.20244, 60.27606, 60.34957, 60.42297, 60.49627, 60.56945, 
    60.64252, 60.71547, 60.78831, 60.86104, 60.93365, 61.00615, 61.07853, 
    61.15078, 61.22292, 61.29494, 61.36683, 61.43861, 61.51026, 61.58178, 
    61.65318, 61.72446, 61.7956, 61.86662, 61.9375, 62.00826, 62.07888, 
    62.14938, 62.21973, 62.28996, 62.36004, 62.42999, 62.4998, 62.56947, 
    62.639, 62.70838, 62.77763, 62.84673, 62.91568, 62.98449, 63.05315, 
    63.12166, 63.19002, 63.25823, 63.32629, 63.39419, 63.46194, 63.52953, 
    63.59697, 63.66424, 63.73135, 63.79831, 63.8651, 63.93172, 63.99818, 
    64.06448, 64.13061, 64.19656, 64.26234, 64.32796, 64.39339, 64.45866, 
    64.52375, 64.58866, 64.65339, 64.71794, 64.7823, 64.84649, 64.91048, 
    64.9743, 65.03793, 65.10136, 65.1646, 65.22765, 65.2905, 65.35316, 
    65.41563, 65.47789, 65.53996, 65.60181, 65.66348, 65.72492, 65.78617, 
    65.84721, 65.90803, 65.96864, 66.02905, 66.08923, 66.1492, 66.20895, 
    66.26848, 66.32779, 66.38687, 66.44573, 66.50436, 66.56276, 66.62093, 
    66.67887, 66.73658, 66.79404, 66.85127, 66.90826, 66.96501, 67.02151, 
    67.07777, 67.13379, 67.18955, 67.24506, 67.30032, 67.35533, 67.41008, 
    67.46457, 67.51879, 67.57276, 67.62646, 67.67989, 67.73306, 67.78596, 
    67.83858, 67.89093, 67.94301, 67.9948, 68.04631, 68.09754, 68.14849, 
    68.19915, 68.24953, 68.29961, 68.3494, 68.39889, 68.44809, 68.49699, 
    68.54559, 68.59388, 68.64187, 68.68954, 68.73692, 68.78398, 68.83073, 
    68.87716, 68.92327, 68.96906, 69.01453, 69.05968, 69.1045, 69.14899, 
    69.19315, 69.23698, 69.28047, 69.32362, 69.36644, 69.40891, 69.45104, 
    69.49283, 69.53426, 69.57535, 69.61608, 69.65646, 69.69649, 69.73615, 
    69.77545, 69.81438, 69.85296, 69.89117, 69.929, 69.96647, 70.00356, 
    70.04028, 70.07661, 70.11257, 70.14815, 70.18333, 70.21814, 70.25256, 
    70.28658, 70.32021, 70.35345, 70.38628, 70.41873, 70.45077, 70.48241, 
    70.51364, 70.54446, 70.57488, 70.60489, 70.63448, 70.66367, 70.69243, 
    70.72077, 70.7487, 70.7762, 70.80328, 70.82993, 70.85616, 70.88196, 
    70.90733, 70.93225, 70.95675, 70.98081, 71.00444, 71.02762, 71.05036, 
    71.07266, 71.09452, 71.11593, 71.13689, 71.1574, 71.17747, 71.19707, 
    71.21623, 71.23493, 71.25318, 71.27097, 71.2883, 71.30517, 71.32157, 
    71.33752, 71.353, 71.36801, 71.38256, 71.39664, 71.41026, 71.4234, 
    71.43608, 71.44828, 71.46001, 71.47127, 71.48205, 71.49236, 71.50219, 
    71.51154, 71.52042, 71.52882, 71.53674, 71.54419, 71.55115, 71.55763, 
    71.56363, 71.56915, 71.57419, 71.57874, 71.58282, 71.58641, 71.58952, 
    71.59214, 71.59428, 71.59593, 71.59711, 71.59779, 71.598, 71.59772, 
    71.59695, 71.5957, 71.59397, 71.59176, 71.58906, 71.58588, 71.58221, 
    71.57806, 71.57343, 71.56831, 71.56271, 71.55664, 71.55008, 71.54305, 
    71.53552, 71.52753, 71.51905, 71.51009, 71.50066, 71.49076, 71.48038, 
    71.46952, 71.45818, 71.44638, 71.4341, 71.42136, 71.40813, 71.39445, 
    71.38029, 71.36567, 71.35058, 71.33502, 71.31901, 71.30253, 71.28558, 
    71.26818, 71.25032, 71.232, 71.21323, 71.194, 71.17432, 71.15419, 
    71.13361, 71.11257, 71.09109, 71.06917, 71.0468, 71.02398, 71.00073, 
    70.97704, 70.9529, 70.92834, 70.90334, 70.87791, 70.85204, 70.82574, 
    70.79903, 70.77188, 70.74431, 70.71632, 70.68791, 70.65908, 70.62984, 
    70.60017, 70.5701, 70.53962, 70.50873, 70.47743, 70.44572, 70.41363, 
    70.38112, 70.34821, 70.31492, 70.28122, 70.24713, 70.21266, 70.1778, 
    70.14254, 70.10691, 70.07089, 70.03449, 69.99772, 69.96057, 69.92304, 
    69.88515, 69.84689, 69.80825, 69.76926, 69.7299, 69.69018, 69.6501, 
    69.60966, 69.56887, 69.52773, 69.48624, 69.4444, 69.40222, 69.35969, 
    69.31682, 69.27361, 69.23006, 69.18619, 69.14198, 69.09743, 69.05256, 
    69.00736, 68.96184, 68.916, 68.86983, 68.82335, 68.77656, 68.72945, 
    68.68202, 68.63429, 68.58626, 68.53792, 68.48927, 68.44032, 68.39108, 
    68.34154, 68.2917, 68.24158, 68.19116, 68.14045, 68.08946, 68.03819, 
    67.98663, 67.93478, 67.88267, 67.83028, 67.77761, 67.72467, 67.67146, 
    67.61798, 67.56424, 67.51023, 67.45596, 67.40144, 67.34664, 67.2916, 
    67.2363, 67.18075, 67.12495, 67.06889, 67.0126, 66.95605, 66.89927, 
    66.84224, 66.78497, 66.72746, 66.66972, 66.61175, 66.55354, 66.4951, 
    66.43643, 66.37754, 66.31842, 66.25908, 66.19952, 66.13973, 66.07973, 
    66.01951, 65.95907, 65.89842, 65.83756, 65.7765, 65.71522, 65.65373, 
    65.59204, 65.53015,
  59.16059, 59.23585, 59.31101, 59.38608, 59.46105, 59.53592, 59.61069, 
    59.68536, 59.75993, 59.8344, 59.90877, 59.98304, 60.0572, 60.13126, 
    60.20521, 60.27906, 60.35279, 60.42643, 60.49995, 60.57336, 60.64666, 
    60.71986, 60.79293, 60.8659, 60.93875, 61.01149, 61.0841, 61.1566, 
    61.22899, 61.30125, 61.3734, 61.44542, 61.51733, 61.58911, 61.66076, 
    61.73229, 61.8037, 61.87497, 61.94612, 62.01714, 62.08803, 62.15879, 
    62.22941, 62.2999, 62.37026, 62.44049, 62.51057, 62.58052, 62.65033, 
    62.71999, 62.78952, 62.85891, 62.92815, 62.99724, 63.06619, 63.13499, 
    63.20365, 63.27216, 63.34051, 63.40871, 63.47676, 63.54465, 63.61239, 
    63.67997, 63.74739, 63.81466, 63.88176, 63.9487, 64.01548, 64.08209, 
    64.14854, 64.21481, 64.28092, 64.34686, 64.41263, 64.47822, 64.54364, 
    64.60888, 64.67394, 64.73883, 64.80354, 64.86806, 64.9324, 64.99656, 
    65.06053, 65.12431, 65.18791, 65.25131, 65.31452, 65.37754, 65.44036, 
    65.50299, 65.56541, 65.62764, 65.68967, 65.75149, 65.8131, 65.87451, 
    65.93571, 65.99671, 66.05749, 66.11806, 66.17841, 66.23855, 66.29846, 
    66.35816, 66.41764, 66.47689, 66.53592, 66.59472, 66.65329, 66.71163, 
    66.76974, 66.82762, 66.88526, 66.94266, 66.99982, 67.05674, 67.11342, 
    67.16985, 67.22604, 67.28197, 67.33766, 67.3931, 67.44827, 67.5032, 
    67.55785, 67.61226, 67.6664, 67.72028, 67.77389, 67.82722, 67.88029, 
    67.9331, 67.98562, 68.03786, 68.08984, 68.14153, 68.19293, 68.24406, 
    68.29489, 68.34544, 68.39569, 68.44566, 68.49532, 68.5447, 68.59377, 
    68.64254, 68.69101, 68.73917, 68.78703, 68.83457, 68.88181, 68.92873, 
    68.97533, 69.02161, 69.06757, 69.11322, 69.15854, 69.20353, 69.24818, 
    69.29252, 69.33652, 69.38017, 69.4235, 69.46648, 69.50912, 69.55141, 
    69.59337, 69.63497, 69.67622, 69.71712, 69.75766, 69.79784, 69.83767, 
    69.87713, 69.91623, 69.95496, 69.99332, 70.03132, 70.06895, 70.10619, 
    70.14306, 70.17955, 70.21566, 70.25139, 70.28673, 70.32169, 70.35625, 
    70.39042, 70.42419, 70.45758, 70.49056, 70.52315, 70.55533, 70.58711, 
    70.61848, 70.64944, 70.68, 70.71014, 70.73987, 70.76918, 70.79808, 
    70.82655, 70.85461, 70.88223, 70.90944, 70.93621, 70.96256, 70.98848, 
    71.01396, 71.03901, 71.06362, 71.0878, 71.11153, 71.13483, 71.15768, 
    71.18008, 71.20204, 71.22356, 71.24461, 71.26523, 71.28539, 71.30509, 
    71.32434, 71.34313, 71.36147, 71.37934, 71.39675, 71.4137, 71.43019, 
    71.44622, 71.46178, 71.47686, 71.49149, 71.50564, 71.51932, 71.53252, 
    71.54527, 71.55753, 71.56931, 71.58063, 71.59147, 71.60183, 71.61171, 
    71.62111, 71.63004, 71.63847, 71.64644, 71.65392, 71.66091, 71.66743, 
    71.67346, 71.67901, 71.68407, 71.68865, 71.69274, 71.69635, 71.69947, 
    71.70211, 71.70426, 71.70592, 71.7071, 71.70779, 71.708, 71.70772, 
    71.70695, 71.7057, 71.70395, 71.70172, 71.69901, 71.69581, 71.69212, 
    71.68796, 71.6833, 71.67816, 71.67254, 71.66643, 71.65984, 71.65276, 
    71.64521, 71.63717, 71.62865, 71.61965, 71.61018, 71.60022, 71.58978, 
    71.57887, 71.56748, 71.55562, 71.54328, 71.53047, 71.51719, 71.50343, 
    71.4892, 71.47451, 71.45934, 71.44371, 71.42762, 71.41106, 71.39403, 
    71.37654, 71.3586, 71.34019, 71.32133, 71.302, 71.28223, 71.26199, 
    71.24131, 71.22018, 71.1986, 71.17657, 71.15409, 71.13117, 71.1078, 
    71.084, 71.05976, 71.03508, 71.00996, 70.98441, 70.95842, 70.93201, 
    70.90517, 70.87789, 70.8502, 70.82207, 70.79353, 70.76457, 70.7352, 
    70.70541, 70.67519, 70.64458, 70.61355, 70.58211, 70.55027, 70.51802, 
    70.48537, 70.45232, 70.41888, 70.38504, 70.35081, 70.31618, 70.28117, 
    70.24577, 70.20998, 70.17381, 70.13725, 70.10033, 70.06302, 70.02534, 
    69.98728, 69.94886, 69.91007, 69.87091, 69.83139, 69.79151, 69.75127, 
    69.71067, 69.66972, 69.62841, 69.58675, 69.54475, 69.5024, 69.4597, 
    69.41666, 69.37329, 69.32957, 69.28553, 69.24114, 69.19643, 69.15139, 
    69.10602, 69.06033, 69.01431, 68.96798, 68.92133, 68.87435, 68.82707, 
    68.77948, 68.73158, 68.68336, 68.63485, 68.58603, 68.53691, 68.48749, 
    68.43777, 68.38776, 68.33746, 68.28687, 68.23598, 68.18482, 68.13337, 
    68.08163, 68.02962, 67.97733, 67.92476, 67.87192, 67.81881, 67.76542, 
    67.71177, 67.65785, 67.60367, 67.54922, 67.49452, 67.43956, 67.38434, 
    67.32887, 67.27314, 67.21717, 67.16094, 67.10447, 67.04775, 66.9908, 
    66.93359, 66.87616, 66.81848, 66.76057, 66.70242, 66.64404, 66.58543, 
    66.5266, 66.46754, 66.40825, 66.34873, 66.289, 66.22905, 66.16888, 
    66.10849, 66.04789, 65.98708, 65.92605, 65.86481, 65.80337, 65.74172, 
    65.67987, 65.61781,
  59.23532, 59.31068, 59.38595, 59.46113, 59.53621, 59.61119, 59.68607, 
    59.76086, 59.83554, 59.91013, 59.98462, 60.05899, 60.13327, 60.20745, 
    60.28152, 60.35548, 60.42934, 60.50309, 60.57673, 60.65027, 60.72369, 
    60.797, 60.8702, 60.94329, 61.01627, 61.08913, 61.16187, 61.2345, 
    61.30701, 61.3794, 61.45167, 61.52382, 61.59586, 61.66776, 61.73955, 
    61.81121, 61.88274, 61.95415, 62.02543, 62.09659, 62.16761, 62.2385, 
    62.30926, 62.37989, 62.45038, 62.52074, 62.59097, 62.66105, 62.731, 
    62.8008, 62.87047, 62.93999, 63.00938, 63.07862, 63.14771, 63.21665, 
    63.28545, 63.3541, 63.4226, 63.49095, 63.55914, 63.62718, 63.69507, 
    63.76279, 63.83037, 63.89778, 63.96503, 64.03212, 64.09904, 64.16581, 
    64.23241, 64.29884, 64.3651, 64.43119, 64.49711, 64.56286, 64.62843, 
    64.69383, 64.75906, 64.8241, 64.88896, 64.95364, 65.01814, 65.08246, 
    65.14659, 65.21053, 65.27428, 65.33785, 65.40122, 65.4644, 65.52739, 
    65.59018, 65.65276, 65.71516, 65.77734, 65.83933, 65.90112, 65.96269, 
    66.02406, 66.08522, 66.14616, 66.2069, 66.26743, 66.32773, 66.38782, 
    66.44769, 66.50733, 66.56675, 66.62595, 66.68492, 66.74367, 66.80218, 
    66.86046, 66.9185, 66.97632, 67.03389, 67.09122, 67.14832, 67.20517, 
    67.26178, 67.31814, 67.37424, 67.43011, 67.48572, 67.54107, 67.59617, 
    67.651, 67.70558, 67.7599, 67.81395, 67.86774, 67.92125, 67.97449, 
    68.02747, 68.08017, 68.1326, 68.18475, 68.23661, 68.28819, 68.33949, 
    68.3905, 68.44122, 68.49165, 68.54179, 68.59164, 68.64118, 68.69043, 
    68.73938, 68.78802, 68.83636, 68.88439, 68.93211, 68.97952, 69.02661, 
    69.07339, 69.11984, 69.16599, 69.21179, 69.25729, 69.30244, 69.34728, 
    69.39178, 69.43594, 69.47977, 69.52327, 69.56642, 69.60923, 69.6517, 
    69.69381, 69.73558, 69.777, 69.81806, 69.85876, 69.89912, 69.9391, 
    69.97873, 70.01799, 70.05688, 70.09541, 70.13356, 70.17134, 70.20875, 
    70.24577, 70.28242, 70.31868, 70.35456, 70.39005, 70.42516, 70.45988, 
    70.49419, 70.52812, 70.56165, 70.59478, 70.62751, 70.65984, 70.69176, 
    70.72327, 70.75437, 70.78506, 70.81535, 70.84521, 70.87465, 70.90368, 
    70.93228, 70.96046, 70.98822, 71.01555, 71.04245, 71.06892, 71.09496, 
    71.12056, 71.14573, 71.17046, 71.19475, 71.2186, 71.242, 71.26496, 
    71.28748, 71.30954, 71.33115, 71.35232, 71.37302, 71.39328, 71.41309, 
    71.43243, 71.45131, 71.46973, 71.48769, 71.5052, 71.52223, 71.5388, 
    71.5549, 71.57053, 71.5857, 71.6004, 71.61462, 71.62836, 71.64164, 
    71.65444, 71.66677, 71.67861, 71.68999, 71.70087, 71.71129, 71.72122, 
    71.73067, 71.73964, 71.74812, 71.75613, 71.76364, 71.77068, 71.77722, 
    71.78328, 71.78886, 71.79395, 71.79855, 71.80267, 71.80629, 71.80943, 
    71.81208, 71.81424, 71.81591, 71.8171, 71.81779, 71.818, 71.81772, 
    71.81694, 71.81568, 71.81393, 71.81169, 71.80897, 71.80575, 71.80205, 
    71.79785, 71.79317, 71.78801, 71.78236, 71.77621, 71.76959, 71.76248, 
    71.75489, 71.74681, 71.73825, 71.7292, 71.71968, 71.70967, 71.69919, 
    71.68822, 71.67677, 71.66485, 71.65245, 71.63957, 71.62622, 71.6124, 
    71.5981, 71.58334, 71.56809, 71.55238, 71.53621, 71.51957, 71.50246, 
    71.48489, 71.46685, 71.44836, 71.4294, 71.40998, 71.39011, 71.36978, 
    71.349, 71.32777, 71.30608, 71.28394, 71.26136, 71.23833, 71.21485, 
    71.19093, 71.16657, 71.14178, 71.11654, 71.09087, 71.06477, 71.03822, 
    71.01126, 70.98386, 70.95604, 70.92779, 70.89912, 70.87003, 70.84051, 
    70.81059, 70.78024, 70.74948, 70.71832, 70.68674, 70.65475, 70.62236, 
    70.58957, 70.55637, 70.52278, 70.48879, 70.45441, 70.41963, 70.38447, 
    70.34892, 70.31297, 70.27665, 70.23994, 70.20285, 70.16539, 70.12755, 
    70.08934, 70.05075, 70.0118, 69.97248, 69.9328, 69.89275, 69.85235, 
    69.81158, 69.77047, 69.729, 69.68717, 69.645, 69.60249, 69.55962, 
    69.51641, 69.47287, 69.42899, 69.38477, 69.34021, 69.29533, 69.25011, 
    69.20457, 69.15871, 69.11252, 69.06601, 69.01918, 68.97204, 68.92458, 
    68.87681, 68.82874, 68.78035, 68.73166, 68.68266, 68.63337, 68.58377, 
    68.53388, 68.4837, 68.43322, 68.38245, 68.33139, 68.28005, 68.22842, 
    68.17651, 68.12432, 68.07185, 68.01911, 67.96609, 67.9128, 67.85925, 
    67.80542, 67.75132, 67.69697, 67.64235, 67.58746, 67.53233, 67.47694, 
    67.42129, 67.36539, 67.30924, 67.25284, 67.1962, 67.13931, 67.08218, 
    67.0248, 66.96719, 66.90934, 66.85126, 66.79294, 66.73439, 66.67561, 
    66.6166, 66.55737, 66.49791, 66.43822, 66.37833, 66.31821, 66.25787, 
    66.19731, 66.13654, 66.07556, 66.01437, 65.95296, 65.89136, 65.82954, 
    65.76752, 65.7053,
  59.30984, 59.38532, 59.4607, 59.53599, 59.61118, 59.68627, 59.76127, 
    59.83617, 59.91097, 59.98567, 60.06026, 60.13476, 60.20916, 60.28345, 
    60.35764, 60.43172, 60.5057, 60.57956, 60.65333, 60.72698, 60.80053, 
    60.87396, 60.94728, 61.02049, 61.09359, 61.16658, 61.23944, 61.3122, 
    61.38483, 61.45735, 61.52975, 61.60203, 61.67419, 61.74623, 61.81815, 
    61.88993, 61.9616, 62.03314, 62.10456, 62.17584, 62.247, 62.31802, 
    62.38892, 62.45968, 62.53031, 62.60081, 62.67117, 62.74139, 62.81148, 
    62.88142, 62.95123, 63.0209, 63.09042, 63.1598, 63.22903, 63.29812, 
    63.36707, 63.43586, 63.5045, 63.57299, 63.64133, 63.70952, 63.77756, 
    63.84543, 63.91315, 63.98071, 64.04812, 64.11536, 64.18243, 64.24935, 
    64.31609, 64.38268, 64.4491, 64.51534, 64.58141, 64.64732, 64.71305, 
    64.7786, 64.84398, 64.90918, 64.97421, 65.03905, 65.10371, 65.16818, 
    65.23247, 65.29658, 65.36049, 65.42422, 65.48775, 65.55109, 65.61424, 
    65.67719, 65.73994, 65.8025, 65.86485, 65.92701, 65.98895, 66.0507, 
    66.11224, 66.17356, 66.23468, 66.29558, 66.35627, 66.41674, 66.477, 
    66.53704, 66.59686, 66.65645, 66.71582, 66.77496, 66.83388, 66.89256, 
    66.95101, 67.00923, 67.06722, 67.12497, 67.18248, 67.23975, 67.29677, 
    67.35355, 67.41009, 67.46637, 67.52241, 67.57819, 67.63372, 67.68899, 
    67.744, 67.79876, 67.85325, 67.90748, 67.96144, 68.01514, 68.06856, 
    68.12171, 68.17458, 68.22719, 68.27951, 68.33155, 68.38332, 68.43479, 
    68.48598, 68.53688, 68.58749, 68.6378, 68.68782, 68.73755, 68.78697, 
    68.8361, 68.88491, 68.93343, 68.98163, 69.02953, 69.07711, 69.12438, 
    69.17133, 69.21796, 69.26427, 69.31026, 69.35593, 69.40126, 69.44627, 
    69.49094, 69.53528, 69.57928, 69.62294, 69.66627, 69.70924, 69.75188, 
    69.79416, 69.8361, 69.87769, 69.91891, 69.95979, 70.0003, 70.04045, 
    70.08024, 70.11966, 70.15872, 70.1974, 70.23572, 70.27366, 70.31122, 
    70.3484, 70.38521, 70.42163, 70.45766, 70.49331, 70.52856, 70.56343, 
    70.59791, 70.63198, 70.66566, 70.69894, 70.73181, 70.76428, 70.79634, 
    70.828, 70.85925, 70.89008, 70.92049, 70.95049, 70.98007, 71.00923, 
    71.03797, 71.06628, 71.09417, 71.12162, 71.14865, 71.17525, 71.2014, 
    71.22713, 71.25241, 71.27726, 71.30167, 71.32562, 71.34914, 71.37221, 
    71.39484, 71.41701, 71.43872, 71.45999, 71.4808, 71.50116, 71.52106, 
    71.54049, 71.55947, 71.57798, 71.59603, 71.61362, 71.63074, 71.64739, 
    71.66357, 71.67928, 71.69453, 71.70929, 71.72359, 71.7374, 71.75075, 
    71.76361, 71.776, 71.7879, 71.79933, 71.81028, 71.82074, 71.83073, 
    71.84023, 71.84924, 71.85777, 71.86581, 71.87336, 71.88043, 71.88701, 
    71.8931, 71.89871, 71.90382, 71.90845, 71.91258, 71.91623, 71.91939, 
    71.92205, 71.92422, 71.9259, 71.92709, 71.92779, 71.928, 71.92771, 
    71.92694, 71.92567, 71.92391, 71.92166, 71.91892, 71.91569, 71.91196, 
    71.90775, 71.90305, 71.89786, 71.89217, 71.886, 71.87935, 71.8722, 
    71.86456, 71.85645, 71.84784, 71.83875, 71.82918, 71.81912, 71.80858, 
    71.79755, 71.78606, 71.77407, 71.7616, 71.74866, 71.73525, 71.72136, 
    71.70699, 71.69215, 71.67683, 71.66104, 71.64479, 71.62806, 71.61087, 
    71.59321, 71.57509, 71.5565, 71.53745, 71.51794, 71.49797, 71.47754, 
    71.45666, 71.43532, 71.41353, 71.39128, 71.36859, 71.34545, 71.32186, 
    71.29784, 71.27336, 71.24844, 71.22308, 71.1973, 71.17107, 71.1444, 
    71.11731, 71.08978, 71.06183, 71.03345, 71.00465, 70.97542, 70.94577, 
    70.91571, 70.88522, 70.85433, 70.82302, 70.7913, 70.75917, 70.72664, 
    70.6937, 70.66035, 70.62662, 70.59248, 70.55795, 70.52302, 70.4877, 
    70.45199, 70.41589, 70.37941, 70.34255, 70.30531, 70.26768, 70.22968, 
    70.19131, 70.15257, 70.11345, 70.07397, 70.03413, 69.99391, 69.95334, 
    69.91241, 69.87112, 69.82949, 69.7875, 69.74516, 69.70247, 69.65943, 
    69.61606, 69.57234, 69.52828, 69.48389, 69.43917, 69.39411, 69.34872, 
    69.30301, 69.25697, 69.21061, 69.16393, 69.11692, 69.0696, 69.02197, 
    68.97403, 68.92577, 68.87721, 68.82835, 68.77917, 68.7297, 68.67993, 
    68.62986, 68.5795, 68.52885, 68.4779, 68.42667, 68.37514, 68.32334, 
    68.27126, 68.21889, 68.16624, 68.11332, 68.06013, 68.00666, 67.95292, 
    67.89892, 67.84465, 67.79012, 67.73532, 67.68027, 67.62495, 67.56938, 
    67.51356, 67.45748, 67.40116, 67.34458, 67.28777, 67.23071, 67.17339, 
    67.11585, 67.05807, 67.00004, 66.94179, 66.88329, 66.82457, 66.76562, 
    66.70644, 66.64703, 66.58741, 66.52756, 66.46748, 66.4072, 66.34669, 
    66.28596, 66.22502, 66.16387, 66.10252, 66.04095, 65.97917, 65.91719, 
    65.855, 65.79262,
  59.38418, 59.45977, 59.53526, 59.61065, 59.68596, 59.76116, 59.83627, 
    59.91128, 59.98619, 60.06101, 60.13572, 60.21033, 60.28484, 60.35925, 
    60.43356, 60.50776, 60.58186, 60.65584, 60.72972, 60.8035, 60.87717, 
    60.95072, 61.02417, 61.0975, 61.17072, 61.24383, 61.31683, 61.3897, 
    61.46247, 61.53511, 61.60764, 61.68005, 61.75233, 61.8245, 61.89655, 
    61.96847, 62.04026, 62.11194, 62.18348, 62.2549, 62.32619, 62.39735, 
    62.46838, 62.53928, 62.61005, 62.68068, 62.75118, 62.82154, 62.89177, 
    62.96185, 63.0318, 63.10161, 63.17127, 63.2408, 63.31017, 63.3794, 
    63.44849, 63.51743, 63.58622, 63.65485, 63.72334, 63.79168, 63.85986, 
    63.92788, 63.99575, 64.06346, 64.13101, 64.1984, 64.26563, 64.3327, 
    64.3996, 64.46634, 64.53291, 64.5993, 64.66553, 64.7316, 64.79748, 
    64.86319, 64.92873, 64.99409, 65.05927, 65.12427, 65.18909, 65.25372, 
    65.31817, 65.38244, 65.44651, 65.5104, 65.5741, 65.6376, 65.70091, 
    65.76403, 65.82695, 65.88967, 65.95219, 66.01451, 66.07662, 66.13853, 
    66.20024, 66.26173, 66.32302, 66.38409, 66.44495, 66.50559, 66.56602, 
    66.62623, 66.68622, 66.74598, 66.80552, 66.86484, 66.92393, 66.98278, 
    67.04141, 67.09981, 67.15797, 67.21589, 67.27357, 67.33101, 67.38821, 
    67.44517, 67.50188, 67.55834, 67.61455, 67.67051, 67.72622, 67.78167, 
    67.83686, 67.89179, 67.94646, 68.00086, 68.055, 68.10888, 68.16248, 
    68.21581, 68.26886, 68.32164, 68.37415, 68.42636, 68.4783, 68.52995, 
    68.58132, 68.6324, 68.68319, 68.73368, 68.78388, 68.83378, 68.88338, 
    68.93269, 68.98168, 69.03037, 69.07876, 69.12682, 69.17458, 69.22203, 
    69.26916, 69.31596, 69.36246, 69.40862, 69.45445, 69.49996, 69.54514, 
    69.58999, 69.6345, 69.67868, 69.72251, 69.76601, 69.80916, 69.85196, 
    69.89442, 69.93652, 69.97827, 70.01967, 70.06071, 70.10139, 70.14171, 
    70.18166, 70.22125, 70.26048, 70.29932, 70.3378, 70.3759, 70.41362, 
    70.45097, 70.48792, 70.5245, 70.56069, 70.5965, 70.6319, 70.66692, 
    70.70155, 70.73578, 70.7696, 70.80302, 70.83605, 70.86867, 70.90087, 
    70.93267, 70.96406, 70.99503, 71.02559, 71.05573, 71.08544, 71.11473, 
    71.14361, 71.17205, 71.20007, 71.22765, 71.25481, 71.28152, 71.30781, 
    71.33366, 71.35906, 71.38403, 71.40855, 71.43262, 71.45625, 71.47943, 
    71.50217, 71.52444, 71.54626, 71.56763, 71.58855, 71.60901, 71.629, 
    71.64854, 71.6676, 71.68621, 71.70435, 71.72202, 71.73923, 71.75597, 
    71.77222, 71.78802, 71.80334, 71.81818, 71.83254, 71.84643, 71.85984, 
    71.87277, 71.88522, 71.89719, 71.90868, 71.91968, 71.93019, 71.94022, 
    71.94977, 71.95883, 71.9674, 71.97549, 71.98308, 71.99019, 71.9968, 
    72.00292, 72.00856, 72.0137, 72.01835, 72.02251, 72.02617, 72.02934, 
    72.03202, 72.0342, 72.03589, 72.03709, 72.03779, 72.038, 72.03771, 
    72.03693, 72.03566, 72.03389, 72.03162, 72.02887, 72.02562, 72.02188, 
    72.01765, 72.01292, 72.0077, 72.00199, 71.99579, 71.9891, 71.98191, 
    71.97424, 71.96608, 71.95743, 71.9483, 71.93867, 71.92856, 71.91797, 
    71.90689, 71.89532, 71.88328, 71.87076, 71.85775, 71.84426, 71.8303, 
    71.81586, 71.80094, 71.78555, 71.76968, 71.75335, 71.73654, 71.71926, 
    71.70152, 71.6833, 71.66462, 71.64548, 71.62587, 71.6058, 71.58527, 
    71.56429, 71.54285, 71.52095, 71.4986, 71.47579, 71.45255, 71.42884, 
    71.40469, 71.3801, 71.35507, 71.3296, 71.30368, 71.27733, 71.25053, 
    71.22331, 71.19566, 71.16758, 71.13907, 71.11013, 71.08076, 71.05099, 
    71.02078, 70.99016, 70.95912, 70.92767, 70.89581, 70.86353, 70.83086, 
    70.79777, 70.76428, 70.73038, 70.6961, 70.66142, 70.62634, 70.59086, 
    70.55499, 70.51875, 70.4821, 70.44508, 70.40768, 70.3699, 70.33173, 
    70.2932, 70.2543, 70.21501, 70.17537, 70.13535, 70.09498, 70.05424, 
    70.01315, 69.97169, 69.92989, 69.88773, 69.84521, 69.80235, 69.75915, 
    69.7156, 69.67171, 69.62749, 69.58292, 69.53802, 69.49279, 69.44723, 
    69.40134, 69.35513, 69.30859, 69.26173, 69.21455, 69.16705, 69.11924, 
    69.07112, 69.02269, 68.97395, 68.9249, 68.87556, 68.8259, 68.77596, 
    68.72572, 68.67517, 68.62434, 68.57322, 68.5218, 68.47011, 68.41812, 
    68.36586, 68.31331, 68.26049, 68.20739, 68.15401, 68.10037, 68.04646, 
    67.99228, 67.93783, 67.88312, 67.82815, 67.77291, 67.71742, 67.66167, 
    67.60567, 67.54942, 67.49293, 67.43617, 67.37918, 67.32195, 67.26446, 
    67.20674, 67.14878, 67.09058, 67.03215, 66.97349, 66.9146, 66.85547, 
    66.79612, 66.73654, 66.67674, 66.61672, 66.55647, 66.49602, 66.43533, 
    66.37444, 66.31334, 66.25202, 66.19049, 66.12875, 66.06681, 66.00467, 
    65.94231, 65.87976,
  59.45832, 59.53402, 59.60962, 59.68512, 59.76054, 59.83585, 59.91108, 
    59.9862, 60.06123, 60.13615, 60.21098, 60.28571, 60.36034, 60.43486, 
    60.50928, 60.5836, 60.65782, 60.73193, 60.80593, 60.87982, 60.95361, 
    61.02729, 61.10086, 61.17431, 61.24766, 61.32089, 61.39401, 61.46701, 
    61.5399, 61.61267, 61.68533, 61.75787, 61.83028, 61.90258, 61.97475, 
    62.04681, 62.11874, 62.19054, 62.26222, 62.33377, 62.4052, 62.47649, 
    62.54766, 62.61869, 62.68959, 62.76036, 62.831, 62.9015, 62.97186, 
    63.04209, 63.11218, 63.18213, 63.25193, 63.32159, 63.39112, 63.46049, 
    63.52972, 63.5988, 63.66774, 63.73652, 63.80516, 63.87364, 63.94197, 
    64.01014, 64.07816, 64.14602, 64.21372, 64.28127, 64.34865, 64.41586, 
    64.48292, 64.5498, 64.61653, 64.68308, 64.74947, 64.81568, 64.88173, 
    64.94759, 65.01329, 65.0788, 65.14414, 65.2093, 65.27428, 65.33908, 
    65.40369, 65.46812, 65.53236, 65.59641, 65.66027, 65.72394, 65.78741, 
    65.85069, 65.91378, 65.97666, 66.03935, 66.10184, 66.16412, 66.2262, 
    66.28807, 66.34973, 66.41119, 66.47243, 66.53345, 66.59427, 66.65487, 
    66.71525, 66.77541, 66.83535, 66.89506, 66.95455, 67.01381, 67.07285, 
    67.13165, 67.19021, 67.24854, 67.30664, 67.3645, 67.42212, 67.4795, 
    67.53663, 67.59351, 67.65015, 67.70654, 67.76268, 67.81857, 67.87419, 
    67.92956, 67.98467, 68.03952, 68.0941, 68.14842, 68.20247, 68.25626, 
    68.30976, 68.363, 68.41595, 68.46864, 68.52103, 68.57315, 68.62498, 
    68.67653, 68.72779, 68.77876, 68.82943, 68.87981, 68.92989, 68.97967, 
    69.02915, 69.07832, 69.1272, 69.17576, 69.22401, 69.27194, 69.31956, 
    69.36687, 69.41386, 69.46052, 69.50686, 69.55287, 69.59856, 69.64391, 
    69.68893, 69.73362, 69.77797, 69.82198, 69.86565, 69.90897, 69.95194, 
    69.99457, 70.03685, 70.07877, 70.12034, 70.16154, 70.20239, 70.24288, 
    70.283, 70.32275, 70.36214, 70.40115, 70.43979, 70.47806, 70.51594, 
    70.55344, 70.59056, 70.6273, 70.66365, 70.69961, 70.73518, 70.77035, 
    70.80512, 70.8395, 70.87348, 70.90706, 70.94022, 70.97299, 71.00534, 
    71.03728, 71.06882, 71.09993, 71.13062, 71.1609, 71.19076, 71.22019, 
    71.24919, 71.27777, 71.30592, 71.33363, 71.36092, 71.38776, 71.41417, 
    71.44014, 71.46567, 71.49075, 71.51539, 71.53958, 71.56333, 71.58662, 
    71.60947, 71.63185, 71.65379, 71.67525, 71.69627, 71.71683, 71.73692, 
    71.75655, 71.77572, 71.79442, 71.81265, 71.83041, 71.8477, 71.86452, 
    71.88087, 71.89674, 71.91213, 71.92705, 71.94148, 71.95544, 71.96893, 
    71.98192, 71.99443, 72.00646, 72.01801, 72.02906, 72.03963, 72.04972, 
    72.05931, 72.06842, 72.07703, 72.08516, 72.0928, 72.09994, 72.10659, 
    72.11274, 72.11841, 72.12357, 72.12825, 72.13242, 72.13611, 72.1393, 
    72.14199, 72.14418, 72.14588, 72.14709, 72.14779, 72.14799, 72.14771, 
    72.14693, 72.14565, 72.14387, 72.14159, 72.13882, 72.13556, 72.1318, 
    72.12754, 72.12279, 72.11755, 72.1118, 72.10557, 72.09884, 72.09162, 
    72.08391, 72.07571, 72.06701, 72.05783, 72.04816, 72.03799, 72.02734, 
    72.01621, 72.00459, 71.99249, 71.9799, 71.96682, 71.95327, 71.93923, 
    71.92472, 71.90973, 71.89426, 71.87831, 71.86189, 71.845, 71.82764, 
    71.8098, 71.7915, 71.77272, 71.75348, 71.73378, 71.71361, 71.69298, 
    71.67189, 71.65034, 71.62834, 71.60588, 71.58297, 71.5596, 71.53579, 
    71.51152, 71.48682, 71.46166, 71.43606, 71.41002, 71.38354, 71.35663, 
    71.32928, 71.30149, 71.27328, 71.24464, 71.21556, 71.18607, 71.15614, 
    71.1258, 71.09504, 71.06386, 71.03226, 71.00025, 70.96783, 70.93501, 
    70.90177, 70.86813, 70.83409, 70.79965, 70.76481, 70.72958, 70.69395, 
    70.65792, 70.62151, 70.58472, 70.54754, 70.50997, 70.47202, 70.4337, 
    70.395, 70.35593, 70.31649, 70.27668, 70.2365, 70.19595, 70.15505, 
    70.11378, 70.07216, 70.03018, 69.98785, 69.94517, 69.90214, 69.85876, 
    69.81504, 69.77097, 69.72658, 69.68184, 69.63676, 69.59135, 69.54562, 
    69.49955, 69.45316, 69.40645, 69.35941, 69.31205, 69.26438, 69.21639, 
    69.16809, 69.11948, 69.07056, 69.02134, 68.97182, 68.92199, 68.87186, 
    68.82143, 68.77071, 68.7197, 68.6684, 68.61681, 68.56493, 68.51276, 
    68.46032, 68.40759, 68.35459, 68.30132, 68.24776, 68.19394, 68.13985, 
    68.08549, 68.03086, 67.97597, 67.92082, 67.86541, 67.80974, 67.75381, 
    67.69764, 67.64121, 67.58453, 67.52761, 67.47044, 67.41302, 67.35536, 
    67.29747, 67.23933, 67.18096, 67.12236, 67.06352, 67.00445, 66.94515, 
    66.88563, 66.82588, 66.76591, 66.70571, 66.6453, 66.58466, 66.52382, 
    66.46275, 66.40148, 66.33999, 66.2783, 66.21639, 66.15428, 66.09196, 
    66.02945, 65.96673,
  59.53227, 59.60807, 59.68378, 59.7594, 59.83492, 59.91035, 59.98569, 
    60.06092, 60.13606, 60.21111, 60.28605, 60.36089, 60.43563, 60.51028, 
    60.58482, 60.65925, 60.73359, 60.80781, 60.88194, 60.95595, 61.02986, 
    61.10366, 61.17735, 61.25093, 61.3244, 61.39775, 61.471, 61.54413, 
    61.61714, 61.69004, 61.76283, 61.83549, 61.90804, 61.98046, 62.05276, 
    62.12495, 62.19701, 62.26894, 62.34076, 62.41244, 62.484, 62.55543, 
    62.62673, 62.6979, 62.76894, 62.83985, 62.91062, 62.98126, 63.05177, 
    63.12213, 63.19236, 63.26245, 63.3324, 63.4022, 63.47187, 63.54139, 
    63.61076, 63.67999, 63.74907, 63.818, 63.88678, 63.95541, 64.02389, 
    64.09221, 64.16038, 64.22839, 64.29624, 64.36394, 64.43147, 64.49884, 
    64.56605, 64.63309, 64.69997, 64.76668, 64.83321, 64.89959, 64.96579, 
    65.03181, 65.09766, 65.16334, 65.22884, 65.29416, 65.3593, 65.42426, 
    65.48903, 65.55362, 65.61802, 65.68224, 65.74625, 65.81009, 65.87373, 
    65.93718, 66.00043, 66.06348, 66.12634, 66.18899, 66.25143, 66.31368, 
    66.37572, 66.43756, 66.49918, 66.56059, 66.6218, 66.68278, 66.74355, 
    66.8041, 66.86443, 66.92455, 66.98443, 67.04409, 67.10353, 67.16273, 
    67.22171, 67.28046, 67.33897, 67.39724, 67.45528, 67.51307, 67.57063, 
    67.62793, 67.685, 67.74181, 67.79838, 67.8547, 67.91076, 67.96657, 
    68.02211, 68.0774, 68.13243, 68.18719, 68.24169, 68.29592, 68.34988, 
    68.40357, 68.45699, 68.51012, 68.56299, 68.61557, 68.66786, 68.71988, 
    68.77161, 68.82304, 68.87419, 68.92505, 68.9756, 69.02586, 69.07583, 
    69.12549, 69.17484, 69.22389, 69.27263, 69.32106, 69.36918, 69.41698, 
    69.46446, 69.51163, 69.55847, 69.60499, 69.65118, 69.69704, 69.74257, 
    69.78777, 69.83263, 69.87716, 69.92134, 69.96518, 70.00867, 70.05183, 
    70.09463, 70.13708, 70.17917, 70.22091, 70.26228, 70.30331, 70.34396, 
    70.38425, 70.42417, 70.46372, 70.5029, 70.5417, 70.58013, 70.61818, 
    70.65585, 70.69312, 70.73002, 70.76653, 70.80264, 70.83837, 70.8737, 
    70.90863, 70.94316, 70.97729, 71.01102, 71.04434, 71.07726, 71.10976, 
    71.14185, 71.17352, 71.20477, 71.23561, 71.26603, 71.29602, 71.32559, 
    71.35474, 71.38345, 71.41173, 71.43958, 71.46698, 71.49396, 71.52049, 
    71.54659, 71.57224, 71.59744, 71.6222, 71.64651, 71.67037, 71.69378, 
    71.71674, 71.73923, 71.76127, 71.78285, 71.80397, 71.82463, 71.84483, 
    71.86456, 71.88381, 71.9026, 71.92093, 71.93878, 71.95615, 71.97306, 
    71.98949, 72.00544, 72.02091, 72.0359, 72.05042, 72.06445, 72.078, 
    72.09106, 72.10364, 72.11572, 72.12733, 72.13844, 72.14907, 72.15921, 
    72.16885, 72.178, 72.18667, 72.19483, 72.20251, 72.20969, 72.21637, 
    72.22256, 72.22825, 72.23344, 72.23814, 72.24234, 72.24605, 72.24925, 
    72.25195, 72.25417, 72.25587, 72.25708, 72.25779, 72.258, 72.25771, 
    72.25692, 72.25563, 72.25385, 72.25156, 72.24878, 72.24549, 72.24171, 
    72.23743, 72.23266, 72.22739, 72.22161, 72.21535, 72.20859, 72.20132, 
    72.19357, 72.18533, 72.17659, 72.16736, 72.15764, 72.14742, 72.13672, 
    72.12553, 72.11385, 72.10168, 72.08902, 72.07588, 72.06226, 72.04816, 
    72.03356, 72.01849, 72.00294, 71.98692, 71.97042, 71.95344, 71.93599, 
    71.91806, 71.89967, 71.8808, 71.86147, 71.84166, 71.8214, 71.80066, 
    71.77947, 71.75781, 71.7357, 71.71313, 71.69011, 71.66663, 71.6427, 
    71.61832, 71.59348, 71.56821, 71.54249, 71.51633, 71.48972, 71.46268, 
    71.4352, 71.40728, 71.37893, 71.35015, 71.32095, 71.29131, 71.26125, 
    71.23076, 71.19986, 71.16853, 71.1368, 71.10464, 71.07207, 71.0391, 
    71.00571, 70.97192, 70.93773, 70.90313, 70.86813, 70.83275, 70.79696, 
    70.76078, 70.72421, 70.68726, 70.64991, 70.61218, 70.57407, 70.53559, 
    70.49673, 70.45749, 70.41788, 70.3779, 70.33755, 70.29684, 70.25576, 
    70.21432, 70.17253, 70.13039, 70.08788, 70.04502, 70.00182, 69.95827, 
    69.91438, 69.87013, 69.82555, 69.78064, 69.73539, 69.6898, 69.64389, 
    69.59765, 69.55108, 69.50419, 69.45697, 69.40944, 69.36159, 69.31342, 
    69.26494, 69.21616, 69.16705, 69.11765, 69.06795, 69.01794, 68.96763, 
    68.91702, 68.86612, 68.81493, 68.76344, 68.71167, 68.65961, 68.60727, 
    68.55464, 68.50174, 68.44855, 68.3951, 68.34137, 68.28736, 68.23309, 
    68.17855, 68.12374, 68.06867, 68.01334, 67.95776, 67.90191, 67.8458, 
    67.78945, 67.73284, 67.67599, 67.61888, 67.56154, 67.50394, 67.44611, 
    67.38804, 67.32973, 67.27118, 67.21239, 67.15339, 67.09414, 67.03467, 
    66.97498, 66.91505, 66.8549, 66.79454, 66.73395, 66.67315, 66.61213, 
    66.5509, 66.48945, 66.42779, 66.36592, 66.30385, 66.24157, 66.17909, 
    66.11641, 66.05352,
  59.60601, 59.68193, 59.75775, 59.83348, 59.90911, 59.98465, 60.0601, 
    60.13545, 60.2107, 60.28586, 60.36092, 60.43587, 60.51073, 60.58549, 
    60.66015, 60.7347, 60.80915, 60.8835, 60.95774, 61.03188, 61.10591, 
    61.17983, 61.25364, 61.32734, 61.40094, 61.47442, 61.54779, 61.62104, 
    61.69418, 61.76721, 61.84012, 61.91291, 61.98559, 62.05814, 62.13058, 
    62.20289, 62.27508, 62.34715, 62.4191, 62.49092, 62.56261, 62.63417, 
    62.70561, 62.77692, 62.84809, 62.91914, 62.99005, 63.06083, 63.13147, 
    63.20198, 63.27234, 63.34258, 63.41267, 63.48261, 63.55242, 63.62209, 
    63.6916, 63.76097, 63.8302, 63.89928, 63.96821, 64.03699, 64.10561, 
    64.17408, 64.2424, 64.31056, 64.37856, 64.44641, 64.5141, 64.58162, 
    64.64898, 64.71618, 64.78321, 64.85007, 64.91678, 64.9833, 65.04966, 
    65.11584, 65.18185, 65.24769, 65.31335, 65.37882, 65.44412, 65.50925, 
    65.57418, 65.63893, 65.7035, 65.76788, 65.83206, 65.89606, 65.95987, 
    66.02348, 66.0869, 66.15012, 66.21313, 66.27596, 66.33858, 66.40099, 
    66.4632, 66.52521, 66.587, 66.64858, 66.70995, 66.77111, 66.83205, 
    66.89278, 66.95329, 67.01357, 67.07363, 67.13347, 67.19308, 67.25246, 
    67.31161, 67.37054, 67.42922, 67.48767, 67.54588, 67.60386, 67.66159, 
    67.71908, 67.77632, 67.83331, 67.89006, 67.94656, 68.0028, 68.05878, 
    68.11451, 68.16998, 68.22519, 68.28014, 68.33482, 68.38922, 68.44337, 
    68.49724, 68.55083, 68.60416, 68.6572, 68.70996, 68.76244, 68.81464, 
    68.86654, 68.91816, 68.96949, 69.02052, 69.07127, 69.12171, 69.17185, 
    69.22169, 69.27123, 69.32046, 69.36938, 69.41799, 69.46629, 69.51427, 
    69.56194, 69.60928, 69.6563, 69.703, 69.74937, 69.79541, 69.84112, 
    69.88649, 69.93153, 69.97623, 70.02059, 70.06461, 70.10828, 70.1516, 
    70.19458, 70.23721, 70.27947, 70.32138, 70.36293, 70.40412, 70.44495, 
    70.4854, 70.52549, 70.56521, 70.60456, 70.64353, 70.68212, 70.72033, 
    70.75816, 70.79561, 70.83266, 70.86933, 70.90561, 70.94149, 70.97698, 
    71.01207, 71.04675, 71.08104, 71.11492, 71.14839, 71.18145, 71.2141, 
    71.24634, 71.27816, 71.30956, 71.34055, 71.3711, 71.40124, 71.43095, 
    71.46022, 71.48907, 71.51749, 71.54546, 71.57301, 71.60011, 71.62677, 
    71.65299, 71.67876, 71.70409, 71.72897, 71.7534, 71.77738, 71.8009, 
    71.82397, 71.84658, 71.86873, 71.89042, 71.91164, 71.9324, 71.9527, 
    71.97253, 71.99188, 72.01077, 72.02919, 72.04713, 72.0646, 72.08158, 
    72.0981, 72.11413, 72.12968, 72.14475, 72.15933, 72.17344, 72.18706, 
    72.20019, 72.21283, 72.22498, 72.23665, 72.24782, 72.2585, 72.26869, 
    72.27838, 72.28758, 72.2963, 72.3045, 72.31222, 72.31944, 72.32615, 
    72.33237, 72.3381, 72.34332, 72.34804, 72.35226, 72.35598, 72.35921, 
    72.36192, 72.36414, 72.36586, 72.36707, 72.36779, 72.368, 72.36771, 
    72.36691, 72.36562, 72.36382, 72.36153, 72.35873, 72.35543, 72.35162, 
    72.34733, 72.34252, 72.33722, 72.33142, 72.32512, 72.31832, 72.31103, 
    72.30324, 72.29494, 72.28616, 72.27689, 72.26711, 72.25684, 72.24609, 
    72.23483, 72.22309, 72.21086, 72.19814, 72.18494, 72.17124, 72.15706, 
    72.1424, 72.12725, 72.11163, 72.09551, 72.07893, 72.06187, 72.04432, 
    72.02631, 72.00781, 71.98885, 71.96942, 71.94952, 71.92915, 71.90832, 
    71.88702, 71.86526, 71.84303, 71.82035, 71.79721, 71.77362, 71.74957, 
    71.72507, 71.70012, 71.67472, 71.64887, 71.62258, 71.59586, 71.56868, 
    71.54107, 71.51302, 71.48454, 71.45562, 71.42627, 71.3965, 71.36629, 
    71.33567, 71.30462, 71.27316, 71.24126, 71.20896, 71.17625, 71.14312, 
    71.10959, 71.07565, 71.0413, 71.00655, 70.97139, 70.93584, 70.89989, 
    70.86356, 70.82683, 70.78971, 70.7522, 70.71432, 70.67604, 70.63739, 
    70.59836, 70.55895, 70.51917, 70.47903, 70.43851, 70.39763, 70.35638, 
    70.31477, 70.2728, 70.23048, 70.18781, 70.14478, 70.10139, 70.05767, 
    70.0136, 69.96918, 69.92443, 69.87934, 69.83391, 69.78815, 69.74206, 
    69.69563, 69.64888, 69.60181, 69.55441, 69.5067, 69.45867, 69.41032, 
    69.36166, 69.31269, 69.26341, 69.21383, 69.16394, 69.11375, 69.06326, 
    69.01247, 68.96139, 68.91002, 68.85835, 68.8064, 68.75416, 68.70163, 
    68.64883, 68.59574, 68.54237, 68.48873, 68.43482, 68.38064, 68.32618, 
    68.27146, 68.21648, 68.16122, 68.10571, 68.04994, 67.99392, 67.93764, 
    67.8811, 67.82432, 67.76728, 67.71, 67.65247, 67.5947, 67.53669, 
    67.47844, 67.41995, 67.36123, 67.30227, 67.24309, 67.18366, 67.12402, 
    67.06415, 67.00405, 66.94373, 66.88319, 66.82243, 66.76145, 66.70026, 
    66.63885, 66.57724, 66.51541, 66.45338, 66.39114, 66.32869, 66.26604, 
    66.20319, 66.14013,
  59.67957, 59.75558, 59.83152, 59.90736, 59.9831, 60.05875, 60.13431, 
    60.20977, 60.28514, 60.36041, 60.43558, 60.51066, 60.58563, 60.66051, 
    60.73528, 60.80995, 60.88452, 60.95899, 61.03335, 61.1076, 61.18176, 
    61.2558, 61.32973, 61.40356, 61.47728, 61.55088, 61.62437, 61.69776, 
    61.77102, 61.84418, 61.91721, 61.99014, 62.06294, 62.13562, 62.20819, 
    62.28064, 62.35296, 62.42516, 62.49724, 62.56919, 62.64101, 62.71272, 
    62.78429, 62.85573, 62.92704, 62.99823, 63.06928, 63.14019, 63.21098, 
    63.28162, 63.35213, 63.4225, 63.49274, 63.56283, 63.63278, 63.70259, 
    63.77225, 63.84177, 63.91114, 63.98037, 64.04944, 64.11837, 64.18714, 
    64.25576, 64.32423, 64.39254, 64.4607, 64.52869, 64.59653, 64.66421, 
    64.73173, 64.79908, 64.86626, 64.93329, 65.00014, 65.06683, 65.13334, 
    65.19968, 65.26585, 65.33185, 65.39767, 65.4633, 65.52876, 65.59405, 
    65.65914, 65.72406, 65.78879, 65.85333, 65.91769, 65.98185, 66.04582, 
    66.1096, 66.17318, 66.23657, 66.29976, 66.36275, 66.42554, 66.48812, 
    66.55051, 66.61268, 66.67464, 66.7364, 66.79794, 66.85928, 66.92039, 
    66.98129, 67.04197, 67.10242, 67.16266, 67.22267, 67.28246, 67.34202, 
    67.40134, 67.46044, 67.51931, 67.57793, 67.63633, 67.69448, 67.75239, 
    67.81006, 67.86748, 67.92465, 67.98158, 68.03825, 68.09468, 68.15085, 
    68.20676, 68.26241, 68.31779, 68.37292, 68.42778, 68.48238, 68.5367, 
    68.59075, 68.64453, 68.69804, 68.75126, 68.80421, 68.85686, 68.90925, 
    68.96134, 69.01314, 69.06465, 69.11587, 69.16679, 69.21742, 69.26775, 
    69.31777, 69.36749, 69.4169, 69.466, 69.51479, 69.56328, 69.61144, 
    69.65929, 69.70681, 69.75401, 69.80089, 69.84744, 69.89366, 69.93955, 
    69.98511, 70.03032, 70.0752, 70.11974, 70.16393, 70.20778, 70.25128, 
    70.29443, 70.33723, 70.37967, 70.42175, 70.46348, 70.50484, 70.54584, 
    70.58646, 70.62672, 70.66662, 70.70613, 70.74527, 70.78403, 70.8224, 
    70.8604, 70.89801, 70.93523, 70.97206, 71.0085, 71.04454, 71.08018, 
    71.11543, 71.15028, 71.18472, 71.21875, 71.25237, 71.28559, 71.31839, 
    71.35078, 71.38274, 71.41429, 71.44542, 71.47612, 71.50639, 71.53624, 
    71.56566, 71.59464, 71.6232, 71.65131, 71.67899, 71.70622, 71.73301, 
    71.75936, 71.78526, 71.81071, 71.83571, 71.86026, 71.88435, 71.908, 
    71.93118, 71.9539, 71.97616, 71.99796, 72.01929, 72.04015, 72.06055, 
    72.08047, 72.09993, 72.11892, 72.13743, 72.15546, 72.17301, 72.19009, 
    72.20669, 72.2228, 72.23843, 72.25358, 72.26824, 72.28242, 72.2961, 
    72.3093, 72.32201, 72.33423, 72.34595, 72.35719, 72.36792, 72.37817, 
    72.38791, 72.39716, 72.40591, 72.41417, 72.42192, 72.42918, 72.43593, 
    72.44218, 72.44794, 72.45319, 72.45793, 72.46218, 72.46592, 72.46915, 
    72.47189, 72.47412, 72.47585, 72.47707, 72.47778, 72.478, 72.47771, 
    72.47691, 72.47561, 72.4738, 72.47149, 72.46868, 72.46536, 72.46154, 
    72.45721, 72.45238, 72.44706, 72.44123, 72.4349, 72.42806, 72.42073, 
    72.4129, 72.40456, 72.39573, 72.3864, 72.37658, 72.36626, 72.35544, 
    72.34413, 72.33233, 72.32003, 72.30725, 72.29397, 72.2802, 72.26595, 
    72.25121, 72.23599, 72.22028, 72.20409, 72.18742, 72.17027, 72.15263, 
    72.13453, 72.11594, 72.09689, 72.07735, 72.05735, 72.03688, 72.01595, 
    71.99454, 71.97266, 71.95033, 71.92754, 71.90429, 71.88058, 71.85641, 
    71.83179, 71.80672, 71.78119, 71.75522, 71.72881, 71.70194, 71.67464, 
    71.64689, 71.61871, 71.59009, 71.56104, 71.53155, 71.50163, 71.47129, 
    71.44052, 71.40932, 71.37772, 71.34568, 71.31322, 71.28036, 71.24709, 
    71.21339, 71.1793, 71.14479, 71.10989, 71.07458, 71.03886, 71.00276, 
    70.96626, 70.92937, 70.89208, 70.85442, 70.81636, 70.77792, 70.73911, 
    70.69991, 70.66033, 70.62038, 70.58006, 70.53938, 70.49832, 70.4569, 
    70.41512, 70.37298, 70.33048, 70.28763, 70.24442, 70.20087, 70.15697, 
    70.11272, 70.06812, 70.02319, 69.97792, 69.93231, 69.88637, 69.8401, 
    69.7935, 69.74657, 69.69931, 69.65174, 69.60384, 69.55563, 69.5071, 
    69.45826, 69.4091, 69.35964, 69.30988, 69.2598, 69.20943, 69.15876, 
    69.10779, 69.05653, 69.00497, 68.95312, 68.90098, 68.84856, 68.79585, 
    68.74286, 68.68959, 68.63605, 68.58222, 68.52813, 68.47376, 68.41912, 
    68.36422, 68.30905, 68.25362, 68.19793, 68.14198, 68.08577, 68.0293, 
    67.9726, 67.91563, 67.85841, 67.80095, 67.74325, 67.6853, 67.62711, 
    67.56868, 67.51001, 67.45111, 67.39198, 67.33261, 67.27302, 67.2132, 
    67.15314, 67.09288, 67.03238, 66.97166, 66.91074, 66.84959, 66.78822, 
    66.72665, 66.66486, 66.60286, 66.54065, 66.47823, 66.41562, 66.3528, 
    66.28978, 66.22655,
  59.75291, 59.82904, 59.90509, 59.98103, 60.05689, 60.13265, 60.20832, 
    60.2839, 60.35938, 60.43476, 60.51005, 60.58524, 60.66033, 60.73532, 
    60.81021, 60.885, 60.95969, 61.03427, 61.10875, 61.18313, 61.2574, 
    61.33157, 61.40562, 61.47957, 61.55341, 61.62714, 61.70076, 61.77427, 
    61.84766, 61.92094, 61.99411, 62.06716, 62.14009, 62.21291, 62.2856, 
    62.35818, 62.43063, 62.50296, 62.57518, 62.64726, 62.71922, 62.79106, 
    62.86277, 62.93435, 63.00579, 63.07711, 63.1483, 63.21936, 63.29028, 
    63.36107, 63.43172, 63.50223, 63.57261, 63.64284, 63.71294, 63.78289, 
    63.8527, 63.92236, 63.99188, 64.06125, 64.13048, 64.19955, 64.26847, 
    64.33724, 64.40586, 64.47433, 64.54263, 64.61078, 64.67877, 64.7466, 
    64.81428, 64.88178, 64.94913, 65.0163, 65.08331, 65.15015, 65.21683, 
    65.28333, 65.34966, 65.41581, 65.48179, 65.54759, 65.61321, 65.67866, 
    65.74392, 65.809, 65.87389, 65.9386, 66.00312, 66.06745, 66.13158, 
    66.19553, 66.25928, 66.32284, 66.3862, 66.44936, 66.51231, 66.57507, 
    66.63762, 66.69997, 66.76211, 66.82404, 66.88575, 66.94726, 67.00854, 
    67.06962, 67.13047, 67.19111, 67.25152, 67.31171, 67.37167, 67.4314, 
    67.49091, 67.55019, 67.60923, 67.66804, 67.72661, 67.78493, 67.84303, 
    67.90087, 67.95847, 68.01583, 68.07294, 68.1298, 68.1864, 68.24275, 
    68.29884, 68.35468, 68.41025, 68.46555, 68.5206, 68.57538, 68.62988, 
    68.68412, 68.73808, 68.79177, 68.84518, 68.89831, 68.95116, 69.00372, 
    69.05599, 69.10798, 69.15968, 69.21107, 69.26218, 69.313, 69.3635, 
    69.41371, 69.46362, 69.51321, 69.5625, 69.61147, 69.66013, 69.70848, 
    69.75651, 69.80421, 69.8516, 69.89866, 69.9454, 69.9918, 70.03786, 
    70.0836, 70.129, 70.17406, 70.21877, 70.26315, 70.30717, 70.35085, 
    70.39418, 70.43716, 70.47977, 70.52203, 70.56393, 70.60546, 70.64664, 
    70.68744, 70.72787, 70.76793, 70.80761, 70.84692, 70.88585, 70.92439, 
    70.96255, 71.00033, 71.03771, 71.07471, 71.11131, 71.14751, 71.18332, 
    71.21873, 71.25372, 71.28832, 71.32251, 71.35629, 71.38966, 71.42261, 
    71.45515, 71.48727, 71.51896, 71.55023, 71.58108, 71.6115, 71.64149, 
    71.67104, 71.70017, 71.72886, 71.75711, 71.78492, 71.81229, 71.8392, 
    71.86568, 71.89171, 71.91729, 71.94241, 71.96708, 71.99129, 72.01505, 
    72.03835, 72.06119, 72.08356, 72.10546, 72.1269, 72.14787, 72.16837, 
    72.1884, 72.20795, 72.22704, 72.24564, 72.26376, 72.28141, 72.29858, 
    72.31526, 72.33146, 72.34717, 72.3624, 72.37714, 72.39138, 72.40514, 
    72.41841, 72.43118, 72.44347, 72.45525, 72.46655, 72.47734, 72.48763, 
    72.49743, 72.50673, 72.51553, 72.52383, 72.53162, 72.53892, 72.54571, 
    72.55199, 72.55778, 72.56305, 72.56783, 72.57209, 72.57585, 72.57911, 
    72.58186, 72.5841, 72.58584, 72.58707, 72.58778, 72.588, 72.58771, 
    72.58691, 72.58559, 72.58378, 72.58146, 72.57863, 72.57529, 72.57145, 
    72.56711, 72.56225, 72.55689, 72.55103, 72.54466, 72.5378, 72.53042, 
    72.52254, 72.51417, 72.50529, 72.49592, 72.48604, 72.47566, 72.46479, 
    72.45342, 72.44156, 72.4292, 72.41634, 72.403, 72.38916, 72.37483, 
    72.36002, 72.34472, 72.32893, 72.31265, 72.29589, 72.27866, 72.26093, 
    72.24273, 72.22405, 72.2049, 72.18526, 72.16516, 72.14458, 72.12354, 
    72.10203, 72.08005, 72.0576, 72.0347, 72.01132, 71.9875, 71.96321, 
    71.93847, 71.91327, 71.88762, 71.86153, 71.83498, 71.80798, 71.78055, 
    71.75267, 71.72435, 71.69559, 71.6664, 71.63677, 71.60671, 71.57623, 
    71.54531, 71.51398, 71.48221, 71.45003, 71.41743, 71.38441, 71.35098, 
    71.31713, 71.28288, 71.24821, 71.21315, 71.17768, 71.14182, 71.10555, 
    71.06889, 71.03183, 70.99438, 70.95654, 70.91832, 70.87971, 70.84073, 
    70.80136, 70.76161, 70.7215, 70.68101, 70.64014, 70.59892, 70.55733, 
    70.51537, 70.47305, 70.43038, 70.38735, 70.34396, 70.30023, 70.25615, 
    70.21172, 70.16695, 70.12184, 70.07639, 70.0306, 69.98447, 69.93803, 
    69.89124, 69.84413, 69.79669, 69.74893, 69.70086, 69.65246, 69.60374, 
    69.55473, 69.50539, 69.45574, 69.40579, 69.35554, 69.30498, 69.25412, 
    69.20296, 69.15152, 69.09978, 69.04774, 68.99542, 68.94281, 68.88992, 
    68.83675, 68.78329, 68.72957, 68.67556, 68.62128, 68.56673, 68.51191, 
    68.45683, 68.40147, 68.34586, 68.28999, 68.23386, 68.17746, 68.12082, 
    68.06393, 68.00677, 67.94938, 67.89174, 67.83385, 67.77573, 67.71735, 
    67.65875, 67.59991, 67.54082, 67.48151, 67.42197, 67.3622, 67.3022, 
    67.24197, 67.18153, 67.12086, 67.05997, 66.99886, 66.93754, 66.876, 
    66.81425, 66.75229, 66.69012, 66.62774, 66.56516, 66.50237, 66.43938, 
    66.37619, 66.3128,
  59.82606, 59.9023, 59.97845, 60.05451, 60.13048, 60.20635, 60.28213, 
    60.35782, 60.43341, 60.50891, 60.58431, 60.65961, 60.73482, 60.80993, 
    60.88494, 60.95985, 61.03465, 61.10936, 61.18396, 61.25845, 61.33284, 
    61.40713, 61.48131, 61.55538, 61.62934, 61.7032, 61.77694, 61.85058, 
    61.9241, 61.99751, 62.0708, 62.14397, 62.21704, 62.28998, 62.36281, 
    62.43551, 62.5081, 62.58057, 62.65291, 62.72513, 62.79723, 62.8692, 
    62.94104, 63.01276, 63.08434, 63.1558, 63.22713, 63.29832, 63.36938, 
    63.44031, 63.5111, 63.58176, 63.65228, 63.72266, 63.79289, 63.86299, 
    63.93295, 64.00275, 64.07242, 64.14194, 64.21131, 64.28053, 64.34961, 
    64.41853, 64.4873, 64.55591, 64.62437, 64.69267, 64.76082, 64.8288, 
    64.89663, 64.96429, 65.03179, 65.09912, 65.16629, 65.23329, 65.30013, 
    65.36678, 65.43327, 65.49959, 65.56573, 65.63169, 65.69747, 65.76308, 
    65.82851, 65.89375, 65.95881, 66.02368, 66.08836, 66.15286, 66.21716, 
    66.28128, 66.3452, 66.40892, 66.47245, 66.53578, 66.59891, 66.66183, 
    66.72456, 66.78708, 66.84939, 66.91149, 66.97338, 67.03506, 67.09652, 
    67.15777, 67.2188, 67.27961, 67.34019, 67.40057, 67.4607, 67.52061, 
    67.5803, 67.63976, 67.69897, 67.75797, 67.81671, 67.87523, 67.93349, 
    67.99152, 68.04931, 68.10685, 68.16414, 68.22118, 68.27796, 68.3345, 
    68.39077, 68.44678, 68.50254, 68.55803, 68.61326, 68.66822, 68.72292, 
    68.77734, 68.83148, 68.88535, 68.93895, 68.99226, 69.0453, 69.09804, 
    69.15051, 69.20267, 69.25455, 69.30614, 69.35744, 69.40843, 69.45913, 
    69.50952, 69.55961, 69.60939, 69.65886, 69.70802, 69.75687, 69.8054, 
    69.85361, 69.9015, 69.94907, 69.99632, 70.04323, 70.08981, 70.13606, 
    70.18198, 70.22756, 70.2728, 70.3177, 70.36225, 70.40646, 70.45032, 
    70.49382, 70.53697, 70.57977, 70.6222, 70.66428, 70.70599, 70.74734, 
    70.78831, 70.82892, 70.86915, 70.909, 70.94848, 70.98758, 71.02629, 
    71.06462, 71.10256, 71.14011, 71.17728, 71.21404, 71.25041, 71.28638, 
    71.32195, 71.3571, 71.39186, 71.42621, 71.46014, 71.49366, 71.52677, 
    71.55946, 71.59172, 71.62357, 71.65499, 71.68598, 71.71655, 71.74668, 
    71.77638, 71.80565, 71.83447, 71.86285, 71.8908, 71.9183, 71.94536, 
    71.97196, 71.99812, 72.02382, 72.04907, 72.07387, 72.0982, 72.12208, 
    72.14549, 72.16844, 72.19093, 72.21294, 72.23449, 72.25557, 72.27617, 
    72.2963, 72.31596, 72.33514, 72.35384, 72.37206, 72.38979, 72.40704, 
    72.42381, 72.44009, 72.45589, 72.4712, 72.48602, 72.50034, 72.51417, 
    72.5275, 72.54035, 72.5527, 72.56454, 72.5759, 72.58675, 72.5971, 
    72.60695, 72.61629, 72.62514, 72.63348, 72.64132, 72.64865, 72.65548, 
    72.6618, 72.66761, 72.67292, 72.67772, 72.68201, 72.68579, 72.68906, 
    72.69183, 72.69408, 72.69582, 72.69706, 72.69778, 72.698, 72.6977, 
    72.6969, 72.69558, 72.69376, 72.69142, 72.68858, 72.68523, 72.68137, 
    72.67699, 72.67211, 72.66673, 72.66084, 72.65443, 72.64752, 72.64011, 
    72.63219, 72.62377, 72.61485, 72.60542, 72.59549, 72.58506, 72.57413, 
    72.56271, 72.55077, 72.53835, 72.52543, 72.51202, 72.49811, 72.4837, 
    72.46881, 72.45343, 72.43755, 72.4212, 72.40435, 72.38702, 72.36921, 
    72.35091, 72.33214, 72.31288, 72.29315, 72.27294, 72.25227, 72.23111, 
    72.20949, 72.1874, 72.16484, 72.14182, 72.11833, 72.09438, 72.06997, 
    72.0451, 72.01978, 71.99401, 71.96778, 71.94111, 71.91398, 71.88641, 
    71.8584, 71.82994, 71.80105, 71.77171, 71.74194, 71.71174, 71.68111, 
    71.65005, 71.61856, 71.58665, 71.55431, 71.52156, 71.48839, 71.4548, 
    71.4208, 71.38639, 71.35157, 71.31635, 71.28072, 71.24468, 71.20825, 
    71.17142, 71.1342, 71.09659, 71.05859, 71.0202, 70.98142, 70.94226, 
    70.90273, 70.86281, 70.82252, 70.78185, 70.74082, 70.69942, 70.65765, 
    70.61552, 70.57302, 70.53017, 70.48696, 70.44341, 70.39949, 70.35522, 
    70.31062, 70.26567, 70.22038, 70.17474, 70.12877, 70.08247, 70.03583, 
    69.98886, 69.94157, 69.89394, 69.84601, 69.79774, 69.74916, 69.70026, 
    69.65105, 69.60153, 69.5517, 69.50157, 69.45113, 69.40038, 69.34934, 
    69.298, 69.24637, 69.19444, 69.14222, 69.08971, 69.03693, 68.98385, 
    68.93049, 68.87685, 68.82294, 68.76875, 68.71428, 68.65955, 68.60455, 
    68.54927, 68.49374, 68.43794, 68.38188, 68.32557, 68.269, 68.21217, 
    68.15509, 68.09776, 68.04018, 67.98236, 67.92429, 67.86598, 67.80743, 
    67.74865, 67.68963, 67.63037, 67.57088, 67.51115, 67.45121, 67.39103, 
    67.33063, 67.27, 67.20916, 67.14809, 67.08681, 67.02531, 66.9636, 
    66.90168, 66.83955, 66.7772, 66.71465, 66.65189, 66.58894, 66.52578, 
    66.46242, 66.39886,
  59.89901, 59.97536, 60.05161, 60.12778, 60.20386, 60.27985, 60.35574, 
    60.43154, 60.50724, 60.58286, 60.65837, 60.73379, 60.80911, 60.88433, 
    60.95946, 61.03448, 61.10941, 61.18423, 61.25895, 61.33357, 61.40808, 
    61.48249, 61.55679, 61.63099, 61.70507, 61.77905, 61.85292, 61.92668, 
    62.00033, 62.07386, 62.14728, 62.22059, 62.29378, 62.36685, 62.43981, 
    62.51265, 62.58537, 62.65796, 62.73044, 62.8028, 62.87502, 62.94713, 
    63.01911, 63.09096, 63.16269, 63.23428, 63.30575, 63.37708, 63.44828, 
    63.51935, 63.59029, 63.66108, 63.73174, 63.80227, 63.87265, 63.94289, 
    64.01299, 64.08295, 64.15276, 64.22243, 64.29195, 64.36131, 64.43054, 
    64.49961, 64.56853, 64.6373, 64.70591, 64.77436, 64.84266, 64.9108, 
    64.97878, 65.0466, 65.11425, 65.18175, 65.24907, 65.31623, 65.38322, 
    65.45004, 65.51669, 65.58316, 65.64947, 65.71559, 65.78154, 65.84731, 
    65.9129, 65.9783, 66.04353, 66.10857, 66.17342, 66.23808, 66.30255, 
    66.36684, 66.43092, 66.49482, 66.55852, 66.62202, 66.68532, 66.74841, 
    66.81131, 66.874, 66.93649, 66.99876, 67.06082, 67.12268, 67.18432, 
    67.24574, 67.30695, 67.36794, 67.4287, 67.48924, 67.54956, 67.60966, 
    67.66952, 67.72916, 67.78855, 67.84772, 67.90665, 67.96535, 68.0238, 
    68.08201, 68.13998, 68.19769, 68.25517, 68.31239, 68.36935, 68.42607, 
    68.48253, 68.53873, 68.59467, 68.65035, 68.70576, 68.76091, 68.81579, 
    68.87039, 68.92473, 68.97878, 69.03257, 69.08607, 69.13928, 69.19222, 
    69.24487, 69.29723, 69.3493, 69.40107, 69.45255, 69.50373, 69.55461, 
    69.60519, 69.65546, 69.70543, 69.75509, 69.80444, 69.85347, 69.90218, 
    69.95058, 69.99866, 70.04641, 70.09384, 70.14094, 70.18771, 70.23415, 
    70.28024, 70.326, 70.37143, 70.41651, 70.46124, 70.50563, 70.54967, 
    70.59335, 70.63669, 70.67966, 70.72227, 70.76453, 70.80641, 70.84794, 
    70.88908, 70.92987, 70.97028, 71.0103, 71.04996, 71.08923, 71.12811, 
    71.16661, 71.20472, 71.24244, 71.27976, 71.3167, 71.35323, 71.38936, 
    71.42509, 71.46041, 71.49532, 71.52983, 71.56392, 71.5976, 71.63086, 
    71.6637, 71.69612, 71.72812, 71.75969, 71.79083, 71.82154, 71.85182, 
    71.88166, 71.91106, 71.94003, 71.96856, 71.99664, 72.02428, 72.05146, 
    72.0782, 72.10448, 72.13032, 72.15569, 72.18061, 72.20507, 72.22906, 
    72.25259, 72.27566, 72.29826, 72.32039, 72.34205, 72.36324, 72.38394, 
    72.40418, 72.42393, 72.44321, 72.46201, 72.48032, 72.49815, 72.5155, 
    72.53236, 72.54872, 72.5646, 72.57999, 72.59488, 72.60928, 72.62318, 
    72.63659, 72.64951, 72.66191, 72.67383, 72.68523, 72.69614, 72.70655, 
    72.71645, 72.72585, 72.73475, 72.74313, 72.75101, 72.75838, 72.76525, 
    72.77161, 72.77745, 72.78278, 72.78761, 72.79192, 72.79572, 72.79901, 
    72.8018, 72.80406, 72.80581, 72.80705, 72.80779, 72.808, 72.8077, 
    72.80689, 72.80557, 72.80373, 72.80138, 72.79853, 72.79516, 72.79128, 
    72.78688, 72.78197, 72.77656, 72.77063, 72.7642, 72.75726, 72.7498, 
    72.74184, 72.73338, 72.7244, 72.71492, 72.70494, 72.69446, 72.68346, 
    72.67197, 72.65998, 72.64749, 72.63451, 72.62102, 72.60703, 72.59256, 
    72.57758, 72.56212, 72.54617, 72.52972, 72.51279, 72.49537, 72.47746, 
    72.45907, 72.4402, 72.42085, 72.40101, 72.3807, 72.35992, 72.33865, 
    72.31692, 72.29472, 72.27204, 72.2489, 72.2253, 72.20123, 72.1767, 
    72.15171, 72.12626, 72.10036, 72.074, 72.04719, 72.01994, 71.99223, 
    71.96407, 71.93548, 71.90645, 71.87697, 71.84706, 71.81671, 71.78593, 
    71.75472, 71.72308, 71.69102, 71.65853, 71.62563, 71.5923, 71.55856, 
    71.5244, 71.48983, 71.45485, 71.41946, 71.38367, 71.34747, 71.31087, 
    71.27389, 71.2365, 71.19872, 71.16055, 71.12199, 71.08304, 71.04371, 
    71.004, 70.96391, 70.92344, 70.8826, 70.84139, 70.79981, 70.75787, 
    70.71556, 70.67288, 70.62985, 70.58647, 70.54272, 70.49863, 70.45419, 
    70.4094, 70.36427, 70.31879, 70.27297, 70.22682, 70.18033, 70.13351, 
    70.08636, 70.03888, 69.99107, 69.94295, 69.8945, 69.84573, 69.79665, 
    69.74725, 69.69755, 69.64753, 69.59721, 69.54659, 69.49565, 69.44443, 
    69.3929, 69.34108, 69.28896, 69.23656, 69.18387, 69.13088, 69.07762, 
    69.02408, 68.97025, 68.91615, 68.86178, 68.80713, 68.7522, 68.69701, 
    68.64156, 68.58585, 68.52986, 68.47362, 68.41712, 68.36036, 68.30335, 
    68.24609, 68.18858, 68.13082, 68.07281, 68.01456, 67.95608, 67.89735, 
    67.83838, 67.77917, 67.71973, 67.66006, 67.60017, 67.54004, 67.47968, 
    67.41911, 67.3583, 67.29728, 67.23604, 67.17458, 67.11291, 67.05102, 
    66.98892, 66.92661, 66.8641, 66.80138, 66.73845, 66.67532, 66.61198, 
    66.54845, 66.48473,
  59.97175, 60.0482, 60.12457, 60.20085, 60.27703, 60.35313, 60.42914, 
    60.50505, 60.58087, 60.65659, 60.73222, 60.80776, 60.88319, 60.95853, 
    61.03378, 61.10892, 61.18396, 61.2589, 61.33374, 61.40848, 61.48312, 
    61.55764, 61.63207, 61.70639, 61.7806, 61.8547, 61.92869, 62.00258, 
    62.07635, 62.15001, 62.22356, 62.29699, 62.37031, 62.44352, 62.51661, 
    62.58957, 62.66242, 62.73515, 62.80777, 62.88025, 62.95262, 63.02486, 
    63.09697, 63.16896, 63.24083, 63.31256, 63.38416, 63.45564, 63.52698, 
    63.59819, 63.66926, 63.7402, 63.811, 63.88167, 63.9522, 64.02258, 
    64.09283, 64.16293, 64.23289, 64.3027, 64.37238, 64.44189, 64.51127, 
    64.58049, 64.64956, 64.71848, 64.78724, 64.85585, 64.9243, 64.9926, 
    65.06073, 65.12871, 65.19652, 65.26417, 65.33165, 65.39897, 65.46612, 
    65.5331, 65.59991, 65.66654, 65.73301, 65.79929, 65.86541, 65.93134, 
    65.99709, 66.06267, 66.12805, 66.19326, 66.25828, 66.32311, 66.38775, 
    66.4522, 66.51646, 66.58053, 66.64439, 66.70806, 66.77154, 66.83481, 
    66.89787, 66.96074, 67.0234, 67.08585, 67.14809, 67.21011, 67.27193, 
    67.33353, 67.39491, 67.45608, 67.51702, 67.57774, 67.63824, 67.69852, 
    67.75856, 67.81837, 67.87795, 67.9373, 67.99641, 68.05529, 68.11392, 
    68.17232, 68.23047, 68.28837, 68.34603, 68.40343, 68.46059, 68.51749, 
    68.57413, 68.63052, 68.68665, 68.74251, 68.79811, 68.85344, 68.90851, 
    68.9633, 69.01782, 69.07207, 69.12603, 69.17972, 69.23312, 69.28625, 
    69.33908, 69.39163, 69.44389, 69.49585, 69.54752, 69.59888, 69.64996, 
    69.70072, 69.75118, 69.80134, 69.85118, 69.90072, 69.94994, 69.99884, 
    70.04742, 70.09569, 70.14363, 70.19124, 70.23853, 70.28548, 70.3321, 
    70.37839, 70.42433, 70.46994, 70.51521, 70.56012, 70.60469, 70.64891, 
    70.69278, 70.73629, 70.77945, 70.82224, 70.86467, 70.90674, 70.94844, 
    70.98977, 71.03072, 71.0713, 71.11151, 71.15134, 71.19077, 71.22984, 
    71.2685, 71.30679, 71.34467, 71.38216, 71.41927, 71.45596, 71.49226, 
    71.52815, 71.56364, 71.59872, 71.63338, 71.66763, 71.70147, 71.73489, 
    71.76788, 71.80045, 71.8326, 71.86433, 71.89561, 71.92648, 71.9569, 
    71.98689, 72.01643, 72.04555, 72.07421, 72.10243, 72.1302, 72.15752, 
    72.18439, 72.21081, 72.23677, 72.26228, 72.28732, 72.3119, 72.33601, 
    72.35966, 72.38285, 72.40556, 72.42781, 72.44958, 72.47087, 72.49169, 
    72.51203, 72.53189, 72.55127, 72.57016, 72.58857, 72.60649, 72.62393, 
    72.64088, 72.65733, 72.67329, 72.68876, 72.70373, 72.71821, 72.73219, 
    72.74567, 72.75864, 72.77113, 72.7831, 72.79457, 72.80554, 72.816, 
    72.82596, 72.83541, 72.84435, 72.85278, 72.8607, 72.86812, 72.87502, 
    72.8814, 72.88728, 72.89265, 72.8975, 72.90183, 72.90565, 72.90897, 
    72.91176, 72.91404, 72.9158, 72.91705, 72.91778, 72.918, 72.9177, 
    72.91689, 72.91556, 72.91371, 72.91135, 72.90848, 72.90508, 72.90118, 
    72.89677, 72.89183, 72.88638, 72.88042, 72.87395, 72.86697, 72.85948, 
    72.85148, 72.84297, 72.83395, 72.82442, 72.81438, 72.80384, 72.79279, 
    72.78124, 72.76918, 72.75662, 72.74357, 72.73001, 72.71595, 72.70139, 
    72.68635, 72.6708, 72.65476, 72.63823, 72.6212, 72.60369, 72.58569, 
    72.56721, 72.54823, 72.52878, 72.50884, 72.48843, 72.46754, 72.44617, 
    72.42432, 72.402, 72.37921, 72.35596, 72.33223, 72.30804, 72.28339, 
    72.25827, 72.2327, 72.20666, 72.18018, 72.15323, 72.12584, 72.09799, 
    72.0697, 72.04097, 72.0118, 71.98217, 71.95212, 71.92162, 71.89069, 
    71.85934, 71.82755, 71.79533, 71.76269, 71.72963, 71.69614, 71.66224, 
    71.62792, 71.59319, 71.55805, 71.5225, 71.48654, 71.45019, 71.41342, 
    71.37627, 71.33871, 71.30076, 71.26241, 71.22368, 71.18456, 71.14506, 
    71.10517, 71.06491, 71.02427, 70.98325, 70.94186, 70.90011, 70.85799, 
    70.8155, 70.77264, 70.72943, 70.68587, 70.64194, 70.59766, 70.55304, 
    70.50806, 70.46275, 70.41709, 70.37109, 70.32475, 70.27808, 70.23107, 
    70.18373, 70.13606, 70.08807, 70.03976, 69.99113, 69.94217, 69.89291, 
    69.84332, 69.79343, 69.74322, 69.69271, 69.6419, 69.59078, 69.53936, 
    69.48765, 69.43564, 69.38334, 69.33074, 69.27786, 69.2247, 69.17125, 
    69.11752, 69.0635, 69.00922, 68.95465, 68.89982, 68.84471, 68.78933, 
    68.73369, 68.67779, 68.62162, 68.56519, 68.50851, 68.45157, 68.39437, 
    68.33692, 68.27923, 68.22128, 68.1631, 68.10467, 68.04599, 67.98708, 
    67.92793, 67.86855, 67.80893, 67.74908, 67.689, 67.62869, 67.56815, 
    67.5074, 67.44642, 67.38522, 67.3238, 67.26217, 67.20032, 67.13825, 
    67.07598, 67.0135, 66.95081, 66.88791, 66.82481, 66.76151, 66.69801, 
    66.6343, 66.5704,
  60.04428, 60.12085, 60.19732, 60.27371, 60.35001, 60.42622, 60.50233, 
    60.57836, 60.65429, 60.73013, 60.80587, 60.88152, 60.95707, 61.03253, 
    61.10789, 61.18315, 61.2583, 61.33337, 61.40833, 61.48318, 61.55794, 
    61.63259, 61.70713, 61.78157, 61.85591, 61.93014, 62.00426, 62.07827, 
    62.15216, 62.22595, 62.29963, 62.37319, 62.44664, 62.51997, 62.59319, 
    62.66629, 62.73927, 62.81214, 62.88488, 62.9575, 63.03, 63.10238, 
    63.17463, 63.24675, 63.31876, 63.39062, 63.46237, 63.53398, 63.60546, 
    63.67682, 63.74803, 63.81911, 63.89006, 63.96087, 64.03154, 64.10207, 
    64.17246, 64.24271, 64.31282, 64.38278, 64.4526, 64.52227, 64.59179, 
    64.66116, 64.73038, 64.79945, 64.86838, 64.93713, 65.00574, 65.0742, 
    65.14249, 65.21062, 65.27858, 65.34639, 65.41403, 65.48151, 65.54881, 
    65.61596, 65.68293, 65.74973, 65.81635, 65.8828, 65.94908, 66.01517, 
    66.08109, 66.14683, 66.21239, 66.27776, 66.34294, 66.40794, 66.47276, 
    66.53738, 66.60181, 66.66604, 66.73008, 66.79392, 66.85757, 66.92101, 
    66.98425, 67.04729, 67.11012, 67.17274, 67.23516, 67.29736, 67.35936, 
    67.42113, 67.4827, 67.54404, 67.60516, 67.66607, 67.72675, 67.78719, 
    67.84742, 67.90742, 67.96718, 68.02671, 68.08601, 68.14507, 68.20388, 
    68.26246, 68.32079, 68.37888, 68.43672, 68.49432, 68.55165, 68.60874, 
    68.66557, 68.72215, 68.77846, 68.8345, 68.8903, 68.94582, 69.00107, 
    69.05605, 69.11076, 69.16519, 69.21935, 69.27322, 69.32681, 69.38013, 
    69.43315, 69.48589, 69.53833, 69.59048, 69.64234, 69.69389, 69.74516, 
    69.79611, 69.84676, 69.8971, 69.94714, 69.99686, 70.04627, 70.09536, 
    70.14413, 70.19259, 70.24072, 70.28851, 70.33599, 70.38313, 70.42994, 
    70.47641, 70.52254, 70.56834, 70.61378, 70.65888, 70.70364, 70.74804, 
    70.79209, 70.83578, 70.87913, 70.9221, 70.96471, 71.00696, 71.04884, 
    71.09035, 71.13148, 71.17224, 71.21262, 71.25262, 71.29224, 71.33147, 
    71.37031, 71.40876, 71.44682, 71.48449, 71.52175, 71.55862, 71.59509, 
    71.63114, 71.66679, 71.70203, 71.73686, 71.77127, 71.80527, 71.83884, 
    71.87199, 71.90472, 71.93703, 71.9689, 72.00034, 72.03135, 72.06192, 
    72.09206, 72.12175, 72.151, 72.17981, 72.20817, 72.23608, 72.26353, 
    72.29054, 72.31709, 72.34319, 72.36881, 72.39398, 72.41869, 72.44293, 
    72.46671, 72.49001, 72.51284, 72.53519, 72.55708, 72.57848, 72.59941, 
    72.61986, 72.63982, 72.65929, 72.67829, 72.6968, 72.71481, 72.73235, 
    72.74937, 72.76592, 72.78197, 72.79752, 72.81257, 72.82713, 72.84118, 
    72.85473, 72.86777, 72.88033, 72.89236, 72.9039, 72.91492, 72.92545, 
    72.93546, 72.94495, 72.95395, 72.96243, 72.97039, 72.97784, 72.98478, 
    72.9912, 72.99712, 73.0025, 73.00739, 73.01174, 73.01559, 73.01891, 
    73.02172, 73.02402, 73.02579, 73.02705, 73.02778, 73.028, 73.02769, 
    73.02688, 73.02554, 73.02369, 73.02132, 73.01842, 73.01501, 73.01109, 
    73.00665, 73.00169, 72.99622, 72.99022, 72.98372, 72.9767, 72.96916, 
    72.96111, 72.95256, 72.94349, 72.93391, 72.92381, 72.91322, 72.90211, 
    72.8905, 72.87837, 72.86575, 72.85262, 72.83899, 72.82485, 72.81022, 
    72.79509, 72.77946, 72.76334, 72.74671, 72.7296, 72.712, 72.6939, 
    72.67532, 72.65625, 72.6367, 72.61665, 72.59613, 72.57513, 72.55365, 
    72.53169, 72.50925, 72.48635, 72.46297, 72.43913, 72.41481, 72.39003, 
    72.36479, 72.33909, 72.31292, 72.2863, 72.25922, 72.23169, 72.20371, 
    72.17529, 72.14641, 72.11708, 72.08732, 72.05711, 72.02647, 71.9954, 
    71.96389, 71.93195, 71.89957, 71.86678, 71.83356, 71.79992, 71.76585, 
    71.73138, 71.69649, 71.66118, 71.62547, 71.58934, 71.55282, 71.51588, 
    71.47855, 71.44083, 71.40271, 71.36419, 71.32529, 71.286, 71.24632, 
    71.20626, 71.16582, 71.125, 71.0838, 71.04224, 71.0003, 70.95799, 
    70.91533, 70.87229, 70.8289, 70.78515, 70.74104, 70.69659, 70.65177, 
    70.60661, 70.56111, 70.51527, 70.46908, 70.42255, 70.37569, 70.3285, 
    70.28098, 70.23312, 70.18494, 70.13644, 70.08762, 70.03848, 69.98902, 
    69.93925, 69.88916, 69.83877, 69.78807, 69.73707, 69.68576, 69.63416, 
    69.58225, 69.53005, 69.47756, 69.42478, 69.37171, 69.31836, 69.26472, 
    69.2108, 69.15659, 69.10212, 69.04737, 68.99234, 68.93705, 68.88148, 
    68.82566, 68.76956, 68.71321, 68.65659, 68.59972, 68.5426, 68.48522, 
    68.42759, 68.36971, 68.31158, 68.2532, 68.1946, 68.13573, 68.07664, 
    68.01731, 67.95774, 67.89794, 67.83791, 67.77765, 67.71716, 67.65645, 
    67.59551, 67.53436, 67.47298, 67.41138, 67.34956, 67.28754, 67.2253, 
    67.16285, 67.1002, 67.03733, 66.97426, 66.91099, 66.84751, 66.78384, 
    66.71996, 66.65589,
  60.11661, 60.19328, 60.26987, 60.34636, 60.42277, 60.49909, 60.57532, 
    60.65145, 60.7275, 60.80345, 60.87931, 60.95507, 61.03074, 61.10631, 
    61.18179, 61.25716, 61.33244, 61.40762, 61.4827, 61.55767, 61.63255, 
    61.70732, 61.78199, 61.85656, 61.93101, 62.00536, 62.07961, 62.15374, 
    62.22777, 62.30168, 62.37548, 62.44918, 62.52275, 62.59622, 62.66957, 
    62.7428, 62.81591, 62.88891, 62.96178, 63.03454, 63.10717, 63.17969, 
    63.25208, 63.32434, 63.39647, 63.46848, 63.54037, 63.61212, 63.68374, 
    63.75523, 63.82659, 63.89782, 63.96891, 64.03986, 64.11067, 64.18135, 
    64.25189, 64.32229, 64.39254, 64.46265, 64.53262, 64.60243, 64.67211, 
    64.74163, 64.811, 64.88023, 64.9493, 65.01822, 65.08698, 65.15558, 
    65.22403, 65.29231, 65.36044, 65.42841, 65.49621, 65.56384, 65.63131, 
    65.69862, 65.76575, 65.8327, 65.89949, 65.96611, 66.03255, 66.09881, 
    66.16489, 66.2308, 66.29652, 66.36206, 66.42741, 66.49258, 66.55756, 
    66.62235, 66.68695, 66.75136, 66.81557, 66.87959, 66.9434, 67.00702, 
    67.07043, 67.13364, 67.19666, 67.25945, 67.32204, 67.38443, 67.4466, 
    67.50855, 67.5703, 67.63182, 67.69312, 67.7542, 67.81506, 67.87569, 
    67.9361, 67.99628, 68.05622, 68.11594, 68.17542, 68.23466, 68.29366, 
    68.35242, 68.41094, 68.46922, 68.52724, 68.58502, 68.64255, 68.69982, 
    68.75684, 68.8136, 68.8701, 68.92634, 68.98232, 69.03802, 69.09346, 
    69.14864, 69.20353, 69.25816, 69.3125, 69.36656, 69.42035, 69.47385, 
    69.52706, 69.57999, 69.63263, 69.68497, 69.73701, 69.78876, 69.84021, 
    69.89136, 69.9422, 69.99274, 70.04296, 70.09287, 70.14247, 70.19175, 
    70.24072, 70.28935, 70.33767, 70.38566, 70.43332, 70.48065, 70.52765, 
    70.5743, 70.62063, 70.6666, 70.71224, 70.75753, 70.80247, 70.84706, 
    70.8913, 70.93517, 70.97869, 71.02185, 71.06464, 71.10708, 71.14913, 
    71.19082, 71.23214, 71.27307, 71.31363, 71.35381, 71.3936, 71.43301, 
    71.47203, 71.51065, 71.54889, 71.58672, 71.62416, 71.66119, 71.69782, 
    71.73405, 71.76987, 71.80527, 71.84026, 71.87484, 71.909, 71.94273, 
    71.97604, 72.00893, 72.04139, 72.07342, 72.10501, 72.13617, 72.16689, 
    72.19717, 72.22701, 72.25641, 72.28535, 72.31386, 72.3419, 72.3695, 
    72.39664, 72.42332, 72.44955, 72.47531, 72.50061, 72.52544, 72.5498, 
    72.5737, 72.59713, 72.62008, 72.64255, 72.66454, 72.68607, 72.7071, 
    72.72765, 72.74772, 72.7673, 72.7864, 72.805, 72.82311, 72.84074, 
    72.85786, 72.87449, 72.89062, 72.90626, 72.92139, 72.93603, 72.95016, 
    72.96378, 72.9769, 72.98951, 73.00162, 73.01321, 73.02431, 73.03488, 
    73.04494, 73.0545, 73.06354, 73.07206, 73.08007, 73.08756, 73.09454, 
    73.101, 73.10694, 73.11237, 73.11727, 73.12165, 73.12552, 73.12887, 
    73.13169, 73.134, 73.13577, 73.13704, 73.13778, 73.138, 73.1377, 
    73.13687, 73.13553, 73.13367, 73.13128, 73.12837, 73.12495, 73.12099, 
    73.11653, 73.11154, 73.10603, 73.10001, 73.09348, 73.08641, 73.07883, 
    73.07075, 73.06214, 73.05302, 73.04339, 73.03324, 73.02258, 73.01141, 
    72.99974, 72.98755, 72.97486, 72.96165, 72.94795, 72.93375, 72.91903, 
    72.90382, 72.88811, 72.87189, 72.85519, 72.83798, 72.82028, 72.80209, 
    72.78341, 72.76424, 72.74458, 72.72443, 72.7038, 72.68269, 72.66109, 
    72.63902, 72.61648, 72.59345, 72.56995, 72.54598, 72.52155, 72.49664, 
    72.47127, 72.44543, 72.41914, 72.39238, 72.36517, 72.3375, 72.30938, 
    72.28081, 72.25179, 72.22232, 72.19241, 72.16206, 72.13127, 72.10004, 
    72.06837, 72.03628, 72.00375, 71.9708, 71.93742, 71.90362, 71.8694, 
    71.83475, 71.7997, 71.76423, 71.72835, 71.69206, 71.65536, 71.61826, 
    71.58076, 71.54286, 71.50457, 71.46588, 71.4268, 71.38734, 71.34748, 
    71.30724, 71.26662, 71.22562, 71.18425, 71.14251, 71.10039, 71.0579, 
    71.01505, 70.97183, 70.92825, 70.88432, 70.84003, 70.79539, 70.75039, 
    70.70505, 70.65936, 70.61332, 70.56695, 70.52023, 70.47319, 70.4258, 
    70.37809, 70.33005, 70.28168, 70.23299, 70.18398, 70.13464, 70.085, 
    70.03503, 69.98476, 69.93418, 69.88329, 69.83209, 69.7806, 69.7288, 
    69.6767, 69.62432, 69.57164, 69.51867, 69.46541, 69.41186, 69.35803, 
    69.30392, 69.24953, 69.19486, 69.13992, 69.08471, 69.02923, 68.97348, 
    68.91746, 68.86118, 68.80463, 68.74783, 68.69078, 68.63346, 68.5759, 
    68.51808, 68.46001, 68.4017, 68.34314, 68.28434, 68.2253, 68.16602, 
    68.10651, 68.04676, 67.98678, 67.92656, 67.86612, 67.80545, 67.74455, 
    67.68344, 67.6221, 67.56055, 67.49877, 67.43678, 67.37457, 67.31216, 
    67.24953, 67.1867, 67.12366, 67.06042, 66.99697, 66.93332, 66.86947, 
    66.80543, 66.74118,
  60.18873, 60.26551, 60.3422, 60.4188, 60.49532, 60.57175, 60.64809, 
    60.72434, 60.8005, 60.87656, 60.95253, 61.02841, 61.10419, 61.17988, 
    61.25547, 61.33097, 61.40636, 61.48166, 61.55686, 61.63196, 61.70695, 
    61.78185, 61.85664, 61.93132, 62.00591, 62.08038, 62.15475, 62.22901, 
    62.30316, 62.3772, 62.45113, 62.52495, 62.59866, 62.67225, 62.74573, 
    62.81909, 62.89234, 62.96547, 63.03848, 63.11137, 63.18414, 63.25678, 
    63.32931, 63.40171, 63.47398, 63.54613, 63.61815, 63.69004, 63.76181, 
    63.83344, 63.90494, 63.97631, 64.04754, 64.11864, 64.1896, 64.26042, 
    64.3311, 64.40165, 64.47205, 64.5423, 64.61243, 64.6824, 64.75222, 
    64.82189, 64.89142, 64.96079, 65.03001, 65.09909, 65.16801, 65.23676, 
    65.30537, 65.37381, 65.44209, 65.51022, 65.57818, 65.64597, 65.7136, 
    65.78107, 65.84836, 65.91548, 65.98244, 66.04921, 66.11581, 66.18224, 
    66.2485, 66.31457, 66.38046, 66.44616, 66.51168, 66.57702, 66.64217, 
    66.70713, 66.7719, 66.83648, 66.90086, 66.96505, 67.02905, 67.09283, 
    67.15643, 67.21981, 67.283, 67.34597, 67.40874, 67.47131, 67.53365, 
    67.59579, 67.65771, 67.71941, 67.78089, 67.84216, 67.90319, 67.96401, 
    68.0246, 68.08496, 68.14509, 68.20499, 68.26465, 68.32407, 68.38326, 
    68.44221, 68.50092, 68.55937, 68.61759, 68.67555, 68.73327, 68.79073, 
    68.84794, 68.90488, 68.96157, 69.01801, 69.07417, 69.13007, 69.1857, 
    69.24106, 69.29614, 69.35096, 69.40549, 69.45975, 69.51373, 69.56742, 
    69.62083, 69.67394, 69.72677, 69.7793, 69.83154, 69.88348, 69.93512, 
    69.98646, 70.03749, 70.08822, 70.13863, 70.18874, 70.23853, 70.288, 
    70.33716, 70.38599, 70.43449, 70.48267, 70.53053, 70.57805, 70.62523, 
    70.67208, 70.71859, 70.76476, 70.81058, 70.85606, 70.90118, 70.94596, 
    70.99038, 71.03445, 71.07815, 71.12149, 71.16447, 71.20708, 71.24933, 
    71.2912, 71.3327, 71.37381, 71.41455, 71.4549, 71.49487, 71.53446, 
    71.57365, 71.61246, 71.65086, 71.68887, 71.72648, 71.76369, 71.80048, 
    71.83688, 71.87286, 71.90844, 71.9436, 71.97833, 72.01265, 72.04655, 
    72.08002, 72.11307, 72.14568, 72.17786, 72.20961, 72.24092, 72.2718, 
    72.30223, 72.33221, 72.36176, 72.39085, 72.41949, 72.44769, 72.47542, 
    72.5027, 72.52952, 72.55588, 72.58177, 72.6072, 72.63216, 72.65665, 
    72.68066, 72.70421, 72.72728, 72.74987, 72.77199, 72.79362, 72.81476, 
    72.83543, 72.8556, 72.87528, 72.89448, 72.91319, 72.9314, 72.94911, 
    72.96632, 72.98305, 72.99927, 73.01498, 73.0302, 73.04491, 73.05912, 
    73.07281, 73.08601, 73.09869, 73.11086, 73.12253, 73.13367, 73.14431, 
    73.15443, 73.16403, 73.17313, 73.18169, 73.18975, 73.19728, 73.2043, 
    73.21079, 73.21677, 73.22222, 73.22716, 73.23156, 73.23545, 73.23882, 
    73.24165, 73.24397, 73.24577, 73.24703, 73.24778, 73.248, 73.2477, 
    73.24686, 73.24551, 73.24364, 73.24124, 73.23832, 73.23487, 73.2309, 
    73.22641, 73.2214, 73.21586, 73.2098, 73.20322, 73.19613, 73.18851, 
    73.18037, 73.17172, 73.16255, 73.15286, 73.14266, 73.13194, 73.12071, 
    73.10897, 73.09672, 73.08395, 73.07069, 73.05691, 73.04262, 73.02782, 
    73.01254, 72.99673, 72.98044, 72.96364, 72.94634, 72.92854, 72.91026, 
    72.89148, 72.8722, 72.85244, 72.83218, 72.81145, 72.79022, 72.76852, 
    72.74633, 72.72366, 72.70052, 72.6769, 72.65281, 72.62824, 72.6032, 
    72.57771, 72.55173, 72.52531, 72.49841, 72.47106, 72.44326, 72.41499, 
    72.38628, 72.35712, 72.3275, 72.29745, 72.26694, 72.236, 72.20462, 
    72.1728, 72.14055, 72.10786, 72.07475, 72.04121, 72.00725, 71.97286, 
    71.93806, 71.90284, 71.8672, 71.83115, 71.79469, 71.75783, 71.72056, 
    71.68288, 71.64481, 71.60635, 71.56748, 71.52822, 71.48858, 71.44855, 
    71.40813, 71.36733, 71.32616, 71.2846, 71.24267, 71.20037, 71.1577, 
    71.11466, 71.07126, 71.0275, 70.98338, 70.9389, 70.89407, 70.84888, 
    70.80335, 70.75748, 70.71126, 70.66469, 70.61779, 70.57055, 70.52298, 
    70.47507, 70.42684, 70.37829, 70.3294, 70.2802, 70.23067, 70.18083, 
    70.13068, 70.08022, 70.02944, 69.97836, 69.92697, 69.87529, 69.8233, 
    69.77101, 69.71843, 69.66556, 69.6124, 69.55894, 69.50521, 69.45119, 
    69.39689, 69.34231, 69.28745, 69.23232, 69.17692, 69.12124, 69.0653, 
    69.00909, 68.95262, 68.8959, 68.83891, 68.78165, 68.72416, 68.6664, 
    68.6084, 68.55015, 68.49165, 68.4329, 68.37392, 68.31469, 68.25523, 
    68.19553, 68.13559, 68.07542, 68.01503, 67.95441, 67.89355, 67.83248, 
    67.77118, 67.70966, 67.64793, 67.58597, 67.5238, 67.46142, 67.39883, 
    67.33602, 67.27302, 67.2098, 67.14638, 67.08276, 67.01894, 66.95491, 
    66.89069, 66.82628 ;

 rlat = -24.032, -23.922, -23.812, -23.702, -23.592, -23.482, -23.372, 
    -23.262, -23.152, -23.042, -22.932, -22.822, -22.712, -22.602, -22.492, 
    -22.382, -22.272, -22.162, -22.052, -21.942, -21.832, -21.722, -21.612, 
    -21.502, -21.392, -21.282, -21.172, -21.062, -20.952, -20.842, -20.732, 
    -20.622, -20.512, -20.402, -20.292, -20.182, -20.072, -19.962, -19.852, 
    -19.742, -19.632, -19.522, -19.412, -19.302, -19.192, -19.082, -18.972, 
    -18.862, -18.752, -18.642, -18.532, -18.422, -18.312, -18.202, -18.092, 
    -17.982, -17.872, -17.762, -17.652, -17.542, -17.432, -17.322, -17.212, 
    -17.102, -16.992, -16.882, -16.772, -16.662, -16.552, -16.442, -16.332, 
    -16.222, -16.112, -16.002, -15.892, -15.782, -15.672, -15.562, -15.452, 
    -15.342, -15.232, -15.122, -15.012, -14.902, -14.792, -14.682, -14.572, 
    -14.462, -14.352, -14.242, -14.132, -14.022, -13.912, -13.802, -13.692, 
    -13.582, -13.472, -13.362, -13.252, -13.142, -13.032, -12.922, -12.812, 
    -12.702, -12.592, -12.482, -12.372, -12.262, -12.152, -12.042, -11.932, 
    -11.822, -11.712, -11.602, -11.492, -11.382, -11.272, -11.162, -11.052, 
    -10.942, -10.832, -10.722, -10.612, -10.502, -10.392, -10.282, -10.172, 
    -10.062, -9.952, -9.842, -9.732, -9.622, -9.512, -9.402, -9.292, -9.182, 
    -9.072, -8.962, -8.852, -8.742, -8.632, -8.522, -8.412, -8.302, -8.192, 
    -8.082, -7.972, -7.862, -7.752, -7.642, -7.532, -7.422, -7.312, -7.202, 
    -7.092, -6.982, -6.872, -6.762, -6.652, -6.542, -6.432, -6.322, -6.212, 
    -6.102, -5.992, -5.882, -5.772, -5.662, -5.552, -5.442, -5.332, -5.222, 
    -5.112, -5.002, -4.892, -4.782, -4.672, -4.562, -4.452, -4.342, -4.232, 
    -4.122, -4.012, -3.902, -3.792, -3.682, -3.572, -3.462, -3.352, -3.242, 
    -3.132, -3.022, -2.912, -2.802, -2.692, -2.582, -2.472, -2.362, -2.252, 
    -2.142, -2.032, -1.922, -1.812, -1.702, -1.592, -1.482, -1.372, -1.262, 
    -1.152, -1.042, -0.932, -0.822, -0.712, -0.602, -0.492, -0.382, -0.272, 
    -0.162, -0.052, 0.058, 0.168, 0.278, 0.388, 0.498, 0.608, 0.718, 0.828, 
    0.938, 1.048, 1.158, 1.268, 1.378, 1.488, 1.598, 1.708, 1.818, 1.928, 
    2.038, 2.148, 2.258, 2.368, 2.478, 2.588, 2.698, 2.808, 2.918, 3.028, 
    3.138, 3.248, 3.358, 3.468, 3.578, 3.688, 3.798, 3.908, 4.018, 4.128, 
    4.238, 4.348, 4.458, 4.568, 4.678, 4.788, 4.898, 5.008, 5.118, 5.228, 
    5.338, 5.448, 5.558, 5.668, 5.778, 5.888, 5.998, 6.108, 6.218, 6.328, 
    6.438, 6.548, 6.658, 6.768, 6.878, 6.988, 7.098, 7.208, 7.318, 7.428, 
    7.538, 7.648, 7.758, 7.868, 7.978, 8.088, 8.198, 8.308, 8.418, 8.528, 
    8.638, 8.748, 8.858, 8.968, 9.078, 9.188, 9.298, 9.408, 9.518, 9.628, 
    9.738, 9.848, 9.958, 10.068, 10.178, 10.288, 10.398, 10.508, 10.618, 
    10.728, 10.838, 10.948, 11.058, 11.168, 11.278, 11.388, 11.498, 11.608, 
    11.718, 11.828, 11.938, 12.048, 12.158, 12.268, 12.378, 12.488, 12.598, 
    12.708, 12.818, 12.928, 13.038, 13.148, 13.258, 13.368, 13.478, 13.588, 
    13.698, 13.808, 13.918, 14.028, 14.138, 14.248, 14.358, 14.468, 14.578, 
    14.688, 14.798, 14.908, 15.018, 15.128, 15.238, 15.348, 15.458, 15.568, 
    15.678, 15.788, 15.898, 16.008, 16.118, 16.228, 16.338, 16.448, 16.558, 
    16.668, 16.778, 16.888, 16.998, 17.108, 17.218, 17.328, 17.438, 17.548, 
    17.658, 17.768, 17.878, 17.988, 18.098, 18.208, 18.318, 18.428, 18.538, 
    18.648, 18.758, 18.868, 18.978, 19.088, 19.198, 19.308, 19.418, 19.528, 
    19.638, 19.748, 19.858, 19.968, 20.078, 20.188, 20.298, 20.408, 20.518, 
    20.628, 20.738, 20.848, 20.958, 21.068, 21.178, 21.288, 21.398, 21.508, 
    21.618, 21.728, 21.838, 21.948, 22.058, 22.168, 22.278, 22.388, 22.498 ;

 rotated_pole = 1 ;

 rlon = -29.0313, -28.9213, -28.8113, -28.7013, -28.5913, -28.4813, -28.3713, 
    -28.2613, -28.1513, -28.0413, -27.9313, -27.8213, -27.7113, -27.6013, 
    -27.4913, -27.3813, -27.2713, -27.1613, -27.0513, -26.9413, -26.8313, 
    -26.7213, -26.6113, -26.5013, -26.3913, -26.2813, -26.1713, -26.0613, 
    -25.9513, -25.8413, -25.7313, -25.6213, -25.5113, -25.4013, -25.2913, 
    -25.1813, -25.0713, -24.9613, -24.8513, -24.7413, -24.6313, -24.5213, 
    -24.4113, -24.3013, -24.1913, -24.0813, -23.9713, -23.8613, -23.7513, 
    -23.6413, -23.5313, -23.4213, -23.3113, -23.2013, -23.0913, -22.9813, 
    -22.8713, -22.7613, -22.6513, -22.5413, -22.4313, -22.3213, -22.2113, 
    -22.1013, -21.9913, -21.8813, -21.7713, -21.6613, -21.5513, -21.4413, 
    -21.3313, -21.2213, -21.1113, -21.0013, -20.8913, -20.7813, -20.6713, 
    -20.5613, -20.4513, -20.3413, -20.2313, -20.1213, -20.0113, -19.9013, 
    -19.7913, -19.6813, -19.5713, -19.4613, -19.3513, -19.2413, -19.1313, 
    -19.0213, -18.9113, -18.8013, -18.6913, -18.5813, -18.4713, -18.3613, 
    -18.2513, -18.1413, -18.0313, -17.9213, -17.8113, -17.7013, -17.5913, 
    -17.4813, -17.3713, -17.2613, -17.1513, -17.0413, -16.9313, -16.8213, 
    -16.7113, -16.6013, -16.4913, -16.3813, -16.2713, -16.1613, -16.0513, 
    -15.9413, -15.8313, -15.7213, -15.6113, -15.5013, -15.3913, -15.2813, 
    -15.1713, -15.0613, -14.9513, -14.8413, -14.7313, -14.6213, -14.5113, 
    -14.4013, -14.2913, -14.1813, -14.0713, -13.9613, -13.8513, -13.7413, 
    -13.6313, -13.5213, -13.4113, -13.3013, -13.1913, -13.0813, -12.9713, 
    -12.8613, -12.7513, -12.6413, -12.5313, -12.4213, -12.3113, -12.2013, 
    -12.0913, -11.9813, -11.8713, -11.7613, -11.6513, -11.5413, -11.4313, 
    -11.3213, -11.2113, -11.1013, -10.9913, -10.8813, -10.7713, -10.6613, 
    -10.5513, -10.4413, -10.3313, -10.2213, -10.1113, -10.0013, -9.8913, 
    -9.7813, -9.6713, -9.5613, -9.4513, -9.3413, -9.2313, -9.1213, -9.0113, 
    -8.9013, -8.7913, -8.6813, -8.5713, -8.4613, -8.3513, -8.2413, -8.1313, 
    -8.0213, -7.9113, -7.8013, -7.6913, -7.5813, -7.4713, -7.3613, -7.2513, 
    -7.1413, -7.0313, -6.9213, -6.8113, -6.7013, -6.5913, -6.4813, -6.3713, 
    -6.2613, -6.1513, -6.0413, -5.9313, -5.8213, -5.7113, -5.6013, -5.4913, 
    -5.3813, -5.2713, -5.1613, -5.0513, -4.9413, -4.8313, -4.7213, -4.6113, 
    -4.5013, -4.3913, -4.2813, -4.1713, -4.0613, -3.9513, -3.8413, -3.7313, 
    -3.6213, -3.5113, -3.4013, -3.2913, -3.1813, -3.0713, -2.9613, -2.8513, 
    -2.7413, -2.6313, -2.5213, -2.4113, -2.3013, -2.1913, -2.0813, -1.9713, 
    -1.8613, -1.7513, -1.6413, -1.5313, -1.4213, -1.3113, -1.2013, -1.0913, 
    -0.9813, -0.8713, -0.7613, -0.6513, -0.5413, -0.4313, -0.3213, -0.2113, 
    -0.1013, 0.0087, 0.1187, 0.2287, 0.3387, 0.4487, 0.5587, 0.6687, 0.7787, 
    0.8887, 0.9987, 1.1087, 1.2187, 1.3287, 1.4387, 1.5487, 1.6587, 1.7687, 
    1.8787, 1.9887, 2.0987, 2.2087, 2.3187, 2.4287, 2.5387, 2.6487, 2.7587, 
    2.8687, 2.9787, 3.0887, 3.1987, 3.3087, 3.4187, 3.5287, 3.6387, 3.7487, 
    3.8587, 3.9687, 4.0787, 4.1887, 4.2987, 4.4087, 4.5187, 4.6287, 4.7387, 
    4.8487, 4.9587, 5.0687, 5.1787, 5.2887, 5.3987, 5.5087, 5.6187, 5.7287, 
    5.8387, 5.9487, 6.0587, 6.1687, 6.2787, 6.3887, 6.4987, 6.6087, 6.7187, 
    6.8287, 6.9387, 7.0487, 7.1587, 7.2687, 7.3787, 7.4887, 7.5987, 7.7087, 
    7.8187, 7.9287, 8.0387, 8.1487, 8.2587, 8.3687, 8.4787, 8.5887, 8.6987, 
    8.8087, 8.9187, 9.0287, 9.1387, 9.2487, 9.3587, 9.4687, 9.5787, 9.6887, 
    9.7987, 9.9087, 10.0187, 10.1287, 10.2387, 10.3487, 10.4587, 10.5687, 
    10.6787, 10.7887, 10.8987, 11.0087, 11.1187, 11.2287, 11.3387, 11.4487, 
    11.5587, 11.6687, 11.7787, 11.8887, 11.9987, 12.1087, 12.2187, 12.3287, 
    12.4387, 12.5487, 12.6587, 12.7687, 12.8787, 12.9887, 13.0987, 13.2087, 
    13.3187, 13.4287, 13.5387, 13.6487, 13.7587, 13.8687, 13.9787, 14.0887, 
    14.1987, 14.3087, 14.4187, 14.5287, 14.6387, 14.7487, 14.8587, 14.9687, 
    15.0787, 15.1887, 15.2987, 15.4087, 15.5187, 15.6287, 15.7387, 15.8487, 
    15.9587, 16.0687, 16.1787, 16.2887, 16.3987, 16.5087, 16.6187, 16.7287, 
    16.8387, 16.9487, 17.0587, 17.1687, 17.2787, 17.3887, 17.4987, 17.6087, 
    17.7187, 17.8287, 17.9387, 18.0487, 18.1587, 18.2687, 18.3787, 18.4887, 
    18.5987, 18.7087, 18.8187 ;
}
